library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;
use ieee.numeric_std.all;    
--USE ieee.std_logic_arith.all;

entity Entropy_encoding is
  generic (
           mult_sum_CL   : string := "sum";
           mult_sum_PCA  : string := "sum";
           N             : integer :=   8; -- input data width
           Huff_wid      : integer :=  12; -- Huffman weight maximum width                   (after change need nedd to update "Huff_code" matrix)
           Wh            : integer :=  16; -- Huffman unit output data width (Note W>=M)
           Wb            : integer := 128; -- output buffer data width
           depth         : integer :=  64; -- buffer depth
           burst         : integer :=  10; -- buffer read burst
 
           PCA_en        : boolean := TRUE; --TRUE; -- PCA Enable/Bypass
           Huff_enc_en   : boolean := TRUE;--FALSE; -- Huffman encoder Enable/Bypass

  	       in_row        : integer := 114;
  	       in_col        : integer := 114
  	       );
  port    (
           clk       : in  std_logic;
           rst       : in  std_logic;

           pca_w_en  : in  std_logic;
           pca_w_num : in  std_logic_vector (6 downto 0);
           pca_w_in  : in  std_logic_vector (7 downto 0);

  	       d_in      : in  std_logic_vector (N-1 downto 0);
  	       en_in     : in  std_logic;
  	       sof_in    : in  std_logic; -- start of frame
  	       --sol     : in  std_logic; -- start of line
  	       --eof     : in  std_logic; -- end of frame

           buf_rd    : in  std_logic;
           buf_num   : in  std_logic_vector (6      downto 0);
           d_out     : out std_logic_vector (Wb  -1 downto 0);
           en_out    : out std_logic_vector (64  -1 downto 0);
           sof_out   : out std_logic);
end Entropy_encoding;

architecture a of Entropy_encoding is

constant PCAweightW   : integer := 8;

component ConvLayer128 is
  generic (
           mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width
           SR            : integer := 8; -- data shift right before output
           --bpp           : integer := 8; -- bit per pixel
           in_row        : integer := 8;
           in_col        : integer := 8
           );
  port    (
           clk     : in std_logic;
           rst     : in std_logic;
           d_in    : in std_logic_vector (N-1 downto 0);
           en_in   : in std_logic;
           sof_in  : in std_logic; -- start of frame
           --sol     : in std_logic; -- start of line
           --eof     : in std_logic; -- end of frame
           w_in    : in std_logic_vector(M-1 downto 0);
           w_num   : in std_logic_vector(  3 downto 0);
           w_en    : in std_logic;

           d_out   : out std_logic_vector (W-1 downto 0);
           en_out  : out std_logic;
           sof_out : out std_logic);
end component;

component PCA_128 is
  generic (
           mult_sum      : string := "sum";
           N             : integer := 8;       -- input data width
           M             : integer := 8;       -- input weight width
           in_row        : integer := 256;
           in_col        : integer := 256
           );
  port    (
           clk     : in std_logic;
           rst     : in std_logic;
          -- d_in      : in std_logic_vector_vector(1 to 64)(N-1 downto 0);
           d01_in    : in std_logic_vector (N-1 downto 0);
           d02_in    : in std_logic_vector (N-1 downto 0);
           d03_in    : in std_logic_vector (N-1 downto 0);
           d04_in    : in std_logic_vector (N-1 downto 0);
           d05_in    : in std_logic_vector (N-1 downto 0);
           d06_in    : in std_logic_vector (N-1 downto 0);
           d07_in    : in std_logic_vector (N-1 downto 0);
           d08_in    : in std_logic_vector (N-1 downto 0);
           d09_in    : in std_logic_vector (N-1 downto 0);
           d10_in    : in std_logic_vector (N-1 downto 0);
           d11_in    : in std_logic_vector (N-1 downto 0);
           d12_in    : in std_logic_vector (N-1 downto 0);
           d13_in    : in std_logic_vector (N-1 downto 0);
           d14_in    : in std_logic_vector (N-1 downto 0);
           d15_in    : in std_logic_vector (N-1 downto 0);
           d16_in    : in std_logic_vector (N-1 downto 0);
           d17_in    : in std_logic_vector (N-1 downto 0);
           d18_in    : in std_logic_vector (N-1 downto 0);
           d19_in    : in std_logic_vector (N-1 downto 0);
           d20_in    : in std_logic_vector (N-1 downto 0);
           d21_in    : in std_logic_vector (N-1 downto 0);
           d22_in    : in std_logic_vector (N-1 downto 0);
           d23_in    : in std_logic_vector (N-1 downto 0);
           d24_in    : in std_logic_vector (N-1 downto 0);
           d25_in    : in std_logic_vector (N-1 downto 0);
           d26_in    : in std_logic_vector (N-1 downto 0);
           d27_in    : in std_logic_vector (N-1 downto 0);
           d28_in    : in std_logic_vector (N-1 downto 0);
           d29_in    : in std_logic_vector (N-1 downto 0);
           d30_in    : in std_logic_vector (N-1 downto 0);
           d31_in    : in std_logic_vector (N-1 downto 0);
           d32_in    : in std_logic_vector (N-1 downto 0);
           d33_in    : in std_logic_vector (N-1 downto 0);
           d34_in    : in std_logic_vector (N-1 downto 0);
           d35_in    : in std_logic_vector (N-1 downto 0);
           d36_in    : in std_logic_vector (N-1 downto 0);
           d37_in    : in std_logic_vector (N-1 downto 0);
           d38_in    : in std_logic_vector (N-1 downto 0);
           d39_in    : in std_logic_vector (N-1 downto 0);
           d40_in    : in std_logic_vector (N-1 downto 0);
           d41_in    : in std_logic_vector (N-1 downto 0);
           d42_in    : in std_logic_vector (N-1 downto 0);
           d43_in    : in std_logic_vector (N-1 downto 0);
           d44_in    : in std_logic_vector (N-1 downto 0);
           d45_in    : in std_logic_vector (N-1 downto 0);
           d46_in    : in std_logic_vector (N-1 downto 0);
           d47_in    : in std_logic_vector (N-1 downto 0);
           d48_in    : in std_logic_vector (N-1 downto 0);
           d49_in    : in std_logic_vector (N-1 downto 0);
           d50_in    : in std_logic_vector (N-1 downto 0);
           d51_in    : in std_logic_vector (N-1 downto 0);
           d52_in    : in std_logic_vector (N-1 downto 0);
           d53_in    : in std_logic_vector (N-1 downto 0);
           d54_in    : in std_logic_vector (N-1 downto 0);
           d55_in    : in std_logic_vector (N-1 downto 0);
           d56_in    : in std_logic_vector (N-1 downto 0);
           d57_in    : in std_logic_vector (N-1 downto 0);
           d58_in    : in std_logic_vector (N-1 downto 0);
           d59_in    : in std_logic_vector (N-1 downto 0);
           d60_in    : in std_logic_vector (N-1 downto 0);
           d61_in    : in std_logic_vector (N-1 downto 0);
           d62_in    : in std_logic_vector (N-1 downto 0);
           d63_in    : in std_logic_vector (N-1 downto 0);
           d64_in    : in std_logic_vector (N-1 downto 0);

           d65_in    : in std_logic_vector (N-1 downto 0);
           d66_in    : in std_logic_vector (N-1 downto 0);
           d67_in    : in std_logic_vector (N-1 downto 0);
           d68_in    : in std_logic_vector (N-1 downto 0);
           d69_in    : in std_logic_vector (N-1 downto 0);
           d70_in    : in std_logic_vector (N-1 downto 0);
           d71_in    : in std_logic_vector (N-1 downto 0);
           d72_in    : in std_logic_vector (N-1 downto 0);
           d73_in    : in std_logic_vector (N-1 downto 0);
           d74_in    : in std_logic_vector (N-1 downto 0);
           d75_in    : in std_logic_vector (N-1 downto 0);
           d76_in    : in std_logic_vector (N-1 downto 0);
           d77_in    : in std_logic_vector (N-1 downto 0);
           d78_in    : in std_logic_vector (N-1 downto 0);
           d79_in    : in std_logic_vector (N-1 downto 0);
           d80_in    : in std_logic_vector (N-1 downto 0);
           d81_in    : in std_logic_vector (N-1 downto 0);
           d82_in    : in std_logic_vector (N-1 downto 0);
           d83_in    : in std_logic_vector (N-1 downto 0);
           d84_in    : in std_logic_vector (N-1 downto 0);
           d85_in    : in std_logic_vector (N-1 downto 0);
           d86_in    : in std_logic_vector (N-1 downto 0);
           d87_in    : in std_logic_vector (N-1 downto 0);
           d88_in    : in std_logic_vector (N-1 downto 0);
           d89_in    : in std_logic_vector (N-1 downto 0);
           d90_in    : in std_logic_vector (N-1 downto 0);
           d91_in    : in std_logic_vector (N-1 downto 0);
           d92_in    : in std_logic_vector (N-1 downto 0);
           d93_in    : in std_logic_vector (N-1 downto 0);
           d94_in    : in std_logic_vector (N-1 downto 0);
           d95_in    : in std_logic_vector (N-1 downto 0);
           d96_in    : in std_logic_vector (N-1 downto 0);
           d97_in    : in std_logic_vector (N-1 downto 0);
           d98_in    : in std_logic_vector (N-1 downto 0);
           d99_in    : in std_logic_vector (N-1 downto 0);
           d100_in    : in std_logic_vector (N-1 downto 0);
           d101_in    : in std_logic_vector (N-1 downto 0);
           d102_in    : in std_logic_vector (N-1 downto 0);
           d103_in    : in std_logic_vector (N-1 downto 0);
           d104_in    : in std_logic_vector (N-1 downto 0);
           d105_in    : in std_logic_vector (N-1 downto 0);
           d106_in    : in std_logic_vector (N-1 downto 0);
           d107_in    : in std_logic_vector (N-1 downto 0);
           d108_in    : in std_logic_vector (N-1 downto 0);
           d109_in    : in std_logic_vector (N-1 downto 0);
           d110_in    : in std_logic_vector (N-1 downto 0);
           d111_in    : in std_logic_vector (N-1 downto 0);
           d112_in    : in std_logic_vector (N-1 downto 0);
           d113_in    : in std_logic_vector (N-1 downto 0);
           d114_in    : in std_logic_vector (N-1 downto 0);
           d115_in    : in std_logic_vector (N-1 downto 0);
           d116_in    : in std_logic_vector (N-1 downto 0);
           d117_in    : in std_logic_vector (N-1 downto 0);
           d118_in    : in std_logic_vector (N-1 downto 0);
           d119_in    : in std_logic_vector (N-1 downto 0);
           d120_in    : in std_logic_vector (N-1 downto 0);
           d121_in    : in std_logic_vector (N-1 downto 0);
           d122_in    : in std_logic_vector (N-1 downto 0);
           d123_in    : in std_logic_vector (N-1 downto 0);
           d124_in    : in std_logic_vector (N-1 downto 0);
           d125_in    : in std_logic_vector (N-1 downto 0);
           d126_in    : in std_logic_vector (N-1 downto 0);
           d127_in    : in std_logic_vector (N-1 downto 0);
           d128_in    : in std_logic_vector (N-1 downto 0);

           en_in     : in std_logic;
           sof_in    : in std_logic; -- start of frame

           w01      : in std_logic_vector(M-1 downto 0); 
           w02      : in std_logic_vector(M-1 downto 0); 
           w03      : in std_logic_vector(M-1 downto 0); 
           w04      : in std_logic_vector(M-1 downto 0); 
           w05      : in std_logic_vector(M-1 downto 0); 
           w06      : in std_logic_vector(M-1 downto 0); 
           w07      : in std_logic_vector(M-1 downto 0); 
           w08      : in std_logic_vector(M-1 downto 0); 
           w09      : in std_logic_vector(M-1 downto 0); 
           w10      : in std_logic_vector(M-1 downto 0); 
           w11      : in std_logic_vector(M-1 downto 0); 
           w12      : in std_logic_vector(M-1 downto 0); 
           w13      : in std_logic_vector(M-1 downto 0); 
           w14      : in std_logic_vector(M-1 downto 0); 
           w15      : in std_logic_vector(M-1 downto 0); 
           w16      : in std_logic_vector(M-1 downto 0); 
           w17      : in std_logic_vector(M-1 downto 0); 
           w18      : in std_logic_vector(M-1 downto 0); 
           w19      : in std_logic_vector(M-1 downto 0); 
           w20      : in std_logic_vector(M-1 downto 0); 
           w21      : in std_logic_vector(M-1 downto 0); 
           w22      : in std_logic_vector(M-1 downto 0); 
           w23      : in std_logic_vector(M-1 downto 0); 
           w24      : in std_logic_vector(M-1 downto 0); 
           w25      : in std_logic_vector(M-1 downto 0); 
           w26      : in std_logic_vector(M-1 downto 0); 
           w27      : in std_logic_vector(M-1 downto 0); 
           w28      : in std_logic_vector(M-1 downto 0); 
           w29      : in std_logic_vector(M-1 downto 0); 
           w30      : in std_logic_vector(M-1 downto 0); 
           w31      : in std_logic_vector(M-1 downto 0); 
           w32      : in std_logic_vector(M-1 downto 0); 
           w33      : in std_logic_vector(M-1 downto 0); 
           w34      : in std_logic_vector(M-1 downto 0); 
           w35      : in std_logic_vector(M-1 downto 0); 
           w36      : in std_logic_vector(M-1 downto 0); 
           w37      : in std_logic_vector(M-1 downto 0); 
           w38      : in std_logic_vector(M-1 downto 0); 
           w39      : in std_logic_vector(M-1 downto 0); 
           w40      : in std_logic_vector(M-1 downto 0); 
           w41      : in std_logic_vector(M-1 downto 0); 
           w42      : in std_logic_vector(M-1 downto 0); 
           w43      : in std_logic_vector(M-1 downto 0); 
           w44      : in std_logic_vector(M-1 downto 0); 
           w45      : in std_logic_vector(M-1 downto 0); 
           w46      : in std_logic_vector(M-1 downto 0); 
           w47      : in std_logic_vector(M-1 downto 0); 
           w48      : in std_logic_vector(M-1 downto 0); 
           w49      : in std_logic_vector(M-1 downto 0); 
           w50      : in std_logic_vector(M-1 downto 0); 
           w51      : in std_logic_vector(M-1 downto 0); 
           w52      : in std_logic_vector(M-1 downto 0); 
           w53      : in std_logic_vector(M-1 downto 0); 
           w54      : in std_logic_vector(M-1 downto 0); 
           w55      : in std_logic_vector(M-1 downto 0); 
           w56      : in std_logic_vector(M-1 downto 0); 
           w57      : in std_logic_vector(M-1 downto 0); 
           w58      : in std_logic_vector(M-1 downto 0); 
           w59      : in std_logic_vector(M-1 downto 0); 
           w60      : in std_logic_vector(M-1 downto 0); 
           w61      : in std_logic_vector(M-1 downto 0); 
           w62      : in std_logic_vector(M-1 downto 0); 
           w63      : in std_logic_vector(M-1 downto 0); 
           w64      : in std_logic_vector(M-1 downto 0); 


           w65      : in std_logic_vector(M-1 downto 0); 
           w66      : in std_logic_vector(M-1 downto 0); 
           w67      : in std_logic_vector(M-1 downto 0); 
           w68      : in std_logic_vector(M-1 downto 0); 
           w69      : in std_logic_vector(M-1 downto 0); 
           w70      : in std_logic_vector(M-1 downto 0); 
           w71      : in std_logic_vector(M-1 downto 0); 
           w72      : in std_logic_vector(M-1 downto 0); 
           w73      : in std_logic_vector(M-1 downto 0); 
           w74      : in std_logic_vector(M-1 downto 0); 
           w75      : in std_logic_vector(M-1 downto 0); 
           w76      : in std_logic_vector(M-1 downto 0); 
           w77      : in std_logic_vector(M-1 downto 0); 
           w78      : in std_logic_vector(M-1 downto 0); 
           w79      : in std_logic_vector(M-1 downto 0); 
           w80      : in std_logic_vector(M-1 downto 0); 
           w81      : in std_logic_vector(M-1 downto 0); 
           w82      : in std_logic_vector(M-1 downto 0); 
           w83      : in std_logic_vector(M-1 downto 0); 
           w84      : in std_logic_vector(M-1 downto 0); 
           w85      : in std_logic_vector(M-1 downto 0); 
           w86      : in std_logic_vector(M-1 downto 0); 
           w87      : in std_logic_vector(M-1 downto 0); 
           w88      : in std_logic_vector(M-1 downto 0); 
           w89      : in std_logic_vector(M-1 downto 0); 
           w90      : in std_logic_vector(M-1 downto 0); 
           w91      : in std_logic_vector(M-1 downto 0); 
           w92      : in std_logic_vector(M-1 downto 0); 
           w93      : in std_logic_vector(M-1 downto 0); 
           w94      : in std_logic_vector(M-1 downto 0); 
           w95      : in std_logic_vector(M-1 downto 0); 
           w96      : in std_logic_vector(M-1 downto 0); 
           w97      : in std_logic_vector(M-1 downto 0); 
           w98      : in std_logic_vector(M-1 downto 0); 
           w99      : in std_logic_vector(M-1 downto 0); 
           w100      : in std_logic_vector(M-1 downto 0); 
           w101      : in std_logic_vector(M-1 downto 0); 
           w102      : in std_logic_vector(M-1 downto 0); 
           w103      : in std_logic_vector(M-1 downto 0); 
           w104      : in std_logic_vector(M-1 downto 0); 
           w105      : in std_logic_vector(M-1 downto 0); 
           w106      : in std_logic_vector(M-1 downto 0); 
           w107      : in std_logic_vector(M-1 downto 0); 
           w108      : in std_logic_vector(M-1 downto 0); 
           w109      : in std_logic_vector(M-1 downto 0); 
           w110      : in std_logic_vector(M-1 downto 0); 
           w111      : in std_logic_vector(M-1 downto 0); 
           w112      : in std_logic_vector(M-1 downto 0); 
           w113      : in std_logic_vector(M-1 downto 0); 
           w114      : in std_logic_vector(M-1 downto 0); 
           w115      : in std_logic_vector(M-1 downto 0); 
           w116      : in std_logic_vector(M-1 downto 0); 
           w117      : in std_logic_vector(M-1 downto 0); 
           w118      : in std_logic_vector(M-1 downto 0); 
           w119      : in std_logic_vector(M-1 downto 0); 
           w120      : in std_logic_vector(M-1 downto 0); 
           w121      : in std_logic_vector(M-1 downto 0); 
           w122      : in std_logic_vector(M-1 downto 0); 
           w123      : in std_logic_vector(M-1 downto 0); 
           w124      : in std_logic_vector(M-1 downto 0); 
           w125      : in std_logic_vector(M-1 downto 0); 
           w126      : in std_logic_vector(M-1 downto 0); 
           w127      : in std_logic_vector(M-1 downto 0); 
           w128      : in std_logic_vector(M-1 downto 0); 
           d_out   : out std_logic_vector (N + M + 5 downto 0);
           en_out  : out std_logic;
           sof_out : out std_logic);
end component;

component Huffman128 is
  generic (
           N             : integer := 4;  -- input data width
           M             : integer := 8;  -- max code width
           Wh            : integer := 16;  -- Huffman unit output data width (Note W>=M)
           Wb            : integer := 512; -- output buffer data width
           Huff_enc_en   : boolean := TRUE; -- Huffman encoder Enable/Bypass
           depth         : integer := 500; -- buffer depth
           burst         : integer := 10   -- buffer read burst
           );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           init_en       : in  std_logic;                         -- initialising convert table
           alpha_data    : in  std_logic_vector(N-1 downto 0);    
           alpha_code    : in  std_logic_vector(M-1 downto 0);    
           alpha_width   : in  std_logic_vector(  3 downto 0);

           d01_in          : in std_logic_vector (N-1 downto 0);
           d02_in          : in std_logic_vector (N-1 downto 0);
           d03_in          : in std_logic_vector (N-1 downto 0);
           d04_in          : in std_logic_vector (N-1 downto 0);
           d05_in          : in std_logic_vector (N-1 downto 0);
           d06_in          : in std_logic_vector (N-1 downto 0);
           d07_in          : in std_logic_vector (N-1 downto 0);
           d08_in          : in std_logic_vector (N-1 downto 0);
           d09_in          : in std_logic_vector (N-1 downto 0);
           d10_in          : in std_logic_vector (N-1 downto 0);
           d11_in          : in std_logic_vector (N-1 downto 0);
           d12_in          : in std_logic_vector (N-1 downto 0);
           d13_in          : in std_logic_vector (N-1 downto 0);
           d14_in          : in std_logic_vector (N-1 downto 0);
           d15_in          : in std_logic_vector (N-1 downto 0);
           d16_in          : in std_logic_vector (N-1 downto 0);
           d17_in          : in std_logic_vector (N-1 downto 0);
           d18_in          : in std_logic_vector (N-1 downto 0);
           d19_in          : in std_logic_vector (N-1 downto 0);
           d20_in          : in std_logic_vector (N-1 downto 0);
           d21_in          : in std_logic_vector (N-1 downto 0);
           d22_in          : in std_logic_vector (N-1 downto 0);
           d23_in          : in std_logic_vector (N-1 downto 0);
           d24_in          : in std_logic_vector (N-1 downto 0);
           d25_in          : in std_logic_vector (N-1 downto 0);
           d26_in          : in std_logic_vector (N-1 downto 0);
           d27_in          : in std_logic_vector (N-1 downto 0);
           d28_in          : in std_logic_vector (N-1 downto 0);
           d29_in          : in std_logic_vector (N-1 downto 0);
           d30_in          : in std_logic_vector (N-1 downto 0);
           d31_in          : in std_logic_vector (N-1 downto 0);
           d32_in          : in std_logic_vector (N-1 downto 0);
           d33_in          : in std_logic_vector (N-1 downto 0);
           d34_in          : in std_logic_vector (N-1 downto 0);
           d35_in          : in std_logic_vector (N-1 downto 0);
           d36_in          : in std_logic_vector (N-1 downto 0);
           d37_in          : in std_logic_vector (N-1 downto 0);
           d38_in          : in std_logic_vector (N-1 downto 0);
           d39_in          : in std_logic_vector (N-1 downto 0);
           d40_in          : in std_logic_vector (N-1 downto 0);
           d41_in          : in std_logic_vector (N-1 downto 0);
           d42_in          : in std_logic_vector (N-1 downto 0);
           d43_in          : in std_logic_vector (N-1 downto 0);
           d44_in          : in std_logic_vector (N-1 downto 0);
           d45_in          : in std_logic_vector (N-1 downto 0);
           d46_in          : in std_logic_vector (N-1 downto 0);
           d47_in          : in std_logic_vector (N-1 downto 0);
           d48_in          : in std_logic_vector (N-1 downto 0);
           d49_in          : in std_logic_vector (N-1 downto 0);
           d50_in          : in std_logic_vector (N-1 downto 0);
           d51_in          : in std_logic_vector (N-1 downto 0);
           d52_in          : in std_logic_vector (N-1 downto 0);
           d53_in          : in std_logic_vector (N-1 downto 0);
           d54_in          : in std_logic_vector (N-1 downto 0);
           d55_in          : in std_logic_vector (N-1 downto 0);
           d56_in          : in std_logic_vector (N-1 downto 0);
           d57_in          : in std_logic_vector (N-1 downto 0);
           d58_in          : in std_logic_vector (N-1 downto 0);
           d59_in          : in std_logic_vector (N-1 downto 0);
           d60_in          : in std_logic_vector (N-1 downto 0);
           d61_in          : in std_logic_vector (N-1 downto 0);
           d62_in          : in std_logic_vector (N-1 downto 0);
           d63_in          : in std_logic_vector (N-1 downto 0);
           d64_in          : in std_logic_vector (N-1 downto 0);

           d65_in          : in std_logic_vector (N-1 downto 0);
           d66_in          : in std_logic_vector (N-1 downto 0);
           d67_in          : in std_logic_vector (N-1 downto 0);
           d68_in          : in std_logic_vector (N-1 downto 0);
           d69_in          : in std_logic_vector (N-1 downto 0);
           d70_in          : in std_logic_vector (N-1 downto 0);
           d71_in          : in std_logic_vector (N-1 downto 0);
           d72_in          : in std_logic_vector (N-1 downto 0);
           d73_in          : in std_logic_vector (N-1 downto 0);
           d74_in          : in std_logic_vector (N-1 downto 0);
           d75_in          : in std_logic_vector (N-1 downto 0);
           d76_in          : in std_logic_vector (N-1 downto 0);
           d77_in          : in std_logic_vector (N-1 downto 0);
           d78_in          : in std_logic_vector (N-1 downto 0);
           d79_in          : in std_logic_vector (N-1 downto 0);
           d80_in          : in std_logic_vector (N-1 downto 0);
           d81_in          : in std_logic_vector (N-1 downto 0);
           d82_in          : in std_logic_vector (N-1 downto 0);
           d83_in          : in std_logic_vector (N-1 downto 0);
           d84_in          : in std_logic_vector (N-1 downto 0);
           d85_in          : in std_logic_vector (N-1 downto 0);
           d86_in          : in std_logic_vector (N-1 downto 0);
           d87_in          : in std_logic_vector (N-1 downto 0);
           d88_in          : in std_logic_vector (N-1 downto 0);
           d89_in          : in std_logic_vector (N-1 downto 0);
           d90_in          : in std_logic_vector (N-1 downto 0);
           d91_in          : in std_logic_vector (N-1 downto 0);
           d92_in          : in std_logic_vector (N-1 downto 0);
           d93_in          : in std_logic_vector (N-1 downto 0);
           d94_in          : in std_logic_vector (N-1 downto 0);
           d95_in          : in std_logic_vector (N-1 downto 0);
           d96_in          : in std_logic_vector (N-1 downto 0);
           d97_in          : in std_logic_vector (N-1 downto 0);
           d98_in          : in std_logic_vector (N-1 downto 0);
           d99_in          : in std_logic_vector (N-1 downto 0);
           d100_in         : in std_logic_vector (N-1 downto 0);
           d101_in         : in std_logic_vector (N-1 downto 0);
           d102_in         : in std_logic_vector (N-1 downto 0);
           d103_in         : in std_logic_vector (N-1 downto 0);
           d104_in         : in std_logic_vector (N-1 downto 0);
           d105_in         : in std_logic_vector (N-1 downto 0);
           d106_in         : in std_logic_vector (N-1 downto 0);
           d107_in         : in std_logic_vector (N-1 downto 0);
           d108_in         : in std_logic_vector (N-1 downto 0);
           d109_in         : in std_logic_vector (N-1 downto 0);
           d110_in         : in std_logic_vector (N-1 downto 0);
           d111_in         : in std_logic_vector (N-1 downto 0);
           d112_in         : in std_logic_vector (N-1 downto 0);
           d113_in         : in std_logic_vector (N-1 downto 0);
           d114_in         : in std_logic_vector (N-1 downto 0);
           d115_in         : in std_logic_vector (N-1 downto 0);
           d116_in         : in std_logic_vector (N-1 downto 0);
           d117_in         : in std_logic_vector (N-1 downto 0);
           d118_in         : in std_logic_vector (N-1 downto 0);
           d119_in         : in std_logic_vector (N-1 downto 0);
           d120_in         : in std_logic_vector (N-1 downto 0);
           d121_in         : in std_logic_vector (N-1 downto 0);
           d122_in         : in std_logic_vector (N-1 downto 0);
           d123_in         : in std_logic_vector (N-1 downto 0);
           d124_in         : in std_logic_vector (N-1 downto 0);
           d125_in         : in std_logic_vector (N-1 downto 0);
           d126_in         : in std_logic_vector (N-1 downto 0);
           d127_in         : in std_logic_vector (N-1 downto 0);
           d128_in         : in std_logic_vector (N-1 downto 0);

           en_in         : in  std_logic;
           sof_in        : in  std_logic;                         -- start of frame
           eof_in        : in  std_logic;                         -- end of frame

           buf_rd        : in  std_logic;
           buf_num       : in  std_logic_vector (6      downto 0);
           d_out         : out std_logic_vector (Wb  -1 downto 0);
           en_out        : out std_logic_vector (128  -1 downto 0);
           eof_out       : out std_logic);                        -- huffman code output
end component;

constant CL_w_width : integer := 8;
type rom_type is array ( 0 to 15 ) of std_logic_vector(CL_w_width-1 downto 0 ) ;

constant weight01 : rom_type := ( 0 => x"00", 1 => x"17", 2 => x"92", 3 => x"14", 4 => x"61", 5 => x"27", 6 => x"53", 7 => x"60", 8 => x"11", 9 => x"61", others => x"00"); 
constant weight02 : rom_type := ( 0 => x"00", 1 => x"35", 2 => x"40", 3 => x"10", 4 => x"87", 5 => x"96", 6 => x"39", 7 => x"66", 8 => x"98", 9 => x"51", others => x"00"); 
constant weight03 : rom_type := ( 0 => x"00", 1 => x"85", 2 => x"48", 3 => x"56", 4 => x"67", 5 => x"82", 6 => x"28", 7 => x"70", 8 => x"72", 9 => x"58", others => x"00"); 
constant weight04 : rom_type := ( 0 => x"00", 1 => x"93", 2 => x"41", 3 => x"26", 4 => x"13", 5 => x"77", 6 => x"10", 7 => x"83", 8 => x"66", 9 => x"44", others => x"00"); 
constant weight05 : rom_type := ( 0 => x"00", 1 => x"88", 2 => x"82", 3 => x"74", 4 => x"24", 5 => x"10", 6 => x"41", 7 => x"99", 8 => x"61", 9 => x"53", others => x"00"); 
constant weight06 : rom_type := ( 0 => x"00", 1 => x"48", 2 => x"64", 3 => x"38", 4 => x"89", 5 => x"84", 6 => x"83", 7 => x"89", 8 => x"58", 9 => x"47", others => x"00"); 
constant weight07 : rom_type := ( 0 => x"00", 1 => x"35", 2 => x"79", 3 => x"73", 4 => x"99", 5 => x"67", 6 => x"26", 7 => x"82", 8 => x"39", 9 => x"49", others => x"00"); 
constant weight08 : rom_type := ( 0 => x"00", 1 => x"24", 2 => x"61", 3 => x"52", 4 => x"55", 5 => x"18", 6 => x"66", 7 => x"46", 8 => x"91", 9 => x"56", others => x"00"); 
constant weight09 : rom_type := ( 0 => x"00", 1 => x"43", 2 => x"16", 3 => x"32", 4 => x"43", 5 => x"81", 6 => x"49", 7 => x"99", 8 => x"51", 9 => x"42", others => x"00"); 
constant weight10 : rom_type := ( 0 => x"00", 1 => x"21", 2 => x"70", 3 => x"90", 4 => x"23", 5 => x"19", 6 => x"36", 7 => x"92", 8 => x"64", 9 => x"34", others => x"00"); 
constant weight11 : rom_type := ( 0 => x"00", 1 => x"19", 2 => x"70", 3 => x"58", 4 => x"17", 5 => x"49", 6 => x"28", 7 => x"34", 8 => x"28", 9 => x"78", others => x"00"); 
constant weight12 : rom_type := ( 0 => x"00", 1 => x"34", 2 => x"54", 3 => x"61", 4 => x"29", 5 => x"42", 6 => x"61", 7 => x"35", 8 => x"90", 9 => x"59", others => x"00"); 
constant weight13 : rom_type := ( 0 => x"00", 1 => x"23", 2 => x"20", 3 => x"51", 4 => x"10", 5 => x"83", 6 => x"64", 7 => x"24", 8 => x"15", 9 => x"69", others => x"00"); 
constant weight14 : rom_type := ( 0 => x"00", 1 => x"33", 2 => x"35", 3 => x"38", 4 => x"42", 5 => x"13", 6 => x"20", 7 => x"52", 8 => x"54", 9 => x"87", others => x"00"); 
constant weight15 : rom_type := ( 0 => x"00", 1 => x"11", 2 => x"11", 3 => x"77", 4 => x"58", 5 => x"54", 6 => x"55", 7 => x"12", 8 => x"13", 9 => x"53", others => x"00"); 
constant weight16 : rom_type := ( 0 => x"00", 1 => x"47", 2 => x"60", 3 => x"59", 4 => x"65", 5 => x"44", 6 => x"70", 7 => x"82", 8 => x"36", 9 => x"92", others => x"00"); 
constant weight17 : rom_type := ( 0 => x"00", 1 => x"35", 2 => x"94", 3 => x"56", 4 => x"40", 5 => x"16", 6 => x"76", 7 => x"46", 8 => x"72", 9 => x"36", others => x"00"); 
constant weight18 : rom_type := ( 0 => x"00", 1 => x"39", 2 => x"84", 3 => x"41", 4 => x"67", 5 => x"62", 6 => x"87", 7 => x"97", 8 => x"67", 9 => x"65", others => x"00"); 
constant weight19 : rom_type := ( 0 => x"00", 1 => x"96", 2 => x"96", 3 => x"12", 4 => x"91", 5 => x"98", 6 => x"46", 7 => x"50", 8 => x"77", 9 => x"60", others => x"00"); 
constant weight20 : rom_type := ( 0 => x"00", 1 => x"89", 2 => x"89", 3 => x"27", 4 => x"56", 5 => x"79", 6 => x"69", 7 => x"20", 8 => x"34", 9 => x"73", others => x"00"); 
constant weight21 : rom_type := ( 0 => x"00", 1 => x"61", 2 => x"79", 3 => x"15", 4 => x"36", 5 => x"10", 6 => x"71", 7 => x"41", 8 => x"35", 9 => x"34", others => x"00"); 
constant weight22 : rom_type := ( 0 => x"00", 1 => x"59", 2 => x"97", 3 => x"32", 4 => x"56", 5 => x"69", 6 => x"70", 7 => x"41", 8 => x"87", 9 => x"40", others => x"00"); 
constant weight23 : rom_type := ( 0 => x"00", 1 => x"32", 2 => x"19", 3 => x"63", 4 => x"12", 5 => x"51", 6 => x"20", 7 => x"30", 8 => x"49", 9 => x"88", others => x"00"); 
constant weight24 : rom_type := ( 0 => x"00", 1 => x"25", 2 => x"58", 3 => x"56", 4 => x"95", 5 => x"92", 6 => x"69", 7 => x"89", 8 => x"76", 9 => x"21", others => x"00"); 
constant weight25 : rom_type := ( 0 => x"00", 1 => x"44", 2 => x"99", 3 => x"99", 4 => x"71", 5 => x"46", 6 => x"39", 7 => x"88", 8 => x"96", 9 => x"19", others => x"00"); 
constant weight26 : rom_type := ( 0 => x"00", 1 => x"69", 2 => x"15", 3 => x"67", 4 => x"53", 5 => x"52", 6 => x"84", 7 => x"30", 8 => x"41", 9 => x"79", others => x"00"); 
constant weight27 : rom_type := ( 0 => x"00", 1 => x"52", 2 => x"91", 3 => x"30", 4 => x"23", 5 => x"11", 6 => x"36", 7 => x"98", 8 => x"32", 9 => x"46", others => x"00"); 
constant weight28 : rom_type := ( 0 => x"00", 1 => x"11", 2 => x"99", 3 => x"67", 4 => x"28", 5 => x"71", 6 => x"99", 7 => x"17", 8 => x"97", 9 => x"56", others => x"00"); 
constant weight29 : rom_type := ( 0 => x"00", 1 => x"77", 2 => x"25", 3 => x"78", 4 => x"63", 5 => x"50", 6 => x"32", 7 => x"33", 8 => x"59", 9 => x"71", others => x"00"); 
constant weight30 : rom_type := ( 0 => x"00", 1 => x"47", 2 => x"66", 3 => x"48", 4 => x"12", 5 => x"84", 6 => x"36", 7 => x"70", 8 => x"31", 9 => x"61", others => x"00"); 
constant weight31 : rom_type := ( 0 => x"00", 1 => x"75", 2 => x"84", 3 => x"84", 4 => x"14", 5 => x"14", 6 => x"62", 7 => x"20", 8 => x"70", 9 => x"94", others => x"00"); 
constant weight32 : rom_type := ( 0 => x"00", 1 => x"99", 2 => x"14", 3 => x"18", 4 => x"81", 5 => x"56", 6 => x"51", 7 => x"23", 8 => x"58", 9 => x"76", others => x"00"); 
constant weight33 : rom_type := ( 0 => x"00", 1 => x"44", 2 => x"77", 3 => x"26", 4 => x"24", 5 => x"50", 6 => x"66", 7 => x"26", 8 => x"36", 9 => x"88", others => x"00"); 
constant weight34 : rom_type := ( 0 => x"00", 1 => x"76", 2 => x"46", 3 => x"82", 4 => x"49", 5 => x"33", 6 => x"98", 7 => x"90", 8 => x"92", 9 => x"16", others => x"00"); 
constant weight35 : rom_type := ( 0 => x"00", 1 => x"31", 2 => x"30", 3 => x"59", 4 => x"30", 5 => x"68", 6 => x"56", 7 => x"70", 8 => x"42", 9 => x"34", others => x"00"); 
constant weight36 : rom_type := ( 0 => x"00", 1 => x"74", 2 => x"90", 3 => x"26", 4 => x"34", 5 => x"85", 6 => x"41", 7 => x"80", 8 => x"50", 9 => x"70", others => x"00"); 
constant weight37 : rom_type := ( 0 => x"00", 1 => x"69", 2 => x"57", 3 => x"57", 4 => x"60", 5 => x"78", 6 => x"62", 7 => x"11", 8 => x"29", 9 => x"36", others => x"00"); 
constant weight38 : rom_type := ( 0 => x"00", 1 => x"40", 2 => x"76", 3 => x"68", 4 => x"54", 5 => x"46", 6 => x"11", 7 => x"24", 8 => x"21", 9 => x"21", others => x"00"); 
constant weight39 : rom_type := ( 0 => x"00", 1 => x"98", 2 => x"58", 3 => x"54", 4 => x"75", 5 => x"93", 6 => x"45", 7 => x"71", 8 => x"82", 9 => x"24", others => x"00"); 
constant weight40 : rom_type := ( 0 => x"00", 1 => x"20", 2 => x"77", 3 => x"26", 4 => x"37", 5 => x"84", 6 => x"98", 7 => x"20", 8 => x"78", 9 => x"43", others => x"00"); 
constant weight41 : rom_type := ( 0 => x"00", 1 => x"64", 2 => x"45", 3 => x"40", 4 => x"31", 5 => x"26", 6 => x"35", 7 => x"74", 8 => x"98", 9 => x"32", others => x"00"); 
constant weight42 : rom_type := ( 0 => x"00", 1 => x"93", 2 => x"63", 3 => x"29", 4 => x"58", 5 => x"30", 6 => x"32", 7 => x"58", 8 => x"47", 9 => x"43", others => x"00"); 
constant weight43 : rom_type := ( 0 => x"00", 1 => x"47", 2 => x"89", 3 => x"14", 4 => x"50", 5 => x"11", 6 => x"65", 7 => x"87", 8 => x"73", 9 => x"23", others => x"00"); 
constant weight44 : rom_type := ( 0 => x"00", 1 => x"69", 2 => x"86", 3 => x"67", 4 => x"41", 5 => x"68", 6 => x"33", 7 => x"92", 8 => x"24", 9 => x"70", others => x"00"); 
constant weight45 : rom_type := ( 0 => x"00", 1 => x"98", 2 => x"95", 3 => x"94", 4 => x"47", 5 => x"67", 6 => x"35", 7 => x"72", 8 => x"19", 9 => x"62", others => x"00"); 
constant weight46 : rom_type := ( 0 => x"00", 1 => x"80", 2 => x"76", 3 => x"15", 4 => x"96", 5 => x"79", 6 => x"35", 7 => x"89", 8 => x"93", 9 => x"29", others => x"00"); 
constant weight47 : rom_type := ( 0 => x"00", 1 => x"49", 2 => x"54", 3 => x"49", 4 => x"37", 5 => x"57", 6 => x"76", 7 => x"51", 8 => x"75", 9 => x"63", others => x"00"); 
constant weight48 : rom_type := ( 0 => x"00", 1 => x"33", 2 => x"56", 3 => x"13", 4 => x"95", 5 => x"90", 6 => x"99", 7 => x"51", 8 => x"22", 9 => x"30", others => x"00"); 
constant weight49 : rom_type := ( 0 => x"00", 1 => x"29", 2 => x"66", 3 => x"72", 4 => x"60", 5 => x"77", 6 => x"83", 7 => x"36", 8 => x"99", 9 => x"58", others => x"00"); 
constant weight50 : rom_type := ( 0 => x"00", 1 => x"72", 2 => x"62", 3 => x"83", 4 => x"77", 5 => x"84", 6 => x"81", 7 => x"13", 8 => x"90", 9 => x"63", others => x"00"); 
constant weight51 : rom_type := ( 0 => x"00", 1 => x"52", 2 => x"74", 3 => x"40", 4 => x"72", 5 => x"86", 6 => x"64", 7 => x"44", 8 => x"63", 9 => x"93", others => x"00"); 
constant weight52 : rom_type := ( 0 => x"00", 1 => x"97", 2 => x"64", 3 => x"95", 4 => x"40", 5 => x"80", 6 => x"75", 7 => x"44", 8 => x"87", 9 => x"37", others => x"00"); 
constant weight53 : rom_type := ( 0 => x"00", 1 => x"39", 2 => x"85", 3 => x"15", 4 => x"19", 5 => x"99", 6 => x"72", 7 => x"92", 8 => x"89", 9 => x"23", others => x"00"); 
constant weight54 : rom_type := ( 0 => x"00", 1 => x"69", 2 => x"81", 3 => x"22", 4 => x"89", 5 => x"16", 6 => x"80", 7 => x"50", 8 => x"75", 9 => x"35", others => x"00"); 
constant weight55 : rom_type := ( 0 => x"00", 1 => x"96", 2 => x"77", 3 => x"69", 4 => x"57", 5 => x"90", 6 => x"26", 7 => x"54", 8 => x"60", 9 => x"15", others => x"00"); 
constant weight56 : rom_type := ( 0 => x"00", 1 => x"19", 2 => x"87", 3 => x"38", 4 => x"53", 5 => x"82", 6 => x"77", 7 => x"44", 8 => x"86", 9 => x"67", others => x"00"); 
constant weight57 : rom_type := ( 0 => x"00", 1 => x"61", 2 => x"95", 3 => x"32", 4 => x"59", 5 => x"68", 6 => x"71", 7 => x"93", 8 => x"24", 9 => x"35", others => x"00"); 
constant weight58 : rom_type := ( 0 => x"00", 1 => x"88", 2 => x"88", 3 => x"98", 4 => x"96", 5 => x"13", 6 => x"52", 7 => x"23", 8 => x"62", 9 => x"67", others => x"00"); 
constant weight59 : rom_type := ( 0 => x"00", 1 => x"80", 2 => x"20", 3 => x"80", 4 => x"34", 5 => x"83", 6 => x"77", 7 => x"76", 8 => x"17", 9 => x"87", others => x"00"); 
constant weight60 : rom_type := ( 0 => x"00", 1 => x"26", 2 => x"69", 3 => x"38", 4 => x"61", 5 => x"34", 6 => x"18", 7 => x"39", 8 => x"10", 9 => x"64", others => x"00"); 
constant weight61 : rom_type := ( 0 => x"00", 1 => x"25", 2 => x"75", 3 => x"60", 4 => x"85", 5 => x"16", 6 => x"81", 7 => x"92", 8 => x"70", 9 => x"47", others => x"00"); 
constant weight62 : rom_type := ( 0 => x"00", 1 => x"11", 2 => x"35", 3 => x"82", 4 => x"83", 5 => x"99", 6 => x"84", 7 => x"75", 8 => x"77", 9 => x"42", others => x"00"); 
constant weight63 : rom_type := ( 0 => x"00", 1 => x"22", 2 => x"47", 3 => x"53", 4 => x"71", 5 => x"19", 6 => x"83", 7 => x"43", 8 => x"53", 9 => x"81", others => x"00"); 
constant weight64 : rom_type := ( 0 => x"00", 1 => x"59", 2 => x"76", 3 => x"96", 4 => x"66", 5 => x"48", 6 => x"67", 7 => x"68", 8 => x"74", 9 => x"72", others => x"00"); 

constant weight65 : rom_type := ( 0 => x"00", 1 => x"9b", 2 => x"6e", 3 => x"6d", 4 => x"f4", 5 => x"09", 6 => x"cf", 7 => x"89", 8 => x"46", 9 => x"c0", others => x"00"); 
constant weight66 : rom_type := ( 0 => x"00", 1 => x"70", 2 => x"db", 3 => x"46", 4 => x"83", 5 => x"49", 6 => x"ed", 7 => x"96", 8 => x"11", 9 => x"42", others => x"00"); 
constant weight67 : rom_type := ( 0 => x"00", 1 => x"c4", 2 => x"80", 3 => x"19", 4 => x"26", 5 => x"70", 6 => x"4a", 7 => x"29", 8 => x"32", 9 => x"eb", others => x"00"); 
constant weight68 : rom_type := ( 0 => x"00", 1 => x"6d", 2 => x"2a", 3 => x"4a", 4 => x"87", 5 => x"d4", 6 => x"8e", 7 => x"b4", 8 => x"15", 9 => x"84", others => x"00"); 
constant weight69 : rom_type := ( 0 => x"00", 1 => x"0e", 2 => x"a9", 3 => x"38", 4 => x"69", 5 => x"69", 6 => x"24", 7 => x"83", 8 => x"9e", 9 => x"36", others => x"00"); 
constant weight70 : rom_type := ( 0 => x"00", 1 => x"44", 2 => x"6d", 3 => x"d1", 4 => x"9a", 5 => x"0d", 6 => x"8f", 7 => x"c1", 8 => x"63", 9 => x"6b", others => x"00"); 
constant weight71 : rom_type := ( 0 => x"00", 1 => x"24", 2 => x"fe", 3 => x"ba", 4 => x"99", 5 => x"91", 6 => x"22", 7 => x"0f", 8 => x"78", 9 => x"a4", others => x"00"); 
constant weight72 : rom_type := ( 0 => x"00", 1 => x"01", 2 => x"19", 3 => x"81", 4 => x"ca", 5 => x"14", 6 => x"1d", 7 => x"82", 8 => x"15", 9 => x"5c", others => x"00"); 
constant weight73 : rom_type := ( 0 => x"00", 1 => x"05", 2 => x"e7", 3 => x"64", 4 => x"f6", 5 => x"16", 6 => x"87", 7 => x"f2", 8 => x"18", 9 => x"ff", others => x"00"); 
constant weight74 : rom_type := ( 0 => x"00", 1 => x"0e", 2 => x"19", 3 => x"93", 4 => x"d4", 5 => x"65", 6 => x"17", 7 => x"65", 8 => x"97", 9 => x"99", others => x"00"); 
constant weight75 : rom_type := ( 0 => x"00", 1 => x"aa", 2 => x"b8", 3 => x"67", 4 => x"5a", 5 => x"34", 6 => x"49", 7 => x"a3", 8 => x"24", 9 => x"c4", others => x"00"); 
constant weight76 : rom_type := ( 0 => x"00", 1 => x"a0", 2 => x"64", 3 => x"58", 4 => x"73", 5 => x"57", 6 => x"a1", 7 => x"f5", 8 => x"74", 9 => x"e1", others => x"00"); 
constant weight77 : rom_type := ( 0 => x"00", 1 => x"40", 2 => x"dd", 3 => x"60", 4 => x"78", 5 => x"5c", 6 => x"6b", 7 => x"9b", 8 => x"20", 9 => x"7b", others => x"00"); 
constant weight78 : rom_type := ( 0 => x"00", 1 => x"e3", 2 => x"32", 3 => x"61", 4 => x"f5", 5 => x"c5", 6 => x"54", 7 => x"93", 8 => x"dc", 9 => x"05", others => x"00"); 
constant weight79 : rom_type := ( 0 => x"00", 1 => x"c4", 2 => x"4c", 3 => x"e3", 4 => x"37", 5 => x"f3", 6 => x"ff", 7 => x"5e", 8 => x"9d", 9 => x"72", others => x"00"); 
constant weight80 : rom_type := ( 0 => x"00", 1 => x"91", 2 => x"37", 3 => x"d0", 4 => x"91", 5 => x"8f", 6 => x"99", 7 => x"a2", 8 => x"13", 9 => x"ff", others => x"00"); 
constant weight81 : rom_type := ( 0 => x"00", 1 => x"f8", 2 => x"97", 3 => x"c6", 4 => x"ad", 5 => x"29", 6 => x"71", 7 => x"04", 8 => x"1f", 9 => x"7e", others => x"00"); 
constant weight82 : rom_type := ( 0 => x"00", 1 => x"2d", 2 => x"cb", 3 => x"1f", 4 => x"1d", 5 => x"a1", 6 => x"83", 7 => x"13", 8 => x"c4", 9 => x"3c", others => x"00"); 
constant weight83 : rom_type := ( 0 => x"00", 1 => x"8c", 2 => x"f0", 3 => x"04", 4 => x"23", 5 => x"dd", 6 => x"84", 7 => x"90", 8 => x"8d", 9 => x"a1", others => x"00"); 
constant weight84 : rom_type := ( 0 => x"00", 1 => x"3b", 2 => x"87", 3 => x"fb", 4 => x"89", 5 => x"95", 6 => x"47", 7 => x"0d", 8 => x"8a", 9 => x"c2", others => x"00"); 
constant weight85 : rom_type := ( 0 => x"00", 1 => x"e7", 2 => x"5e", 3 => x"8e", 4 => x"f0", 5 => x"f9", 6 => x"5f", 7 => x"26", 8 => x"c2", 9 => x"47", others => x"00"); 
constant weight86 : rom_type := ( 0 => x"00", 1 => x"f1", 2 => x"ec", 3 => x"76", 4 => x"41", 5 => x"d4", 6 => x"5c", 7 => x"22", 8 => x"b7", 9 => x"47", others => x"00"); 
constant weight87 : rom_type := ( 0 => x"00", 1 => x"ab", 2 => x"33", 3 => x"8c", 4 => x"8d", 5 => x"da", 6 => x"1d", 7 => x"98", 8 => x"4a", 9 => x"d2", others => x"00"); 
constant weight88 : rom_type := ( 0 => x"00", 1 => x"03", 2 => x"90", 3 => x"69", 4 => x"1f", 5 => x"ca", 6 => x"53", 7 => x"f0", 8 => x"ef", 9 => x"61", others => x"00"); 
constant weight89 : rom_type := ( 0 => x"00", 1 => x"41", 2 => x"b4", 3 => x"19", 4 => x"bf", 5 => x"b5", 6 => x"a2", 7 => x"5b", 8 => x"d0", 9 => x"6d", others => x"00"); 
constant weight90 : rom_type := ( 0 => x"00", 1 => x"dc", 2 => x"da", 3 => x"81", 4 => x"74", 5 => x"03", 6 => x"38", 7 => x"c9", 8 => x"2a", 9 => x"44", others => x"00"); 
constant weight91 : rom_type := ( 0 => x"00", 1 => x"c5", 2 => x"89", 3 => x"61", 4 => x"b0", 5 => x"a3", 6 => x"ad", 7 => x"ee", 8 => x"7a", 9 => x"81", others => x"00"); 
constant weight92 : rom_type := ( 0 => x"00", 1 => x"ab", 2 => x"b3", 3 => x"e6", 4 => x"59", 5 => x"d8", 6 => x"05", 7 => x"16", 8 => x"ef", 9 => x"a7", others => x"00"); 
constant weight93 : rom_type := ( 0 => x"00", 1 => x"3e", 2 => x"89", 3 => x"bf", 4 => x"7d", 5 => x"b5", 6 => x"7a", 7 => x"0a", 8 => x"37", 9 => x"37", others => x"00"); 
constant weight94 : rom_type := ( 0 => x"00", 1 => x"47", 2 => x"ba", 3 => x"6e", 4 => x"a1", 5 => x"18", 6 => x"a0", 7 => x"79", 8 => x"b3", 9 => x"cb", others => x"00"); 
constant weight95 : rom_type := ( 0 => x"00", 1 => x"0c", 2 => x"3b", 3 => x"aa", 4 => x"6b", 5 => x"d3", 6 => x"eb", 7 => x"c9", 8 => x"51", 9 => x"2a", others => x"00"); 
constant weight96 : rom_type := ( 0 => x"00", 1 => x"b2", 2 => x"2f", 3 => x"a8", 4 => x"fa", 5 => x"dd", 6 => x"40", 7 => x"c0", 8 => x"f1", 9 => x"2c", others => x"00"); 
constant weight97 : rom_type := ( 0 => x"00", 1 => x"dc", 2 => x"f5", 3 => x"84", 4 => x"68", 5 => x"59", 6 => x"1d", 7 => x"8d", 8 => x"9f", 9 => x"66", others => x"00"); 
constant weight98 : rom_type := ( 0 => x"00", 1 => x"78", 2 => x"76", 3 => x"a0", 4 => x"2b", 5 => x"16", 6 => x"6f", 7 => x"ae", 8 => x"58", 9 => x"12", others => x"00"); 
constant weight99 : rom_type := ( 0 => x"00", 1 => x"e5", 2 => x"0c", 3 => x"ac", 4 => x"c1", 5 => x"7e", 6 => x"55", 7 => x"80", 8 => x"e5", 9 => x"48", others => x"00"); 
constant weight100: rom_type := ( 0 => x"00", 1 => x"55", 2 => x"55", 3 => x"28", 4 => x"2e", 5 => x"65", 6 => x"05", 7 => x"0d", 8 => x"3d", 9 => x"a8", others => x"00"); 
constant weight101: rom_type := ( 0 => x"00", 1 => x"25", 2 => x"2e", 3 => x"ba", 4 => x"c5", 5 => x"53", 6 => x"a8", 7 => x"d3", 8 => x"64", 9 => x"13", others => x"00"); 
constant weight102: rom_type := ( 0 => x"00", 1 => x"2b", 2 => x"78", 3 => x"fe", 4 => x"27", 5 => x"57", 6 => x"32", 7 => x"41", 8 => x"7a", 9 => x"20", others => x"00"); 
constant weight103: rom_type := ( 0 => x"00", 1 => x"01", 2 => x"8f", 3 => x"9d", 4 => x"ba", 5 => x"a2", 6 => x"29", 7 => x"db", 8 => x"47", 9 => x"32", others => x"00"); 
constant weight104: rom_type := ( 0 => x"00", 1 => x"31", 2 => x"a7", 3 => x"89", 4 => x"07", 5 => x"d0", 6 => x"a6", 7 => x"aa", 8 => x"60", 9 => x"85", others => x"00"); 
constant weight105: rom_type := ( 0 => x"00", 1 => x"5f", 2 => x"48", 3 => x"8a", 4 => x"ce", 5 => x"df", 6 => x"fe", 7 => x"42", 8 => x"77", 9 => x"aa", others => x"00"); 
constant weight106: rom_type := ( 0 => x"00", 1 => x"ff", 2 => x"27", 3 => x"75", 4 => x"fc", 5 => x"af", 6 => x"8d", 7 => x"a5", 8 => x"da", 9 => x"20", others => x"00"); 
constant weight107: rom_type := ( 0 => x"00", 1 => x"0a", 2 => x"fd", 3 => x"6e", 4 => x"20", 5 => x"fc", 6 => x"bd", 7 => x"d0", 8 => x"b1", 9 => x"03", others => x"00"); 
constant weight108: rom_type := ( 0 => x"00", 1 => x"a8", 2 => x"d3", 3 => x"ee", 4 => x"dc", 5 => x"75", 6 => x"87", 7 => x"cf", 8 => x"11", 9 => x"bd", others => x"00"); 
constant weight109: rom_type := ( 0 => x"00", 1 => x"c7", 2 => x"04", 3 => x"33", 4 => x"60", 5 => x"27", 6 => x"41", 7 => x"df", 8 => x"ec", 9 => x"fb", others => x"00"); 
constant weight110: rom_type := ( 0 => x"00", 1 => x"02", 2 => x"d4", 3 => x"32", 4 => x"f5", 5 => x"7f", 6 => x"39", 7 => x"e3", 8 => x"3b", 9 => x"b2", others => x"00"); 
constant weight111: rom_type := ( 0 => x"00", 1 => x"20", 2 => x"55", 3 => x"ce", 4 => x"6f", 5 => x"26", 6 => x"67", 7 => x"35", 8 => x"05", 9 => x"c7", others => x"00"); 
constant weight112: rom_type := ( 0 => x"00", 1 => x"44", 2 => x"6a", 3 => x"37", 4 => x"9f", 5 => x"84", 6 => x"91", 7 => x"57", 8 => x"5d", 9 => x"67", others => x"00"); 
constant weight113: rom_type := ( 0 => x"00", 1 => x"87", 2 => x"27", 3 => x"8a", 4 => x"1e", 5 => x"a2", 6 => x"2d", 7 => x"b0", 8 => x"87", 9 => x"e5", others => x"00"); 
constant weight114: rom_type := ( 0 => x"00", 1 => x"06", 2 => x"d5", 3 => x"3f", 4 => x"aa", 5 => x"8b", 6 => x"6f", 7 => x"5f", 8 => x"7e", 9 => x"6b", others => x"00"); 
constant weight115: rom_type := ( 0 => x"00", 1 => x"49", 2 => x"e3", 3 => x"eb", 4 => x"d2", 5 => x"bb", 6 => x"d7", 7 => x"2c", 8 => x"de", 9 => x"e3", others => x"00"); 
constant weight116: rom_type := ( 0 => x"00", 1 => x"6f", 2 => x"79", 3 => x"70", 4 => x"b6", 5 => x"8b", 6 => x"b9", 7 => x"43", 8 => x"2c", 9 => x"93", others => x"00"); 
constant weight117: rom_type := ( 0 => x"00", 1 => x"56", 2 => x"9d", 3 => x"6d", 4 => x"03", 5 => x"ad", 6 => x"bd", 7 => x"8a", 8 => x"1b", 9 => x"f6", others => x"00"); 
constant weight118: rom_type := ( 0 => x"00", 1 => x"b5", 2 => x"b6", 3 => x"7e", 4 => x"1b", 5 => x"93", 6 => x"8a", 7 => x"58", 8 => x"87", 9 => x"7b", others => x"00"); 
constant weight119: rom_type := ( 0 => x"00", 1 => x"7d", 2 => x"45", 3 => x"40", 4 => x"58", 5 => x"16", 6 => x"61", 7 => x"68", 8 => x"3d", 9 => x"4a", others => x"00"); 
constant weight120: rom_type := ( 0 => x"00", 1 => x"2e", 2 => x"2f", 3 => x"71", 4 => x"37", 5 => x"5b", 6 => x"87", 7 => x"f5", 8 => x"d4", 9 => x"75", others => x"00"); 
constant weight121: rom_type := ( 0 => x"00", 1 => x"6f", 2 => x"2e", 3 => x"5e", 4 => x"db", 5 => x"5d", 6 => x"ad", 7 => x"9e", 8 => x"aa", 9 => x"a3", others => x"00"); 
constant weight122: rom_type := ( 0 => x"00", 1 => x"c8", 2 => x"61", 3 => x"ff", 4 => x"da", 5 => x"35", 6 => x"72", 7 => x"17", 8 => x"38", 9 => x"0d", others => x"00"); 
constant weight123: rom_type := ( 0 => x"00", 1 => x"8e", 2 => x"9e", 3 => x"36", 4 => x"a1", 5 => x"42", 6 => x"c4", 7 => x"2a", 8 => x"17", 9 => x"86", others => x"00"); 
constant weight124: rom_type := ( 0 => x"00", 1 => x"41", 2 => x"69", 3 => x"a3", 4 => x"12", 5 => x"cf", 6 => x"26", 7 => x"49", 8 => x"72", 9 => x"7a", others => x"00"); 
constant weight125: rom_type := ( 0 => x"00", 1 => x"83", 2 => x"d3", 3 => x"c6", 4 => x"a2", 5 => x"28", 6 => x"0c", 7 => x"09", 8 => x"1b", 9 => x"21", others => x"00"); 
constant weight126: rom_type := ( 0 => x"00", 1 => x"be", 2 => x"90", 3 => x"7e", 4 => x"30", 5 => x"9c", 6 => x"89", 7 => x"b2", 8 => x"f7", 9 => x"92", others => x"00"); 
constant weight127: rom_type := ( 0 => x"00", 1 => x"25", 2 => x"ad", 3 => x"c3", 4 => x"0a", 5 => x"81", 6 => x"06", 7 => x"eb", 8 => x"13", 9 => x"7c", others => x"00"); 
constant weight128: rom_type := ( 0 => x"00", 1 => x"bd", 2 => x"11", 3 => x"ff", 4 => x"96", 5 => x"bb", 6 => x"2e", 7 => x"c3", 8 => x"19", 9 => x"66", others => x"00"); 

-- weight init 

signal  w01_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w02_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w03_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w04_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w05_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w06_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w07_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w08_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w09_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w10_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w11_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w12_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w13_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w14_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w15_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w16_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w17_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w18_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w19_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w20_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w21_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w22_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w23_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w24_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w25_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w26_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w27_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w28_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w29_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w30_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w31_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w32_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w33_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w34_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w35_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w36_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w37_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w38_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w39_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w40_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w41_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w42_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w43_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w44_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w45_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w46_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w47_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w48_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w49_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w50_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w51_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w52_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w53_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w54_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w55_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w56_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w57_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w58_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w59_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w60_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w61_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w62_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w63_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w64_in    : std_logic_vector(CL_w_width-1 downto 0);

signal  w65_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w66_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w67_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w68_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w69_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w70_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w71_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w72_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w73_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w74_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w75_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w76_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w77_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w78_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w79_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w80_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w81_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w82_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w83_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w84_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w85_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w86_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w87_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w88_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w89_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w90_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w91_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w92_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w93_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w94_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w95_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w96_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w97_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w98_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w99_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w100_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w101_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w102_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w103_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w104_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w105_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w106_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w107_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w108_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w109_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w110_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w111_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w112_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w113_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w114_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w115_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w116_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w117_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w118_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w119_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w120_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w121_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w122_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w123_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w124_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w125_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w126_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w127_in    : std_logic_vector(CL_w_width-1 downto 0);
signal  w128_in    : std_logic_vector(CL_w_width-1 downto 0);

signal  w_num       : std_logic_vector(  3 downto 0);
signal  w_en        : std_logic;
signal  w_count     : std_logic_vector(  3 downto 0);
signal  w_count_en  : std_logic;
signal  w_count_en2 : std_logic;

-- conv layer
constant CL_W       : integer := N+CL_w_width+4; -- output data width
constant CL_SR      : integer := 0; -- data shift right before output
signal  cl_en_out, cl_sof_out: std_logic;
signal  d01_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d02_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d03_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d04_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d05_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d06_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d07_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d08_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d09_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d10_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d11_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d12_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d13_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d14_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d15_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d16_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d17_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d18_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d19_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d20_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d21_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d22_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d23_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d24_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d25_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d26_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d27_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d28_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d29_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d30_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d31_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d32_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d33_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d34_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d35_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d36_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d37_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d38_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d39_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d40_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d41_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d42_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d43_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d44_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d45_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d46_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d47_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d48_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d49_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d50_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d51_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d52_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d53_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d54_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d55_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d56_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d57_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d58_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d59_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d60_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d61_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d62_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d63_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d64_out1       : std_logic_vector (CL_W-1 downto 0);

signal  d65_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d66_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d67_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d68_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d69_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d70_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d71_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d72_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d73_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d74_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d75_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d76_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d77_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d78_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d79_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d80_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d81_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d82_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d83_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d84_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d85_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d86_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d87_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d88_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d89_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d90_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d91_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d92_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d93_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d94_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d95_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d96_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d97_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d98_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d99_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d100_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d101_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d102_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d103_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d104_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d105_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d106_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d107_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d108_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d109_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d110_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d111_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d112_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d113_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d114_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d115_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d116_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d117_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d118_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d119_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d120_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d121_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d122_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d123_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d124_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d125_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d126_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d127_out1       : std_logic_vector (CL_W-1 downto 0);
signal  d128_out1       : std_logic_vector (CL_W-1 downto 0);

constant PCA_data_w   : integer := 8; -- PCA data width
signal  d01_out       : std_logic_vector (CL_W-1 downto 0);
signal  d02_out       : std_logic_vector (CL_W-1 downto 0);
signal  d03_out       : std_logic_vector (CL_W-1 downto 0);
signal  d04_out       : std_logic_vector (CL_W-1 downto 0);
signal  d05_out       : std_logic_vector (CL_W-1 downto 0);
signal  d06_out       : std_logic_vector (CL_W-1 downto 0);
signal  d07_out       : std_logic_vector (CL_W-1 downto 0);
signal  d08_out       : std_logic_vector (CL_W-1 downto 0);
signal  d09_out       : std_logic_vector (CL_W-1 downto 0);
signal  d10_out       : std_logic_vector (CL_W-1 downto 0);
signal  d11_out       : std_logic_vector (CL_W-1 downto 0);
signal  d12_out       : std_logic_vector (CL_W-1 downto 0);
signal  d13_out       : std_logic_vector (CL_W-1 downto 0);
signal  d14_out       : std_logic_vector (CL_W-1 downto 0);
signal  d15_out       : std_logic_vector (CL_W-1 downto 0);
signal  d16_out       : std_logic_vector (CL_W-1 downto 0);
signal  d17_out       : std_logic_vector (CL_W-1 downto 0);
signal  d18_out       : std_logic_vector (CL_W-1 downto 0);
signal  d19_out       : std_logic_vector (CL_W-1 downto 0);
signal  d20_out       : std_logic_vector (CL_W-1 downto 0);
signal  d21_out       : std_logic_vector (CL_W-1 downto 0);
signal  d22_out       : std_logic_vector (CL_W-1 downto 0);
signal  d23_out       : std_logic_vector (CL_W-1 downto 0);
signal  d24_out       : std_logic_vector (CL_W-1 downto 0);
signal  d25_out       : std_logic_vector (CL_W-1 downto 0);
signal  d26_out       : std_logic_vector (CL_W-1 downto 0);
signal  d27_out       : std_logic_vector (CL_W-1 downto 0);
signal  d28_out       : std_logic_vector (CL_W-1 downto 0);
signal  d29_out       : std_logic_vector (CL_W-1 downto 0);
signal  d30_out       : std_logic_vector (CL_W-1 downto 0);
signal  d31_out       : std_logic_vector (CL_W-1 downto 0);
signal  d32_out       : std_logic_vector (CL_W-1 downto 0);
signal  d33_out       : std_logic_vector (CL_W-1 downto 0);
signal  d34_out       : std_logic_vector (CL_W-1 downto 0);
signal  d35_out       : std_logic_vector (CL_W-1 downto 0);
signal  d36_out       : std_logic_vector (CL_W-1 downto 0);
signal  d37_out       : std_logic_vector (CL_W-1 downto 0);
signal  d38_out       : std_logic_vector (CL_W-1 downto 0);
signal  d39_out       : std_logic_vector (CL_W-1 downto 0);
signal  d40_out       : std_logic_vector (CL_W-1 downto 0);
signal  d41_out       : std_logic_vector (CL_W-1 downto 0);
signal  d42_out       : std_logic_vector (CL_W-1 downto 0);
signal  d43_out       : std_logic_vector (CL_W-1 downto 0);
signal  d44_out       : std_logic_vector (CL_W-1 downto 0);
signal  d45_out       : std_logic_vector (CL_W-1 downto 0);
signal  d46_out       : std_logic_vector (CL_W-1 downto 0);
signal  d47_out       : std_logic_vector (CL_W-1 downto 0);
signal  d48_out       : std_logic_vector (CL_W-1 downto 0);
signal  d49_out       : std_logic_vector (CL_W-1 downto 0);
signal  d50_out       : std_logic_vector (CL_W-1 downto 0);
signal  d51_out       : std_logic_vector (CL_W-1 downto 0);
signal  d52_out       : std_logic_vector (CL_W-1 downto 0);
signal  d53_out       : std_logic_vector (CL_W-1 downto 0);
signal  d54_out       : std_logic_vector (CL_W-1 downto 0);
signal  d55_out       : std_logic_vector (CL_W-1 downto 0);
signal  d56_out       : std_logic_vector (CL_W-1 downto 0);
signal  d57_out       : std_logic_vector (CL_W-1 downto 0);
signal  d58_out       : std_logic_vector (CL_W-1 downto 0);
signal  d59_out       : std_logic_vector (CL_W-1 downto 0);
signal  d60_out       : std_logic_vector (CL_W-1 downto 0);
signal  d61_out       : std_logic_vector (CL_W-1 downto 0);
signal  d62_out       : std_logic_vector (CL_W-1 downto 0);
signal  d63_out       : std_logic_vector (CL_W-1 downto 0);
signal  d64_out       : std_logic_vector (CL_W-1 downto 0);

signal  d65_out       : std_logic_vector (CL_W-1 downto 0);
signal  d66_out       : std_logic_vector (CL_W-1 downto 0);
signal  d67_out       : std_logic_vector (CL_W-1 downto 0);
signal  d68_out       : std_logic_vector (CL_W-1 downto 0);
signal  d69_out       : std_logic_vector (CL_W-1 downto 0);
signal  d70_out       : std_logic_vector (CL_W-1 downto 0);
signal  d71_out       : std_logic_vector (CL_W-1 downto 0);
signal  d72_out       : std_logic_vector (CL_W-1 downto 0);
signal  d73_out       : std_logic_vector (CL_W-1 downto 0);
signal  d74_out       : std_logic_vector (CL_W-1 downto 0);
signal  d75_out       : std_logic_vector (CL_W-1 downto 0);
signal  d76_out       : std_logic_vector (CL_W-1 downto 0);
signal  d77_out       : std_logic_vector (CL_W-1 downto 0);
signal  d78_out       : std_logic_vector (CL_W-1 downto 0);
signal  d79_out       : std_logic_vector (CL_W-1 downto 0);
signal  d80_out       : std_logic_vector (CL_W-1 downto 0);
signal  d81_out       : std_logic_vector (CL_W-1 downto 0);
signal  d82_out       : std_logic_vector (CL_W-1 downto 0);
signal  d83_out       : std_logic_vector (CL_W-1 downto 0);
signal  d84_out       : std_logic_vector (CL_W-1 downto 0);
signal  d85_out       : std_logic_vector (CL_W-1 downto 0);
signal  d86_out       : std_logic_vector (CL_W-1 downto 0);
signal  d87_out       : std_logic_vector (CL_W-1 downto 0);
signal  d88_out       : std_logic_vector (CL_W-1 downto 0);
signal  d89_out       : std_logic_vector (CL_W-1 downto 0);
signal  d90_out       : std_logic_vector (CL_W-1 downto 0);
signal  d91_out       : std_logic_vector (CL_W-1 downto 0);
signal  d92_out       : std_logic_vector (CL_W-1 downto 0);
signal  d93_out       : std_logic_vector (CL_W-1 downto 0);
signal  d94_out       : std_logic_vector (CL_W-1 downto 0);
signal  d95_out       : std_logic_vector (CL_W-1 downto 0);
signal  d96_out       : std_logic_vector (CL_W-1 downto 0);
signal  d97_out       : std_logic_vector (CL_W-1 downto 0);
signal  d98_out       : std_logic_vector (CL_W-1 downto 0);
signal  d99_out       : std_logic_vector (CL_W-1 downto 0);
signal  d100_out       : std_logic_vector (CL_W-1 downto 0);
signal  d101_out       : std_logic_vector (CL_W-1 downto 0);
signal  d102_out       : std_logic_vector (CL_W-1 downto 0);
signal  d103_out       : std_logic_vector (CL_W-1 downto 0);
signal  d104_out       : std_logic_vector (CL_W-1 downto 0);
signal  d105_out       : std_logic_vector (CL_W-1 downto 0);
signal  d106_out       : std_logic_vector (CL_W-1 downto 0);
signal  d107_out       : std_logic_vector (CL_W-1 downto 0);
signal  d108_out       : std_logic_vector (CL_W-1 downto 0);
signal  d109_out       : std_logic_vector (CL_W-1 downto 0);
signal  d110_out       : std_logic_vector (CL_W-1 downto 0);
signal  d111_out       : std_logic_vector (CL_W-1 downto 0);
signal  d112_out       : std_logic_vector (CL_W-1 downto 0);
signal  d113_out       : std_logic_vector (CL_W-1 downto 0);
signal  d114_out       : std_logic_vector (CL_W-1 downto 0);
signal  d115_out       : std_logic_vector (CL_W-1 downto 0);
signal  d116_out       : std_logic_vector (CL_W-1 downto 0);
signal  d117_out       : std_logic_vector (CL_W-1 downto 0);
signal  d118_out       : std_logic_vector (CL_W-1 downto 0);
signal  d119_out       : std_logic_vector (CL_W-1 downto 0);
signal  d120_out       : std_logic_vector (CL_W-1 downto 0);
signal  d121_out       : std_logic_vector (CL_W-1 downto 0);
signal  d122_out       : std_logic_vector (CL_W-1 downto 0);
signal  d123_out       : std_logic_vector (CL_W-1 downto 0);
signal  d124_out       : std_logic_vector (CL_W-1 downto 0);
signal  d125_out       : std_logic_vector (CL_W-1 downto 0);
signal  d126_out       : std_logic_vector (CL_W-1 downto 0);
signal  d127_out       : std_logic_vector (CL_W-1 downto 0);
signal  d128_out       : std_logic_vector (CL_W-1 downto 0);
-- PCA weights

type pca_mem_type is array ( 0 to 127 ) of std_logic_vector(CL_w_width-1 downto 0 ) ;
signal pca_mem : pca_mem_type;
signal pca_w01,pca_w02,pca_w03,pca_w04,pca_w05,pca_w06,pca_w07,pca_w08,pca_w09,pca_w10,pca_w11,pca_w12,pca_w13,pca_w14,pca_w15,pca_w16 : std_logic_vector (7 downto 0);
signal pca_w17,pca_w18,pca_w19,pca_w20,pca_w21,pca_w22,pca_w23,pca_w24,pca_w25,pca_w26,pca_w27,pca_w28,pca_w29,pca_w30,pca_w31,pca_w32 : std_logic_vector (7 downto 0);
signal pca_w33,pca_w34,pca_w35,pca_w36,pca_w37,pca_w38,pca_w39,pca_w40,pca_w41,pca_w42,pca_w43,pca_w44,pca_w45,pca_w46,pca_w47,pca_w48 : std_logic_vector (7 downto 0);
signal pca_w49,pca_w50,pca_w51,pca_w52,pca_w53,pca_w54,pca_w55,pca_w56,pca_w57,pca_w58,pca_w59,pca_w60,pca_w61,pca_w62,pca_w63,pca_w64 : std_logic_vector (7 downto 0);
signal pca_w65,pca_w66,pca_w67,pca_w68,pca_w69,pca_w70,pca_w71,pca_w72,pca_w73,pca_w74,pca_w75,pca_w76,pca_w77,pca_w78,pca_w79,pca_w80 : std_logic_vector (7 downto 0);
signal pca_w81,pca_w82,pca_w83,pca_w84,pca_w85,pca_w86,pca_w87,pca_w88,pca_w89,pca_w90,pca_w91,pca_w92,pca_w93,pca_w94,pca_w95,pca_w96 : std_logic_vector (7 downto 0);
signal pca_w97,pca_w98,pca_w99,pca_w100, pca_w101,  pca_w102,  pca_w103,  pca_w104,  pca_w105,  pca_w106,  pca_w107,  pca_w108,  pca_w109,  pca_w110,  pca_w111  : std_logic_vector (7 downto 0);
signal pca_w112,  pca_w113,  pca_w114,  pca_w115,  pca_w116,  pca_w117,  pca_w118,  pca_w119,  pca_w120,  pca_w121,  pca_w122,  pca_w123,  pca_w124,  pca_w125,  pca_w126,  pca_w127,  pca_w128 : std_logic_vector (7 downto 0);

type PCArom_type is array ( 0 to 127 ) of std_logic_vector(128*8-1 downto 0 ) ;
constant Pw: --PCAweight64 : 
PCArom_type := 
(  0 => x"64bc1efb896a67a20e171d4f69967628b785fd1b8225ea5cc81832d5c9a9be0c2ae30eb9146aa502dd8587708ff1b753790483cf6733f2182529bc72537085b2969fb178e9ce4d0166e4983c39739d66ea98f6e3a31f9fd44cf261c37fce041c824105477e56eb35886cd73e1e2723e319d09d774fa96afbff7d4ea65f7d9d81", 
   1 => x"987a6d88e79b980037f1d45f6a927370ab11057ae29065b0b2dd3838a92041ea54b73cb2aed4010fec63ecea9cfbc51db016af32240b3d853fd586dd6eabd765a8e01d27e8711e14e1ed6da847fd2e34a3d1fda6eb20ae4134e2a4cfba38c7d01a1a29303f78071c24a0b97412f74e1ab507aecf702c89347d05935ae0221dae", 
   2 => x"8b0e6d137288b3a7837af181bcbb527c26f9ae682e903707e4882a6394983d0bed2621dffe7d93bea8f92d7a166b76cfeb1bf849cbfa99421b296f0bc5d626e2a16820d93c0376db6e44aaa417ef39928eda35467152584800854dbb1bfd7f50ae4eb474a3ee36ed24594df7d5c32501bc2b614b9221bcf0a6aa1ac3cb7c9dee", 
   3 => x"d03e3d48194d1c12406fc5eeb705c9a90b3ec67298a8d725bbfc848d5fd351936696cba1d25dfaef23a29ae45db9a8f498544fbb35459a8121716c0e766704b267f218069765a39d0e15c4ed87b3dceaa76ddde98ca36bee295e02aad1b23852f6e75ba829c8b5dbcc29da3fcae948a9bf95a60619af9662cb007c96ac2e8e6f", 
   4 => x"528d439deed19fdfdd8c2ab90808de3bb27bdda6a0281b766e9d1dc0a7cc74fb13e0bfbe4b13f7bce276bc01e8d616f75fc8919c3d54298db07a1f23a62553aa1824036f7a746be723135be09e1c21526b7f9ed7f5c119332f30e0072dc21402352359d6824285fbcab7d091bd89d26945d5b07334ed0e326808480cb55a917d", 
   5 => x"4411bbc64f5d361f04d1180ded230bbb15aa57f00a5b816c7c7b4600a12c6b8af53efe667c35a2ede68765763ebe888a548a0270c6e1f98dad93677b8344ce62c31fde91b725d305ef4d03511e18f97771646e82c7727386c21486a7b5f313bdb42d1ae14675c0321af8cedb0a303df1c0283f789ec058175a9066f75bee7e56", 
   6 => x"d782cbab61559e0f84a8e67df88b66059cf5ba5547ce1b157559740d4d1ae75d555906136d2b138364c125f233dcf84dcddfbf0064ca7ff496e42fb0903184076c93b6e7d645cb909fa684ebcb0eed2d48efef72141ef7025379414f94874085ff0b69822d38055c1ed7cf0300a3c3f957b182893dcb01e46d097821eeeacf6f", 
   7 => x"5fd8470d2a240f6a08b008e176bd6dd7ffc270f8d7587dee1b19021e32114aaee344063c2f444a92cd7474a58de14f457bd5cbaff480beb497464ac762519e3e1cd8eb7d6dc148d6c39e4346e42a83329866de6aad0aa82fa02b0c9125d79cfe18c80227d0230aa336fa2e5093fdeb64bcaf54a2432d65760fa571f4f06802b3", 
   8 => x"7100de74ba0a1f69cb418887941651e540c1d17bf94d432f6e8a5025263c68097c35e16a6c9f496d0c26ed77dde01dbae951d9e1d35a75a373a458448f1e82b0fddc1aea5d218b8936794219c3960ae7edfb912166ce33033c33914fe975a6fdb3021337664c26c581c651f39541d2fcffb937a0a289fc2cd5cd4b5eab29fd3d", 
   9 => x"d4d0e3b52615cca8266b0a22e0181ade9b93ddd7034e026161fddecfe4149243de01eb1806d739d06bd243976a8c38e43a9c56ade309fdbfe9a14df15a3fcec208780cd0ef9a4d4c490c2507981695770185f45d99c8b59b1f358a2d25b7ea484173438a7999088be89fc76db861206cf0427fab708ce77ebba4c539bf571a2b",
  10 => x"ab1a999238da5c718613bc81a0d0b2c53e446238cf8401e11afe5c213bd5ab334a3bab9e66e0b1b786f367d143e9833b47d629efc078ab9e0632741aca373c37d50af855b57325ff140efe492605bf63c1f0983dc7f48fd84f3fd35eef4499b9e802fc8abe01e26848221da66109d22e6b372a5eec87ebfa66a48737c99b67c6", 
  11 => x"7cd20cdce5be969bcfb2f946d938bb43ff53b2bea3646603842b71c7d38d4660dbe9c761c24f68bfa1ab6d367b85bdc0838e293d935b7c44de7ff3b720038d9871a2e880a6889230d8e46545b513e6e9d7d01d58260c7a321eef640b3e9556c25718dbf8672a69fe9ce7d6564a1816e7dbc9817e64aec93522df2b8a5876904d", 
  12 => x"7ac338f8a773b22b78e5596bc7fd328d99c7092eea96a9bbd3b57fa32b26c12cea0e8d48bed593fe1270caf59d4b1b304dcaf7993733d61231eb01b9232c4a47245ce66ae86ad64736b1c2139115b13ace7d9cbda2d35ac0e82c08a380150e66c60030924c852c3ef843d8d037b08d06813230ed8d97da5b99becc1123220a47", 
  13 => x"b94a3e439c246fa1382074036c57e95dae129d05dbe26ec4a7835e34513b7f164d20680fa2186a5c31c545f469356c0500d67272aa79edca6aba26cd408c3a930d51b168d85b0357230106466d731f75712fcec319123450d0269c0715871b889021f64347a102d62e41198b611c27b8ffb9cecd0fa0b8829ef46f7dbf6d7ed2", 
  14 => x"eab3a050c84bc77b698ea16afce348d9da36957af8572571deea75dd9b4847529861ab99e11b5a6a8d288dec23c16275d3307d0661847c228b0958dbe93b9e5cc5762600e6915419a027331985fe3cddc11e09ed72f5157e7761e0b6cb019366e5aa1bd40829537aaa064b20d2ff0dcbf87daf03847ef5061bb17e6d6e13b507", 
  15 => x"13caf19e29fc9a8243a6f749abad98b5d5d8b85e88175118bc9448c207c098341978f1da83c82c8950fb4dafb8b62d62477ea586994e432a211744b231acc1e65b62705be8e7219be7d2a45737a9d14d6071280e02a89a04efff5307f99ab71abdd601fd544945d56d332205e0887016c0014d66099dd6f695751c4dc4b6d478", 
  16 => x"407643c9319c396158681ceb4b47da1effc12da36f24b86010cbe1a5e1e7e304b9cab1d5a9553a80bce27e57ce306055078a79052d9bdbac91567d7a73c5d23dcd5ba5129dcdc4da9470bdd189e8d18da7891fca82ca44cb7a28d8abb42f83ae6c76cf36a2c87a498076bd44b174d016698d110fd1231911558a5edcbc7a7a1d", 
  17 => x"cb8e284c089316104a17ad702717b83621137171472c14bde0e1843aa30850ee70084d74764b6dd05a7d58a83fe11502404110fbb50b20a679d500e56e4442085dba148e1c16406278b35a929443704de528101c70676aa29c07e844094f3e74f74aa1604a1ddfaf3e51491365c64425880161384d39d052d6e7490f3bf869cb", 
  18 => x"86213ddee81deda67d7d976150c55e296ff5dc2054b646a553bdc176ed609e3a605056a26f0d3e960e1d534d7d661370131ddf8d8753176d0e639882c9402989cb79c8cca80bd97c336b01fb3b71eca02f202a0e928cfb6c48a9336f6218d2f429fe8c024d86856d2b890b2445be9ed79ff275de1c9f2a238a04a6ef0663efca", 
  19 => x"b3b7b9ed04580c13f89a844641eb61979216b10e76415397434ad4dbe4c631ac09b518a54c50b18c540989a9d715a094dc145477907224e465d36fbddf3b4608947830d43b5ee6cdce5c8da58a887921767f6cadc7b646e9aefcad40a64c808e6bac12380ecdf423f05f42716cffe585fe4902c7689fa2811a19ee4bf0b93d7f",
  20 => x"3592c47b7ddcb26018d734082cf81ed07e9632722cc7f59ea2842b5fbaa297cbe1d778aa59796a3d8243d24d7e072243f3af20acbb4960cd5b3c23830413bc60d26aa8e0517e8e6c241f51f32db4e93ceec39014b6110f87077a2adc0fb24d3b902baf6e7626f6190804998d4162a97a62328b1bcff94e6fa2ac13d6630a3072", 
  21 => x"09935d7337cfaa2a596fcc44a391a2bedbb8d83b58c03983dacfb3f49d559717aad6c7e15b523e22516d111be17d4408c2a622856116facd6079cf749c0db54d6d38c335964cb94a9fb47d4a706bf3fadc633c0266e0dbc58737bb3e5ecad1d1f4588a8a33a8d873ee53647671542a11727ef48bd455ecba6a82140d263143cb", 
  22 => x"a23f196e9499d68c88224586f8ec67f121fd73fd17d12fe672821f108613689d263c7c388ac542823390a139a8d96f7f3c19be5381efa1aea49a6e345f5423026adfb4cc1c5cb0e9297a1c5876f835ba3ffe2134dd8f87cd0068c5e53fe4c1819b0da82ae8e5af0a4c701ecca2874e6e3adf384b19bc63e59866783b6f992037", 
  23 => x"bd2f6a6a85133557969ba6dc678be7b2e4142712066bc127182887a23840c8f2c15b650c786052f5013fe38a6ed8e70274c4943dbbafb4767346d6512e3b8aeae408f07ff01c53a31608d21200c8ea881c7f5b14c3a1a256775b15f0df16da04bab4477bf22b484322909096d1d751860aadd5c79a2634669f9aed0bd08300ae", 
  24 => x"45fa0aa376f55f4451a69a3577b55a3b47fbf21503eba32e315c280385803b5801bb32384dc7b61abfaa45f586c30f279a61d97ca18ffcd67dc2573bc928cf9f91064b0ac98782d86d2f37e54413244d5c6067e26255a79522d8166e214c264b0068fbd3e2c4078bbdcf0a7f441afb48e486f57223d0fb84daa48a3ae67474fa", 
  25 => x"48757fa78ef6079b7864ed43450dc0f67ffbddb20ab9542388249cdd5da3a5b672c991e3fb9dec3db104e85a80fd8553a2ac3ad6e020c5616c16f5924abb48d6bee8e5603ee8020ba1dc68bef6fd6e469627f271ff4d119d7b69fa13a734dfa62da66b1ba5da8209731c2098dd8eb4a010892fcc282f3e7f0299241b66deb6cb", 
  26 => x"31d8b965bccb532ce81221e1692c68bd7aacc9d9110f0596ca1fb86f56c789a7155c1f251b0590fc51912a4d8734887274978e6a050d9d2913e7a94b8a8c69ca42c82631b36b2aec37e4b323f2390de3bb687c395bf93bc77ff5533485b50cdcd79b0ea0c68a5e4484bd71ff465fceed33b9530165d2a521023a56c1759cb9b7", 
  27 => x"19402fc218ddb1af8f54e7365c9702595b351d37bcbfb7a9cea4f31c50f22e6a8834c112537f7ccd10bbdc6d8d7c6caa292dfab1b30a4373df9d0378f7260ead1dc2fcebc74229231f5ad188d49a02c6e23f2e8189da2631dc9a7bb3c7212abb16fe93ff85a59f50ecfb3a4d1f69d76b84a324916936418ffd5eaa0c8598e6ff", 
  28 => x"7233386e766d3a7baad3aa0a4b8b7ba8fa255256bd8b3e01510548ae2a3e8c329ee5cac0ff86d36dc45079b43c32da7cb081a63cd79d13f70148fb72785780ef03d454bae21a86da07703f12c18e1b4428e6872a862d2a3e7e369a3a629806cf3da54915c5d3b985a35d010bd7984f49a5d8a7386c131acecea3ed7193b4de78", 
  29 => x"86ffad88296fbfa9d187490674999bee6b41d91f372d707e8da1861d09caee9e589c3f0854adac449a7372c79258418f2d74ef6d0e510a3b0016da2c13eec26c168be62bf2db96a8011f2959bd049dfa179209a25b3a79bd351f20c3b5f9d840ed9b6e416371026f44a43e91a319b3d7f754bbdc8ac3d222da5b5512bef431b3", 
  30 => x"931242718d9409645923def1df56c4b8e32ddee8c05f2e4ac226fe5d1d4767d31a80a407170e2875494fe25068f0bce31ddec8d317faa01b9a59cc36700449014752292f7aa82364765dea1cc8e5f7b2e61669d0b32cd3d977ad15e4ed9267fe19191ed8a06ccf00c18cb27c007d0a1aeaf4c33472ac48eab58bd651b97a4fed", 
  31 => x"ce5467bdb436188fec68d7beb4d5d9a241b78bbc8c24457d7ed4486d65d02ad134931ddd1ab947fb144dac56fdb1c3633697f23ed630a520ae39c9835c91c04dfb54fe98f38f5eeb89bd76ab4a49d625e18bf810aefa7e321a1ede5861ccaaf156193aae710fc486a8253604df3526a52c228e4334300b9541a5258e1d841b57", 
  32 => x"d4af7c18538c40ea4deab1395b537fa588f7ca2c6933b8d4e02dae0f5d8ea1b08a0c0d437da39ca1f352d7b30362d90710da0360c027c298453a1c69700e04a9c944703eadf5fff0c92e0ee4ea505195c431445018d16171c6bdf73d48a3ed3f61c3e50f3ebe94b8811d6056ead52cf0316b9c528d7b43001dce5d258935e0c0", 
  33 => x"148ff70a403deba177ed78198abfc23166d15428e64d0355b7d4fe866962095ac947579ea912d4f754cc9f474222dc74cd976eb84ad9125eb290fcad1ae37cb3f3b6f814f9c937e8b54e6658ee81be4db8f6bb3a5e3cb1d98217301561bea34979288690504b66cfeba869d49cd3b66747e38c3563f0958988c4840ce4b1d5b5", 
  34 => x"5666366804b5de6428bc04dfd2c5202d6153a8218dcbe98a71e622eb3e3b2bfab76abd1334195583fff4ddacde8d8cdfee5f316242ec2ead49785754d41404dad8bbdeb88bd618c71d14dc30a6cf9ad16c382aba6a314b8b7d4d9c023e541c36599a3f4c6b39adc58a2a04a29fe4af95ad72eea5efa1b36958b1ef31a2238b57", 
  35 => x"5db9ef757358e054cba6048e37122b70529cc71cfa647684355abe13b5f13f6a7d9eae6f2df1496ec51060d998a029b5e23619b0d0178d7fe4f85bf2b877c89a6b7b0c99a4b494192a43810f4b265207d756e3c6959d8e38aacbe02120e202d354f9dea138cb699ef1b89217b516b84007db95bfa848c8a4a746277d931226c7", 
  36 => x"0dd8319d995e1e79222463cd3f6e0360a233976edd61994990e81c9a840e167eba92397b1b019eeca9368a49183d29433c810b704ea576c0d0416eed788457268e34be15472eab1860696bc8aeb6844ab17994be4b05a7095a1634a98f681734b09c1ceb3954e3fd17eb42170062f97430ffb069b23ca4c6803beb1df60cfe91", 
  37 => x"82b67f6c63cd53187bfa7ec4ebfecfc7fdd53b4814dde80b99c19141ad4c9abb2595771584820948719e4fab6a013a677971ddf3e3a084cf1cd4a4f5bd923fa1bc45684c9c18a171ff5ef88fd3bffcdf292171ceef89bbbbff5f76879dd13161b16d3d2e065fab8c8e6649221acf5984b160ced7e514d633fa0e255ac392a271", 
  38 => x"e52e8702ab6521d27415b26bf9942e8b6f82185ddc487e621e8f22205cf0bc533d5c0868c405e866b5de49aa84b253c144eafec4214ed7f3020fd422763d223f0b097503745db133f735a51ed254e34a94ebe49ae66aafedbaebf7ba3910806db6c44e0169a6ab1fb4a9a36922366aab900cf0e8ffcbbd5d75e9d51714f6d4f3", 
  39 => x"55de09081c13d06dc4b0c5ec03e89531ca314996a851ece3fc543d8dd9d998169cae07230e5ad2038147e8f4e73d3c95b059586246d02cc292d19faaf409be436db0364954cd88f9f69489793811320b5a4ad1b06b913e00e76541e8bd455efc1a1e41be555fa059b86b5f236f62d08ecf8b58588610a64bfc5549d9951a59e4", 
  40 => x"31c61669dddf50d55ec6d5fedad62e9d19611da38c44e179868ca9541af3330e28d98946a03587ca7f8031cfa0b6b7a61a752ad31cd4214c86bc606d6ca803331585f16e644cfdbff958fc3165b532d30fa178b72803594234d9916eee8f3ef4ce676b13d658ba13644cd964e04cc024d1a1465dbea8291d2834e99861bde419", 
  41 => x"75a44c4551978b2caed19d009ffc0ebfb05df79f2d9447d82abaa399645b2d3a842e1bd3cd5a7e10d6d38f3c0eceaab404c19c1ab6687c97de4a9c8d8e4fc534a2924396ba6a3c85643bf690ae98beee586bc2f20f57ff31b1652936711ee2da95d11c31668229472660bcc849b72ff4248b63a77481cdc22329379c6714781a", 
  42 => x"87e5b37d59ea8cb90d8827fb05c40508635cd943617922992b14e0579078da27b7adbe289b9210ad3b2f644a4573f77b0245c4641e860b378fbe6c87367e141ccbae972c2dd448a519b0bf8dccc222f207f574134794e7af1be845f79df9acddd9fe7fb55b3c38b54cb4131749540f314ccac5a8a16e2608607d38b37b51968c", 
  43 => x"7ddb57b14492f4841cadd5bdcbea2100f9a88eb25f0b30285bc0856923c69538fe736708f3643787542d45d919697172f24ffc921c85a3da34cc75c2d6450d5617f5a80bb3758d1dd38d179a695bd10d30688878b15f1daef7d17b28df687b5c0cab3a9817a5dc8ad9b534626e1f9fd358d4c00c0a7e6ee4cc53848897708501", 
  44 => x"5d01772160fe5a2eb55d03eef15dd8fadad3fb4e1828ab36e1508efdb64f1e81fb614d3a0f1bc1cf8cd707aa763eeb0a344133da78fbbce36fe93a4043cee3107636620e985a7f77f030be3fb97a8b48ccc99126f3b167bd7fbffdd6dca83fcfff848c6e823056a0426490cd5fd6aeeb2e6e08b9b43d176faa0b68957fd12d70", 
  45 => x"e4d41833518273d5c42a3791639fe695d5ce84829215171d08cc77834973fb9a5dd5ac5ef333eb0b99b7bf27d0fc412a2c0bc20276070942606e7fbca8cb0f512ab36d078050801e62cf1358386e8f08c886fd1608d7e1e324d48d31e18c34ec873cceb0ba28e2a1fb37306d7b583fd23c95f17c465a413f63733b1e76e2da3f", 
  46 => x"209912127386b80e2ed6c2d7225d697ca02aaf0e060eeeac57746c5faf958c2ac118c0e24396539e3e11882abaae33f0e906811bf6a0477442e3a4b236011487d2dd33d3741a792702060af788a0d7aa19a3b4b9ceb2f44f97d440d0ea6c698e2e503baa5164781849e9eb3e85ad0f26c8df3aad5b57aa2ecdec9cceb4874fea", 
  47 => x"b258264007054ede6dc9a79cd947e8a244c93b5982c26ba743a4604003d3ac3ddf27a9261c018354286fc936bbdbef85f53d0f0b727eba25987780f2c122a58b113886b6b9992c1e1b20130d5b0dec5fc4c26fe1c4ee9b6d029b60b1c324563438d22deb65e080c8cd8c0bc872b916d8760ee4613276fa77239b3657c73bb607", 
  48 => x"5b2f74e3c5d7cedfd36078568f764144ce656ef3c26999d82206b0bb74987b10a9710b19304a618123e42191f9c63fb5fa8340aaab0af65c5e552dd638afb49d69f780a5395f5ddc349792359ca053f42081a02427af1dc1360b1633d3479d4ad8b2d96d3884c0c51742922346eac8ac29b702440071d38829692e455a33023e", 
  49 => x"8fd8dc48d553888a27dcc1ecdc6a65aa9361e14b3bbd52761e4c1ba47d3b969ed10e3b260e2398bd2837c720932605e99ab173bf47698fd9e1f011a1293f09814af081800c944a50a19b0b60f75962a0771bf0b792164213cd8c7906995f6993c4ebe926064c4101c64794b14fa6b934eb5e44ebed361c5233f5e34ddb6c0709", 
  50 => x"3b941f583e2ef49f09172bdc53e380e6fc6b96bedd29932d730bfa59739384dbc836f32347748ab8bb131d4c3f9bb72a481a7f4487d6f25543dd46d9f21026ab2b8f6e2dd333cd873d45a43838d0adfc06f3d754be6f9747ebd49aa5349d82fb692dc36b95a35d0eb258e043e6e00828817573ab745a730c87dd16b95809451b", 
  51 => x"a9ec322ae057156e62ba4dbe5d5d4adb4a835543c6c7cf9831e7b971e3dc5409bf40596d90d4e92736e8b03431dede184f6dda7eb8d7d8683962cf0d356b2f52c22a9cba667417469a38c77544adf9ad6948bc4af6879b92c83f56f43e5075e48c97c32dbda3fc5ce200df14325e9cc0bc6a8272f7100a7b68193fde2e59b683", 
  52 => x"31d010ca172d3e1f88e37074d71e80975fb7b0fc37a866ca4a629a3a1e811d1a60851dde7909d162cad31523e5e1dabda20c1517019ed1ca7354fa4132f59c3a375af8e93041faa047ae1e33116d6c0a2766fb620254b2d79596f9d7521045357f40d325a2046d86570660b558a4352dad09718b3b12544de1ec4c4db122b6df", 
  53 => x"cfdb072359cd55912014f7e3de2c5bc909f3b76ad23ad0da122c7a2681a3ebd6488985871f400ac893d7e057849510a19d082d47a064eb64a3969e28528b87b9e378ac0d581530d4777c775be9bfb4835f0996fad0259aae27ebbe93002caa5b9420fa2184b3aeab3518994d872de71c90089cda9f62cca6991999b9078a8ba5", 
  54 => x"8672569ed0533692beb951dffe33e9b16d7e712b14e150e1abe8f3c4d7b44f5c544fdfb1a27246c2b0adc0d28e0380d2642645ed73423cfb043f7da5828d4d95e949dac74eee01b09604a061568fad3ca85aed4baa86571ee7cd485017dd4f3bd1da9c4ba1748996484a1c23d8a6b60b634bb5238cee96e043fcdfe40ef4f5aa", 
  55 => x"ad8b6aa916d2e8a5a71644e51194441a1158cc52ac0d1c57eebf69d3ec2679632b5bb2aef236c9778392a1388a61fa52be46a6ed7dc327b83bee16a30316ae3eb44b7819f0329fe52c726cc294790f75bfc87af20352e9c94e6d6b00fe9398015fab2ea3fd99cd561a65bfb9a994b07c13db67091f42535276e893d1a0d52223", 
  56 => x"7657433bcb9a199e7e5af682020564f1590bb49d1d59520c94102f83363ff6dbc19d54325be4f52f273605232b050e1fe0a87e1ff5c13e68df38f400e2d59a6edb86625369db0d2e4029cfe56ee9f3fdee24a190673063d892b849cfa9785ae093f4b312b7554f3be91dd3bf4a0567203fa7cbdfe69fc6f59183351e45e288d6", 
  57 => x"cdf8cffb87798a20bb0fd067d835eece6be0626d0dc7b182971dc4e7510af205cfc31145917f68cc900fd504c60681c0fb970b1e2d470e599efe14f46fc32ecad4d0a1a4256a7175145c5823c5f81d45976ea299b9fabe7807d36cb487dfe7cbaafea5c952cb254d42f718e3613d10b044ded3a35e55009af2a749131dd76245", 
  58 => x"c9271e655e96cbedfd0d4e2e6a854074a0596a3a180af4d3ed98120170fdc902017a1ea87fd021dc15d6dc1f17a22d81921811512655f2ff95ae7b2a12ecfeee6367e01c5452e0580d749ed591a4c474b721b86e9e57d07504cadb9fd8bcee4e7904a121bd479af8429e02cab030efae52144d7983f3deb04b03e6f20ff49b0e", 
  59 => x"68db8e5757f3df72de6b3c0178b65c492d866b652fad05f9230358c8906df08d729a34c78ed7da2e7a3a4d33955589d9eadb477ca0f899e45e00547ace77599420099e16c97442dff1da3c6855ed00343d6a1f0ab69df92b0704c30741c09a68edfb865641e55ebb15821c8347fdd73b408ece65397df3bec97c9c0771ad2e5a", 
  60 => x"5d2178ba0a86a8c9215e4200d3eb80b239bcc5f50d9ba9a19e89ffba00dca8a42510e0bfea03fe686eb9e84a50ac45f347c08f72867239a069eeaaedfc292171d6526bdc0b9ff09d69d9fcdd79bc95f9956874939c1d4d1d89e02d1174e02e363b5dc552d8144fc135fd49c94f8043e46e0b646097d742be9219bb2ccbe62e08", 
  61 => x"7e835c35e9aed6982b573678ec4ec989c50cfb69244d83f20262b3722bd48a12edf83f3896c12cabce132573e88e029d83b1e45475816fb7cd3693fb93710b59f3cb03e5b316ae2f05e8964eb2b1884890011c99c4bc129039c10b95e48d9ceace69b141872b1d64957202e36fb4aa0172724493eedb8524f70e9753dbd5d118", 
  62 => x"58476d76a38a22811b88dcd887d4a4e21863a05660c7a1329c4c8de86ea142a9b8593b3911d11eef3332b92cc6f2639072e7a3cf890cd38e61824bd424cea5d0ad2e185537ba0f7654958dd93942eae26d7e6ace184074a7f3104888675fc00859673d1104b4772593a43f452e413963c3d5b8b57cb134f1d7bbc527bb577ebf", 
  63 => x"436863034df353cf401d32bbbef1a6d1752101a69157010fe3b3e16c6855580b2da52582b52bf0cce2e979b644a44f53a3cc1847864a0d28cc039a4af6812dcd6c25b16a05584cdc3574fc53b29bfa46336234f70a696319cb7540cb9427acb3e8fb02dffe80386a734b317066b3092925d0fb1d38f6b622d0119bcbe7c3b464",
  64 => x"c8d0b58762a6fb273c385cf2b50f141494fc920ad05ca3c443641fdf5ab6c2653c35420237bf46b7485fefda05a3a0f4d52eb4abdecda1385d9a84d94b47c51eb1d01cfb3da1319a43eeecc895aadec611add19a259af46f3e3fd60ed5e801a7e82140dda098914aa083785cdd73110312fb382835d64c335ff73011dc5cf548", 
  65 => x"dcd2c35b49faad1fd07f000ba90a89959ba74f97d10a953672aaa667bc17e8eae7fa3208c55b4c6360019d84bfa39a2b3ec6ae04deda5b9743fd87e4c727552ca7971ab83eb413745b8d0528efa5a71ba033cb257dfa7d6e2d270c533a027911ae4d3d60d5457a7d30583418a857ce84a7562a9b1741cc6097547072ba8dc6f1", 
  66 => x"2b5545668eb84e626347ee5b0ea54b08de48b9a45ee0acbba385a66e765ae26a0841f98e1b01cc2bccc2400d23ad5d06c558847fcbb6080f4eef4317ef55a4516c1f2c971206ecc0733338250a2793818cf587a169fc76d1220c6bc39512ba3aa190a2e21c78c704bba9e05c6ec3601b70f4d34b0634ad27429f42d0d8d952cf", 
  67 => x"3e5267e96eff534ee7a59dc1e00eb892f365e8a9d58466de38fc7f953574070b9d187b41b32dc6e7fd3247054507239dbc3330645beaa1d76e048653f4a86d722d815d9d1a92b90046b3964ff8796bd08a370ca09a5789eb52e42a79f14d93465fe8f87c56beca43308d82d91825c0803c448b2857dbb65f5db22a76ecfac132", 
  68 => x"9ed003216761b668d0c1dc664122bc1940eebd85c9a45ae2730a5580aecefd8c5ba0d68182c8c909120c622514a36dc9ff85d2566195972fd5efd80479c0310206fee5dcc74ee2b664c67d50a400650bb98a90a767c01ab9262f0d324a207a69d60eec3dd570b4ab79d8d246921648512a00c789795a0654effbbf7646f78c8d", 
  69 => x"1c047f948ea9a9b3e1c2bc39d2665b4a92a9e0196b61e1be3121177f375d865cbdf06ee963612b43bac01945e7689ff7c183ee9b6023d1ee6fea583a14a457c5c53f795fccf834038772d5ea2b2260af98f69609ecace421510d3501864fbd8b7b192094b28a5e0d97754ce12d6db214899381427e08ec567f22cea3621d70be", 
  70 => x"343533bc769db73e60a4b66d65f04697c70254f7dd4f7e77464be4518dc481b0aff049b682f0ceb270d1a50a88d51002e35667c2b1de0a8a7092b8a72ff17d87096515c262dc9bd4085a02c88899422b6419f6dcc104b5bd2d3c67f8d17a0cd176874ebc47cd896df7ad72a891ac81e85e0fa90a4835be78004b94cb6fd0398c", 
  71 => x"e5859f83482b83d493f4801bb3d8cd4643785e0c05989539778fe23a35d94978d59be3030b038686f2ed115d666c55c1ea11417fc05a4f758de4e4ac1b28704e494f741bfb165aa62ad40c5a3f8c276fc5a9ef6bcc1288240ffede624911286e668a88b732197bf41a69f75147b9d4ac078af2af001c12a26de791ca0a7bee2e", 
  72 => x"829e466bddb021d62874ddde7afa85aab5ab00672fdcf3e25bcd6b9c7034342efb81d39e81bbd475934fc5a8ddf80a7eaf4af430db16c5c1a9e022192576727dd29c8040e1e56b69880ddf9148433d090b6eb714f6b0abb121280a8146734c6633e12a4d619e70ed17210aab505c7eb15ce9f67e916cbcfb9f09d9bb8ee4690e", 
  73 => x"e5a4705354fed6b876eefcf8f2a6af11ac44f65517078c5da8133ad27e3e5ac2d6637bcd114a56f9fe31d2ca6894edaa4145d5dfacead207d51b51e471534312fb4074450e2e36b28af1aed278725b323f8636d4a9ac352c35d19d90df8fd490ef7b00ccc81ca83b4b698bde0c1e14778a1cc04725b9de407687d3e6d0e69f71",
  74 => x"760f709ab2c9d5378e45aa604ccced6465fa97067179f4d388394324baadb3678ad37870d1c7948edfddc77761724808e5337073e082aafb605963a1badcdc7bd3f0e9e2b23a2bbaa5d068495a862f7fa487652b829adbe5b322eb7c7cbcb431f20d4df5b56b0b4997ac23ec6c130e67354b328d1634f27dda694eefecb410f3", 
  75 => x"d3c5e3c4d7261b14037b49fcccdc37a9fe52fc821f52b81f9675cd682c0984a8d792b6897eb694a88f5a6ba28766aad96996344b53151e25b6239d3592cb15d37c2572b1c5cd744fff894dd676cc60e47d8157854a686e71cd127832e3c16ed6717eb237cf002b48b941edf1d1996ca3fa9fe4ccd5fe995817d4881dba5767c4", 
  76 => x"1dbc7e7d7172fd6e61b91120eac2d76caef81c7b6833d08fd44e1d932d3181aa5b318222b621fb419f3ae8df896003abf80b42f8731300636881ba87fb355860a8544a5cdeac791c5708bc6135d4ba4b362f1de8a77b4135ff2b9825fef13aeab9dab6612d41eaaa705ce0c358f0d3728d568ce63c778d1e23d0bf75e4aa01f9", 
  77 => x"1f800ae2d1d8e6615d3a3e3d45d5621487a0ae173035a77714bdca2657e37dec7b91da31f8b23ed32cf42e97fd60dac16a9f5adf6e328f1ac77cf958c558bd176611954589f97184ef80eb1d119627c3651389d720d2a2e2f959ccf468fe565b51bd6621b29a6f2d204ee262a70d2991694f5a80c45e74edc8a1eb52ba7a2819", 
  78 => x"18f3487096b49506a55c41ba54cf1c6f7ff08095cbe42ef2a360cd27dcfe7e79115adebb7a5bbcc625a859eb322b6e79e24dbd5745896296316d6303d3b458334af11d652476026aa5f7d986401d1ccb228657746c54acc398e962c5c379c20d2467cb391b18d72199cc795ebb6ee73ee50607b9dc8a9d4f2c61c8f627f742b2", 
  79 => x"9cc194ad4c91732414d565b7c7cb5b7eddf820c03dedb380052664ad404caea32c9fadaae3aabc6cf33e80f7b5c2921bce03c22a888b388d747ee0ee618f9aad3d9125bceee80867af5616df32e2fd4ec72eff788cec8e3b309d855ad685b388d9dd78dc9ccaab2285815ef04e9a91595cb60907f44eb24438801d468536e0d8", 
  80 => x"a84b696ef6bbd1e3f0ed31bffd9fb60cfeca9d7766c7937dd4e3c1a1c23a57baf96f6a3256fae6f0cc18d6548147b8ea28cda1cfe68f2d2277d693ea233826a4334ed9f6c7fc2b5ea7b37d6ce375c9028c13243c47653fb8fc8383c5b180d90814e7d498cad09c0a77c46086a272f65d76b4e8081f7c7bec0774ef84714d5016", 
  81 => x"8c083020c337adb02bd0c42d9e6616b43f1034536e2d8ad878dbc2fb3519414e2f96f4d346a541fe81a33cd42478ac11766f354eb827bd39670fa692c46fac9b363ade69b286e498aa1a5157090b3d3bb79ec3e12d0234291a1fde6f070715f17894f3c8247f84f903a6d68b9afb27a0683f7a1dfffc0935fa7e6f3b84339722", 
  82 => x"c67a54d6ed7839617fb7a1c1214e37a6e0342205635a2596a34856271479be09c14319a0420faeff04490089e4b2f4e0b104e959d0f1f4ca4b75861cf666bd2ab782a8734c962a1697a70218047989000c03db4d83775018d6a161473192561a26d85970d88de4a15e60fc207d3dfbfd3b84ccc72502999850876e9426086ca7", 
  83 => x"eea2a2646bbb38dbd3294a65f6c0dffb9315b6314ed3b711a3f1ffb6ad632915181a8679d5d958d8fc64458539c1bef846dae18d949ef1af5e64eb09bbde640cb7ce879a7489933b230e8079d0a4da07263f90c0d9ba5978ad244744192fdbbee21eabab12c38f0242043c2d14359722acb12b5eb2904bc6900ea142cc620700", 
  84 => x"60899132aed77c24c9d3927cd8a2490c55e9b24a2b03f32e7c95f8a6b493ccc89e49d5946f9e932ba4b9c507c5e00da2530e76a003d367225bb25f65b527aebd186d003cc4d3419e429568c6d522771084b611694924d2a01af0a25d3487409b69fe641849a7a1bef644b3b799c478ae2f59793a595959428c5fb40e3fb3fdf1", 
  85 => x"67447a32cab26d1d7be62a319ccd239d92b2b6cd84ed466af7fb33fd4243d8f34cff1a72069e22afee3a842eaf6a17a1490f87549352c278220b8c49825b30a695b89c02480b0ae1ebda08f8d917cfd43e705c4cf1e6f20c82c597f073f910fd29d74a18bd47cbd8d5abf6e27b89ab0c6ead3145f879b6fc7a004e5d5b6926bb", 
  86 => x"b8609733f52947b9b36733970b9fa70b4df15e9b44d55c4c1361c4ed671e20bad45cf18de18c667c737e83fecb8b9d308c73a297d9cab8c49e3404c0ec6ed4560c4392ad6acc2278cfaa123edb1ce21553e35bd8fce966ef65f2a56e8926dc398e138990b1debca3974d7d7b7a1eb0fb7edad92ea041962b7d388ea41196c234", 
  87 => x"72f9a5455e40f910a3dff2464bdce1fab6809ee5816de796fe7c832aa463693291aec6b5e3409bf497ca8f74c23502ea56d7a86ee3a503550c207b42c70f4c6c4c09b3202e494e967d8bc0d63672559e1722905ab5ad4ada0af4b9a8ccd7d043f9b25c95a0d477e3f76b7ceda576e8a5ed380a3ae1121def9986b91673a27362", 
  88 => x"079f83f4db5d5729dd32c0030ec8a1f57cb91b8127893702fd22b54b5bf2004aa2229f3cb395d4a586236ebbcc0965a1426a80798629137e291f055209df236e8e7012078e0087302dbcbb893331b00c8e5ac9fc5caa40a5fb8aa54c61d005258fd785de193642536d942644c3f1d860a20f6da89bf62b85827e699cdc5655a0", 
  89 => x"53d7d822b0c42d8161e2b99bee279bb30db8199c21180701039700cad44f8a5d5b6ad95d9f5ff57c044399037f480174ed510fcdb0b90ade63c30e3cd34c0073203ed9cb8b854aab3ce0439c4f3b9f6abcb4421aec84324a409902d995f5a786b79dd0ea45d0dbc36bba08c0e3470a9108f82b2e31b3618890a5d951e5cd824b", 
  90 => x"5016748de4f12a088af4d02b4ae8691309c7bd9b6e059eed2267f5c1214623f67610e3614ffbfefa25bfabb76ebdb59a7e018a1421a268accda9b625facb162184eba422a63eedbcf162cdaf8885cd3ba15e6eb27f01f96a937c8695780a1ef0d245d4b680846a5d7b8e1ff341532db9b8b3b425ad36b525edb6b4e1d1b56abd", 
  91 => x"53b27adeb6ca1e06622dedc6b4bfdbac23f1c63dc6cb34956b5c8535ba6ba76225b2025519d4160dc2e894d4b242b338a04c7278791b9bdf493ddb7e4445b0d6f9a8d8947c6c0d2b2e41bd09d456b1f4732dd6d80f542f7b8ba9aeb47973ed46dbf3cbbe2798f90b41c00b6a6633fa33ba4e85598128647ef67b9ad90ba90db7", 
  92 => x"d3ae0a67a278cb3d3afd5ef8502db31e7e3ad51253afdd28678f0b4a0dfa0fc87fad57db66a4fb0a5201e3935eaba1f0fc304623711d0e59e8ce17aac4a03b40c029f8f8a43c027a1c13128669f8b20dc89d55629f7b2b049fe694c170831ea1f18b54fd4a0ec34585c89e3b7e759d54ffcbc9dd5f7f3828a929053a4dca3818", 
  93 => x"3c05aebabda22b6ed2f63713c9057cc489362ef318efd7e0232916705ec3e1f684a20fe8f6e2136041aa6c1336bc0547583347a27170f28eded8833bbc389ac34fd059fb89552d6cc3c5cf7b3df82847bf4bce360c20c52ecd9e2ac715b44f558287fb1b4c44424e6815fe32bf2f2ab55223cf309202645265225bfb8e1ddd7e", 
  94 => x"4cc8fc0907e6aa741f609b376243bb1d6155a08edd00d78ebdeb7c106988209640a7a01c118bd06f60ca64dcbc596c7fd14a1cb8b69c8b737e5c9058422ed8457f8b9909006bb166a4c22faef11860512d8e4213b47fe15a74cb11eb838ed9406387bde66a0cd1a6c35b53416c789e3a17c9ffc0df2522e96a0e072d479e1476", 
  95 => x"174e3571d284eac82ab68840dc8d96b3aac43d74d806ea478d1d8ce24be76c2bc1a3da2138312d541f1558bf2b24d0ad81094a6642bf96e254db06eafdf9eb203a5d671170b2edc8c1207d1d508b9d3b97bcf175d31d899ccbfe340c2b3ac501b329bb87f1bf3051543839a337f9ce4dcd4f602afe4e44157ac3a8c3d5c52cae", 
  96 => x"7cb61f071e00e93f2a542a876fdea4ddfdc60f85be7a4c3fe32d76cf726c351e0d47dc32d0c3eb01f0db05c103c04603ce60dc5c33fe4701684175f1c18fb9335803454d99ad2330188431cb2769ed325a8b9f374fcceae5c096a0fbc539591ba30ab7b7e2523e8b620814631338a29d2813d598dd861984e2bf3b179aed22ae", 
  97 => x"941c78eb8cca60af9786ce4ae8d0584107f71b40b83c05ab240f7b5ac8d13caa770b50ae4cf1e2b172473e1d960df3ed04aa522e5e93860e5aa826a0fb5bb0d38dbb003db4f7d12253c6952175237c8dc40676453ad7bd5e1e5e91dc7bb742bf89b788c9ce157c77e3a97345b2d98ef711de1120f386509234826c974c42e70f", 
  98 => x"6b4c3eaab9721e2d489da02d9f10554ef2bbfb615328ffe87e826e63b2b315764476c32a873c42c6b471b085a2483a3e1dd50c8aa3b70ac7cf31e3cafafb572869b413f99ee7a49a34d23dc2618ca0913997c0a700736b0d7b7ed26c1276242923bb18e5dd63bd94f0b42deb95016798a56e2dc0bd48f6191431c10c332dd113", 
  99 => x"d2a6dc9a6c1ee2da21ed42c109ad9c6c40409c58a5c87e4a8ed8411f1e528e932377ed05625260223ab9bec78a914451c9826a233efa729d40fc7f0a5a444168525c1a543ded2a6690c65ecad414f3758f248665d68c93bee8103858d9fbd538f1a5bb750680bcd8abd580fce74cb171e19cb70d24d90c53021eb36e0b9805b3", 
 100 => x"9b806adb44a9515f6a0c85fb5250520e44e6032b3b0419f361032e0e37f61f10e05478bcfd38f2b3e68bed927bec9ecb157aa4dbc72b14d8c001cf88989fbe1e2689e42a68e3bd7101e2ce12932dc0fb9b68b95962eb9054e04fa3388fe23412bb941130f48d039f47ee317ee8c68587e9b00410e3447e3f726e75093ec36c72", 
 101 => x"27b6ecfa06ad5b437e9d74e6536d06e8ac2c950442bd73d09d94be878eb5a5838a4675c3b36b7b9e8aa093701acbcfbdf3ba91f61c2290c295351025a6123997097a3e58c271bd1dbf0994f4c72d798bd32fd105cb6698a50e82043277f6155be4c8e3482f5c0f24acd24e6f6ef767931bedbce50ec68e74b5d45c4a85ad9b17", 
 102 => x"60b378006a65300507385ed6fda42d0cc2330d9b34c6eac34415c6c982cc4113fb63dd32951e245ab91e8b4349a8c73b07c21e6addf1a68f602100f8555b369a591545b284ed172722304128ebe40448b9548cc2551837c05c163e6b43c5b94047cae4bd3ab5439eae1e7fbcdd411534d1b2e93d59372132a09a0cb033f37c58", 
 103 => x"358e40764928a75bce8a6876107f31211158249f081d68edfa9e121c06c0dc42402c8b5092693116304fc69b2ad530e8fe0466704bcda73425fd6803cbe70554c7d2e20ea340713b55654d90570f13dab36232e2debaedd03337d44503db1c4722c684687876920a2bcfdd5cbf7f96ab3e9288e9b4b8c5171d0711c49fdb258d", 
 104 => x"8b4566869080908ddb385b2ef80a4ac769fa275bba2089f00ad3c20910e4a0db780a0db53c690ceda41dca1ed2642eacdbd27b73d45910bec0a6c077ae33dc8c1c6d672603cc06a4aa15bacee26f6dc08a18070af91908543ec560a4dde250e623f825165fbaab821dc011fc8adb99fef0273ccaa35be32c9338484bf50c8713", 
 105 => x"6b184d3cadf5357cd2a5ecfeb2d27b8b319bd4e4c74ab252bcf285dc326e2840aeaf407fd8f50693435c2e96e0784fdbd38d56800c84d45d915f33e2f5c24e781cd1d03b4d8006f36769d5133d656200ac2b7e70f2a21ae135f761db883021d9431196be272f4e9bf2599b1007a2ad8be39f5ebb2f881b45c9d53101b54a031f", 
 106 => x"8cb9f2eba4d71c8cc963d7a975ef1d3aeb3d60b272e2310e81ef33138ccfef670a1f02ab82ef77caa1014d293e395cec1818ded69391774ee8a5098b631eea953e61bc3d86ec03d7559ea544fb6d39ba222e248cb6f2634ba407d49190f68fa4a6c8205dd65198eefd81c042e5989455dfa43744998e9a28edfd91070dbdc3b3", 
 107 => x"7420b73677b344673aac53f30e66cc8fd0628bef81373dd95bc4190413b746a69846afcddcd4ddcd666914fd9c98a69ec6a6eaaf6a01f7b54310e23b3f2acc4d8f95fe0217f711afd75e42e6ce37055e0ccb185ef1b0507f7303aca8dcf14a57b25b42fef2555e2302dedf602ac1691092bf93bf9867097414a0bf8dc498e250", 
 108 => x"8bf4c96b2592c88ff7031cbd77d62ef224ac4e98b28704c8d0b94ffe63720f6ef8a91da56ba8dd43cf8a822459d931b85d8f44d3a3ffe3b046b03028e5a01d85a8b69ee5cde0efeb92a052c3ec7c2f6fa33c25eeacfae1d746644ddb5fef02a764d1a9b0073f55852296bf9b3b9bdad3beee31832a4cda69258f96dbb93ae244", 
 109 => x"6e58e16dd4367a00211a85969c2c0a41c05bf9d6fb38c5311395abc0de06ce116a07719e6f622bd0e192990d8dacb542e89181c3deefedb309c10c44d943dc5fcc5e5c37ca7313cf7799aa09354f5d826769eade545f0c98ad9b87e8c90eb7b40707b446085620f1cd6034699e5fc854b9764340614355fc857553f306b21d23", 
 110 => x"9aada4f64c3329601ac8963c37efba533703ebc96d3d9ef4a9dde528ebd0be96efd04abdbf06056d59d9d8d6554d7683fc93b9539b263cff7b5b3e5ad7110695c71d79c87c73909a7039e60a58acba6423b6dd617eb96623cffca67f298bbff3c929e306da0ab79f0db5b5ab62d1f6fe01468ed862b57aa4ff8825157f3d2b62", 
 111 => x"eb6c1d37344b21e6b17511b797a32b632e638507099d756f0a2ad49a66e57d44462fc84c9cf14a2024b55f2b9e527ea55853263ab61962f643f2fc8c1f666cd21010673baf4f58df47d9f2afdbc8572fd23c74101efbd22177937d23736a5666912b7e12d9cc73a9e73200e2df6d7f42347b30e9e8d7ec855b3116d9ff711fcf", 
 112 => x"8ce197b99405224f2f1a2b57f71b14c9b48a310062d765218587c074cba51d987ca1404fd9389ac592f136484a0b212012c1f5a053f08a93177ebffe92c451a3980bdece7425ec43052ca703927c74c530c4556b303686483f65ba2fb2a23779a47ea7bd6a104c7aec695a2388a4f97dccfec10cd6074c1a11e815f2a2d79ef5", 
 113 => x"bf6116a7c453a95ab074d2228e523900be316d56792ea40d3143705ba8dae34ac0ad35d399ce4ef9561c4397ce0e6842618f8f753a7ec99a21676500b51f2333a8562d0b09dcdcba691058069bc48fff9059b16e3123e86d6a13460e991c15039f1b3edababe2b75f60c13086df34813e64d857b98f7c995d1cbe74746d0b5a9", 
 114 => x"380cfe7b9d170d915ca56d3954469126c8ad83bf012aaaf626eff12a8ef67ea89a845da53e1b248e810f6933cc6dc03c4373a023eb5149bddfa3981b270a1ac90c25a920e60802b60de783f2095a5e8d54a37fb915afc7139acd1c0eb13a0d434c6e6edc31880ec5183df2c76fe34aaebad099abcc6b309f8bf5558ff03b38cd", 
 115 => x"ef6cd209687e278904e67c02fb7fa0c11a44aa531aa6040a4acc8bbd058e426a58878bd8d5c1f8197063220a2b00fdb9309c3cfc0c358a09a668ede55b134fcfdfed9215a2478a9d088ed272578d37fd8967ec7a989a97360977fe8842f7acc634a8dba04d6a2edcf6b652c87c27e0d6a5f4808257c1be208d5567c4734e8639", 
 116 => x"7913edb2141ff39acbf23369c1e57a5cddbc3f3dbdb5f531f3de648f0d7c7926438bb66bf39b1380901376193e0b9d80d1144a9ba895e3e569591e6cadc79d23e67336a64b1970bbc3d5a2c022eb84b84731c1d1afe88907d85f3c223c2c03386d76eebdbc9b36f06bce2980407be98e3baf00a2524ac0d3e29369f6046da38c", 
 117 => x"808dcc92c54988de538adc61acea4452003c1ee3ed076879e2747f4048eb8a54bb1b42d5e8608ee72bc33a0349a975b127be07472614ce03b0ff9e6b366c6f1d2ae9c9263484972931f87dc168fe67784d74bc8d32d02b5ade0003a437ad5b873dcd2d9c377e903d4b4a089509fc82f32d95cb87cd02ab0af8964a1eeb748406", 
 118 => x"7096e908b9482be0ceb0f48a7f09c09fca2da0d21dca3b170ed3426c346a3e6cb88ea3ba323e6a296c32d200bed9ea601f3e42d5728391c53c6960b2b80242e21152b99454fa94c459d4abfd3aa59ef70a85161067a9499f4a57a74d16ea088eea9e20b5e70de67f46f051e8097fec1e5cb3804d3e9e0a763b7be894ebf8b935", 
 119 => x"4e0d618e382b28ecb9724b92f8f964bd77d4ec723e54f31bd08d261db36073ca26214e3eb5bdb5952edddd0d78d721dc842fab576042977b362ba2729559e894c166076534a84b43beb761255e3d9311b3d8a4eeabc912048bfdc125147cbd835421f0ab86d9fac1d3f4145dec22b5dc3006ec7ab18914f2a83d6d9895ad4115", 
 120 => x"9d3b07085ecc504f513a48edcfeed0aee89e36eb19b188169691080467c40d5c8a652142e3f5463faf8aa99dbd46828a978ebf1a91b0951cbb89766a664dc7170359dd4071400ad28231a72601c5f5b26ee8b01609bcdd606a82c835b8f2a14a3a90884c0051f234b907f2ecb7d9bb668304dd71fa3010060d59573c258c296d", 
 121 => x"ac31d028c595d5647328ea735316cfbaa966f20a7b00ccdd57d81f90d94f9ec832191f4b3f431bdfc50a1fb9fc80850506eb8c19a0f6352b2c21ffc5b142905924fa5b61550e042d0827c47ce574c49113ece559a19a2a1e6342e7620030bb59e4f4eca33e16616e7058a2916b44ba0e7f320a5fe6c61bec39ce9c1b8d2e779a", 
 122 => x"bbf2a751e7e0f830003db3a39acf3c5a4b553174695ac0f07189fcd1d0b7a3aba104bbaf484f2cfb742c7e2be6c3d055b044c37c399dbfb17228ad09c96fbbaa899a9ece47305dfc925d238ad094b4ab3dcdada740f547a9b01f98c87c24168d89fc719dc2e36898db8387bb807b444cc169c72192ccde8ddfb6b7eb8bb23d84", 
 123 => x"b8c2654c52b7b0ea20ee3956e587d026a205caadcc0ba50a29b3d635ca30ce90e2cb14079d60caee351daa5a1c869e153baf06b6eb34af88aa99ef0e0ee312da6e1c591a782142aeae317eb6125f77a25e46248654cba8c917c90aac01eb5ea6b67d91eae974eec9784ca5f69c3022fe79af0c80a09bb7d436a447bbfb70638d", 
 124 => x"e50c7fe496ce37cf35dc67e5c4fec0b1624db7c1b467025f0b204814561c01cb7293750ec68df656bbbca2b5ca57914f13c82daf68bc9d21af5370d633d282b6d5864b8c399a9b8f75ed26984fde69fed3a7b8d2be7d352d16ef2533720b0fa9ee929d6711ceca5b0c31a7f50a80b504002999d1c201573991633f06b9d1cdfe", 
 125 => x"6a043e569f4c8bdc2e205774a1fa001124ea006bea4d5377375ad800876cfc67425e5f74b30507df2960597113467e1954ed45496ccda25134090c288d20afbc27366b3b551be4212ff7f81ab17200784693adc2a920b79670014c9e54a7bc65ad7dc391d43244aa8ea4fc3c82ccbdac3574e46269294883b22154200536d609", 
 126 => x"ca1b0fe269abd1380ed6fb661a03bc0a951c71d81638847cecaeea9ba7ed16b79b3b31726fc3115cb2418f1e3e651e7d07037b4495cba234190034ca4c79f35a3a9623062dd4b6a95373ba6251e7635c6848d5fa3bc270c39b94ea5d71965dc0a227449b00519bdd223d45960646dd2b939fe07ccd87004d4d6724e810c5bd79", 
 127 => x"d3d1af79aa0ea3c747a2c68c72e0106bca05b8a66d5232aad30361922f15fcf10428b95f42f2b073daf865423d7080ee22662d0db5cee2061c97e88298d0f662afff213781066b96e71aaa2008f0bf1024d03e55ea5a77b5afa7a80e65d4ebd75309f0241365946a5968a23350a864f5d410e5da1cfbf1d9c27414e3744767ad"
  ); 
--signal pca_w01  : std_logic_vector(7 downto 0); 
--signal pca_w02  : std_logic_vector(7 downto 0); 
--signal pca_w03  : std_logic_vector(7 downto 0); 
--signal pca_w04  : std_logic_vector(7 downto 0); 
--signal pca_w05  : std_logic_vector(7 downto 0); 
--signal pca_w06  : std_logic_vector(7 downto 0); 
--signal pca_w07  : std_logic_vector(7 downto 0); 
--signal pca_w08  : std_logic_vector(7 downto 0); 
--signal pca_w09  : std_logic_vector(7 downto 0); 
--signal pca_w10  : std_logic_vector(7 downto 0); 
--signal pca_w11  : std_logic_vector(7 downto 0); 
--signal pca_w12  : std_logic_vector(7 downto 0); 
--signal pca_w13  : std_logic_vector(7 downto 0); 
--signal pca_w14  : std_logic_vector(7 downto 0); 
--signal pca_w15  : std_logic_vector(7 downto 0); 
--signal pca_w16  : std_logic_vector(7 downto 0); 
--signal pca_w17  : std_logic_vector(7 downto 0); 
--signal pca_w18  : std_logic_vector(7 downto 0); 
--signal pca_w19  : std_logic_vector(7 downto 0); 
--signal pca_w20  : std_logic_vector(7 downto 0); 
--signal pca_w21  : std_logic_vector(7 downto 0); 
--signal pca_w22  : std_logic_vector(7 downto 0); 
--signal pca_w23  : std_logic_vector(7 downto 0); 
--signal pca_w24  : std_logic_vector(7 downto 0); 
--signal pca_w25  : std_logic_vector(7 downto 0); 
--signal pca_w26  : std_logic_vector(7 downto 0); 
--signal pca_w27  : std_logic_vector(7 downto 0); 
--signal pca_w28  : std_logic_vector(7 downto 0); 
--signal pca_w29  : std_logic_vector(7 downto 0); 
--signal pca_w30  : std_logic_vector(7 downto 0); 
--signal pca_w31  : std_logic_vector(7 downto 0); 
--signal pca_w32  : std_logic_vector(7 downto 0); 
--signal pca_w33  : std_logic_vector(7 downto 0); 
--signal pca_w34  : std_logic_vector(7 downto 0); 
--signal pca_w35  : std_logic_vector(7 downto 0); 
--signal pca_w36  : std_logic_vector(7 downto 0); 
--signal pca_w37  : std_logic_vector(7 downto 0); 
--signal pca_w38  : std_logic_vector(7 downto 0); 
--signal pca_w39  : std_logic_vector(7 downto 0); 
--signal pca_w40  : std_logic_vector(7 downto 0); 
--signal pca_w41  : std_logic_vector(7 downto 0); 
--signal pca_w42  : std_logic_vector(7 downto 0); 
--signal pca_w43  : std_logic_vector(7 downto 0); 
--signal pca_w44  : std_logic_vector(7 downto 0); 
--signal pca_w45  : std_logic_vector(7 downto 0); 
--signal pca_w46  : std_logic_vector(7 downto 0); 
--signal pca_w47  : std_logic_vector(7 downto 0); 
--signal pca_w48  : std_logic_vector(7 downto 0); 
--signal pca_w49  : std_logic_vector(7 downto 0); 
--signal pca_w50  : std_logic_vector(7 downto 0); 
--signal pca_w51  : std_logic_vector(7 downto 0); 
--signal pca_w52  : std_logic_vector(7 downto 0); 
--signal pca_w53  : std_logic_vector(7 downto 0); 
--signal pca_w54  : std_logic_vector(7 downto 0); 
--signal pca_w55  : std_logic_vector(7 downto 0); 
--signal pca_w56  : std_logic_vector(7 downto 0); 
--signal pca_w57  : std_logic_vector(7 downto 0); 
--signal pca_w58  : std_logic_vector(7 downto 0); 
--signal pca_w59  : std_logic_vector(7 downto 0); 
--signal pca_w60  : std_logic_vector(7 downto 0); 
--signal pca_w61  : std_logic_vector(7 downto 0); 
--signal pca_w62  : std_logic_vector(7 downto 0); 
--signal pca_w63  : std_logic_vector(7 downto 0); 
--signal pca_w64  : std_logic_vector(7 downto 0); 

signal pca_w_data     : std_logic_vector(64*8-1 downto 0);
signal pca_w_addr     : std_logic_vector(5 downto 0);
signal pca_col_count  : std_logic_vector(7 downto 0); --max 265 columns

signal pca_d01_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d02_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d03_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d04_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d05_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d06_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d07_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d08_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d09_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d10_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d11_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d12_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d13_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d14_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d15_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d16_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d17_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d18_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d19_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d20_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d21_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d22_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d23_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d24_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d25_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d26_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d27_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d28_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d29_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d30_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d31_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d32_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d33_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d34_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d35_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d36_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d37_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d38_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d39_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d40_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d41_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d42_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d43_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d44_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d45_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d46_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d47_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d48_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d49_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d50_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d51_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d52_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d53_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d54_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d55_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d56_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d57_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d58_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d59_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d60_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d61_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d62_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d63_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d64_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);


signal pca_d65_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d66_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d67_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d68_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d69_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d70_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d71_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d72_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d73_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d74_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d75_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d76_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d77_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d78_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d79_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d80_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d81_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d82_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d83_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d84_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d85_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d86_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d87_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d88_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d89_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d90_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d91_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d92_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d93_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d94_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d95_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d96_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d97_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d98_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d99_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d100_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d101_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d102_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d103_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d104_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d105_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d106_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d107_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d108_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d109_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d110_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d111_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d112_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d113_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d114_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d115_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d116_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d117_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d118_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d119_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d120_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d121_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d122_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d123_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d124_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d125_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d126_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d127_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);
signal pca_d128_out   : std_logic_vector(CL_W + PCAweightW + 5 downto 0);

signal pca_en_out  : std_logic;
signal pca_sof_out : std_logic;

signal d_tmp_1_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_2_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_3_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_4_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_5_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_6_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_7_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_8_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_9_out   : std_logic_vector (Wb-1 downto 0);
signal d_tmp_10_out  : std_logic_vector (Wb-1 downto 0);
signal d_tmp_11_out  : std_logic_vector (Wb-1 downto 0);
signal d_tmp_12_out  : std_logic_vector (Wb-1 downto 0);
signal d_tmp_13_out  : std_logic_vector (Wb-1 downto 0);
signal d_tmp_14_out  : std_logic_vector (Wb-1 downto 0);
signal d_tmp_15_out  : std_logic_vector (Wb-1 downto 0);
signal d_tmp_16_out  : std_logic_vector (Wb-1 downto 0);


type Huff_code_type  is array ( 0 to 255 ) of std_logic_vector(Huff_wid-1 downto 0);
type Huff_width_type is array ( 0 to 255 ) of std_logic_vector(         3 downto 0);

constant Huff_code  : Huff_code_type  := ( 0 => x"003", 1 => x"037", 2 => x"932", 3 => x"124", 4 => x"611", 5 => x"027", 6 => x"523", 7 => x"630", 8 => x"121", 9 => x"361", others => x"BAD"); 
constant Huff_width : Huff_width_type := ( 0 => x"4", 1 => x"8",  2 => x"C",   3 => x"C",   4 => x"C",   5 => x"8",  6 => x"C",   7 => x"C",   8 => x"C",   9 => x"C",   others => x"C"); 

signal h_en          : std_logic;
signal h_count_en    : std_logic;
signal h_count_en2   : std_logic;
signal h_count       : std_logic_vector(         7 downto 0);
signal alpha_data    : std_logic_vector(         7 downto 0);
signal alpha_code    : std_logic_vector(Huff_wid-1 downto 0);
signal alpha_width   : std_logic_vector(         3 downto 0);



signal huff_out      : std_logic_vector (Wb-1 downto 0);

-- PCA disable signals
signal PCA_dis1, PCA_dis2, PCA_dis3, PCA_dis4, PCA_dis5, PCA_dis6, PCA_dis7, PCA_dis8, PCA_dis9 , PCA_dis10, PCA_dis11, PCA_dis12, PCA_dis13, PCA_dis14, PCA_dis15, PCA_dis16  : std_logic_vector(7 downto 0);
begin

-- weight init

  p_weight1 : process (clk,rst)
  begin
    if rst = '1' then
       w_en        <= '0';
       w_count_en  <= '1';
       w_count_en2 <= '0';
       w_count     <= (others => '0');
    elsif rising_edge(clk) then
       if w_count_en = '1' then
          w_num   <= w_count;
          w_count <= w_count + 1;
       end if;
       if w_count = (2**(w_count'left+1) - 1) then
          w_count_en <= '0';
       end if;
       w_count_en2 <= w_count_en;
       w_en        <= w_count_en2;
    end if;
  end process p_weight1;

  p_weight2 : process (clk)
  begin
    if rising_edge(clk) then
       w01_in <=  weight01(conv_integer('0' & w_count));
       w02_in <=  weight02(conv_integer('0' & w_count));
       w03_in <=  weight03(conv_integer('0' & w_count));
       w04_in <=  weight04(conv_integer('0' & w_count));
       w05_in <=  weight05(conv_integer('0' & w_count));
       w06_in <=  weight06(conv_integer('0' & w_count));
       w07_in <=  weight07(conv_integer('0' & w_count));
       w08_in <=  weight08(conv_integer('0' & w_count));
       w09_in <=  weight09(conv_integer('0' & w_count));
       w10_in <=  weight10(conv_integer('0' & w_count));
       w11_in <=  weight11(conv_integer('0' & w_count));
       w12_in <=  weight12(conv_integer('0' & w_count));
       w13_in <=  weight13(conv_integer('0' & w_count));
       w14_in <=  weight14(conv_integer('0' & w_count));
       w15_in <=  weight15(conv_integer('0' & w_count));
       w16_in <=  weight16(conv_integer('0' & w_count));
       w17_in <=  weight17(conv_integer('0' & w_count));
       w18_in <=  weight18(conv_integer('0' & w_count));
       w19_in <=  weight19(conv_integer('0' & w_count));
       w20_in <=  weight20(conv_integer('0' & w_count));
       w21_in <=  weight21(conv_integer('0' & w_count));
       w22_in <=  weight22(conv_integer('0' & w_count));
       w23_in <=  weight23(conv_integer('0' & w_count));
       w24_in <=  weight24(conv_integer('0' & w_count));
       w25_in <=  weight25(conv_integer('0' & w_count));
       w26_in <=  weight26(conv_integer('0' & w_count));
       w27_in <=  weight27(conv_integer('0' & w_count));
       w28_in <=  weight28(conv_integer('0' & w_count));
       w29_in <=  weight29(conv_integer('0' & w_count));
       w30_in <=  weight30(conv_integer('0' & w_count));
       w31_in <=  weight31(conv_integer('0' & w_count));
       w32_in <=  weight32(conv_integer('0' & w_count));
       w33_in <=  weight33(conv_integer('0' & w_count));
       w34_in <=  weight34(conv_integer('0' & w_count));
       w35_in <=  weight35(conv_integer('0' & w_count));
       w36_in <=  weight36(conv_integer('0' & w_count));
       w37_in <=  weight37(conv_integer('0' & w_count));
       w38_in <=  weight38(conv_integer('0' & w_count));
       w39_in <=  weight39(conv_integer('0' & w_count));
       w40_in <=  weight40(conv_integer('0' & w_count));
       w41_in <=  weight41(conv_integer('0' & w_count));
       w42_in <=  weight42(conv_integer('0' & w_count));
       w43_in <=  weight43(conv_integer('0' & w_count));
       w44_in <=  weight44(conv_integer('0' & w_count));
       w45_in <=  weight45(conv_integer('0' & w_count));
       w46_in <=  weight46(conv_integer('0' & w_count));
       w47_in <=  weight47(conv_integer('0' & w_count));
       w48_in <=  weight48(conv_integer('0' & w_count));
       w49_in <=  weight49(conv_integer('0' & w_count));
       w50_in <=  weight50(conv_integer('0' & w_count));
       w51_in <=  weight51(conv_integer('0' & w_count));
       w52_in <=  weight52(conv_integer('0' & w_count));
       w53_in <=  weight53(conv_integer('0' & w_count));
       w54_in <=  weight54(conv_integer('0' & w_count));
       w55_in <=  weight55(conv_integer('0' & w_count));
       w56_in <=  weight56(conv_integer('0' & w_count));
       w57_in <=  weight57(conv_integer('0' & w_count));
       w58_in <=  weight58(conv_integer('0' & w_count));
       w59_in <=  weight59(conv_integer('0' & w_count));
       w60_in <=  weight60(conv_integer('0' & w_count));
       w61_in <=  weight61(conv_integer('0' & w_count));
       w62_in <=  weight62(conv_integer('0' & w_count));
       w63_in <=  weight63(conv_integer('0' & w_count));
       w64_in <=  weight64(conv_integer('0' & w_count));


       w65_in <=  weight01(conv_integer('0' & w_count));
       w66_in <=  weight02(conv_integer('0' & w_count));
       w67_in <=  weight03(conv_integer('0' & w_count));
       w68_in <=  weight04(conv_integer('0' & w_count));
       w69_in <=  weight05(conv_integer('0' & w_count));
       w70_in <=  weight06(conv_integer('0' & w_count));
       w71_in <=  weight07(conv_integer('0' & w_count));
       w72_in <=  weight08(conv_integer('0' & w_count));
       w73_in <=  weight09(conv_integer('0' & w_count));
       w74_in <=  weight10(conv_integer('0' & w_count));
       w75_in <=  weight11(conv_integer('0' & w_count));
       w76_in <=  weight12(conv_integer('0' & w_count));
       w77_in <=  weight13(conv_integer('0' & w_count));
       w78_in <=  weight14(conv_integer('0' & w_count));
       w79_in <=  weight15(conv_integer('0' & w_count));
       w80_in <=  weight16(conv_integer('0' & w_count));
       w81_in <=  weight17(conv_integer('0' & w_count));
       w82_in <=  weight18(conv_integer('0' & w_count));
       w83_in <=  weight19(conv_integer('0' & w_count));
       w84_in <=  weight20(conv_integer('0' & w_count));
       w85_in <=  weight21(conv_integer('0' & w_count));
       w86_in <=  weight22(conv_integer('0' & w_count));
       w87_in <=  weight23(conv_integer('0' & w_count));
       w88_in <=  weight24(conv_integer('0' & w_count));
       w89_in <=  weight25(conv_integer('0' & w_count));
       w90_in <=  weight26(conv_integer('0' & w_count));
       w91_in <=  weight27(conv_integer('0' & w_count));
       w92_in <=  weight28(conv_integer('0' & w_count));
       w93_in <=  weight29(conv_integer('0' & w_count));
       w94_in <=  weight30(conv_integer('0' & w_count));
       w95_in <=  weight31(conv_integer('0' & w_count));
       w96_in <=  weight32(conv_integer('0' & w_count));
       w97_in <=  weight33(conv_integer('0' & w_count));
       w98_in <=  weight34(conv_integer('0' & w_count));
       w99_in <=  weight35(conv_integer('0' & w_count));
       w100_in <=  weight36(conv_integer('0' & w_count));
       w101_in <=  weight37(conv_integer('0' & w_count));
       w102_in <=  weight38(conv_integer('0' & w_count));
       w103_in <=  weight39(conv_integer('0' & w_count));
       w104_in <=  weight40(conv_integer('0' & w_count));
       w105_in <=  weight41(conv_integer('0' & w_count));
       w106_in <=  weight42(conv_integer('0' & w_count));
       w107_in <=  weight43(conv_integer('0' & w_count));
       w108_in <=  weight44(conv_integer('0' & w_count));
       w109_in <=  weight45(conv_integer('0' & w_count));
       w110_in <=  weight46(conv_integer('0' & w_count));
       w111_in <=  weight47(conv_integer('0' & w_count));
       w112_in <=  weight48(conv_integer('0' & w_count));
       w113_in <=  weight49(conv_integer('0' & w_count));
       w114_in <=  weight50(conv_integer('0' & w_count));
       w115_in <=  weight51(conv_integer('0' & w_count));
       w116_in <=  weight52(conv_integer('0' & w_count));
       w117_in <=  weight53(conv_integer('0' & w_count));
       w118_in <=  weight54(conv_integer('0' & w_count));
       w119_in <=  weight55(conv_integer('0' & w_count));
       w120_in <=  weight56(conv_integer('0' & w_count));
       w121_in <=  weight57(conv_integer('0' & w_count));
       w122_in <=  weight58(conv_integer('0' & w_count));
       w123_in <=  weight59(conv_integer('0' & w_count));
       w124_in <=  weight60(conv_integer('0' & w_count));
       w125_in <=  weight61(conv_integer('0' & w_count));
       w126_in <=  weight62(conv_integer('0' & w_count));
       w127_in <=  weight63(conv_integer('0' & w_count));
       w128_in <=  weight64(conv_integer('0' & w_count));

    end if;
  end process p_weight2;

CL01: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w01_in, w_num => w_num, w_en => w_en, d_out => d01_out1, en_out => cl_en_out, sof_out => cl_sof_out);
CL02: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w02_in, w_num => w_num, w_en => w_en, d_out => d02_out1, en_out => open, sof_out => open);
CL03: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w03_in, w_num => w_num, w_en => w_en, d_out => d03_out1, en_out => open, sof_out => open);
CL04: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w04_in, w_num => w_num, w_en => w_en, d_out => d04_out1, en_out => open, sof_out => open);
CL05: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w05_in, w_num => w_num, w_en => w_en, d_out => d05_out1, en_out => open, sof_out => open);
CL06: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w06_in, w_num => w_num, w_en => w_en, d_out => d06_out1, en_out => open, sof_out => open);
CL07: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w07_in, w_num => w_num, w_en => w_en, d_out => d07_out1, en_out => open, sof_out => open);
CL08: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w08_in, w_num => w_num, w_en => w_en, d_out => d08_out1, en_out => open, sof_out => open);
CL09: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w09_in, w_num => w_num, w_en => w_en, d_out => d09_out1, en_out => open, sof_out => open);
CL10: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w10_in, w_num => w_num, w_en => w_en, d_out => d10_out1, en_out => open, sof_out => open);
CL11: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w11_in, w_num => w_num, w_en => w_en, d_out => d11_out1, en_out => open, sof_out => open);
CL12: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w12_in, w_num => w_num, w_en => w_en, d_out => d12_out1, en_out => open, sof_out => open);
CL13: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w13_in, w_num => w_num, w_en => w_en, d_out => d13_out1, en_out => open, sof_out => open);
CL14: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w14_in, w_num => w_num, w_en => w_en, d_out => d14_out1, en_out => open, sof_out => open);
CL15: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w15_in, w_num => w_num, w_en => w_en, d_out => d15_out1, en_out => open, sof_out => open);
CL16: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w16_in, w_num => w_num, w_en => w_en, d_out => d16_out1, en_out => open, sof_out => open);
CL17: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w17_in, w_num => w_num, w_en => w_en, d_out => d17_out1, en_out => open, sof_out => open);
CL18: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w18_in, w_num => w_num, w_en => w_en, d_out => d18_out1, en_out => open, sof_out => open);
CL19: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w19_in, w_num => w_num, w_en => w_en, d_out => d19_out1, en_out => open, sof_out => open);
CL20: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w20_in, w_num => w_num, w_en => w_en, d_out => d20_out1, en_out => open, sof_out => open);
CL21: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w21_in, w_num => w_num, w_en => w_en, d_out => d21_out1, en_out => open, sof_out => open);
CL22: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w22_in, w_num => w_num, w_en => w_en, d_out => d22_out1, en_out => open, sof_out => open);
CL23: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w23_in, w_num => w_num, w_en => w_en, d_out => d23_out1, en_out => open, sof_out => open);
CL24: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w24_in, w_num => w_num, w_en => w_en, d_out => d24_out1, en_out => open, sof_out => open);
CL25: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w25_in, w_num => w_num, w_en => w_en, d_out => d25_out1, en_out => open, sof_out => open);
CL26: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w26_in, w_num => w_num, w_en => w_en, d_out => d26_out1, en_out => open, sof_out => open);
CL27: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w27_in, w_num => w_num, w_en => w_en, d_out => d27_out1, en_out => open, sof_out => open);
CL28: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w28_in, w_num => w_num, w_en => w_en, d_out => d28_out1, en_out => open, sof_out => open);
CL29: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w29_in, w_num => w_num, w_en => w_en, d_out => d29_out1, en_out => open, sof_out => open);
CL30: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w30_in, w_num => w_num, w_en => w_en, d_out => d30_out1, en_out => open, sof_out => open);
CL31: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w31_in, w_num => w_num, w_en => w_en, d_out => d31_out1, en_out => open, sof_out => open);
CL32: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w32_in, w_num => w_num, w_en => w_en, d_out => d32_out1, en_out => open, sof_out => open);
CL33: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w33_in, w_num => w_num, w_en => w_en, d_out => d33_out1, en_out => open, sof_out => open);
CL34: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w34_in, w_num => w_num, w_en => w_en, d_out => d34_out1, en_out => open, sof_out => open);
CL35: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w35_in, w_num => w_num, w_en => w_en, d_out => d35_out1, en_out => open, sof_out => open);
CL36: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w36_in, w_num => w_num, w_en => w_en, d_out => d36_out1, en_out => open, sof_out => open);
CL37: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w37_in, w_num => w_num, w_en => w_en, d_out => d37_out1, en_out => open, sof_out => open);
CL38: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w38_in, w_num => w_num, w_en => w_en, d_out => d38_out1, en_out => open, sof_out => open);
CL39: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w39_in, w_num => w_num, w_en => w_en, d_out => d39_out1, en_out => open, sof_out => open);
CL40: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w40_in, w_num => w_num, w_en => w_en, d_out => d40_out1, en_out => open, sof_out => open);
CL41: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w41_in, w_num => w_num, w_en => w_en, d_out => d41_out1, en_out => open, sof_out => open);
CL42: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w42_in, w_num => w_num, w_en => w_en, d_out => d42_out1, en_out => open, sof_out => open);
CL43: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w43_in, w_num => w_num, w_en => w_en, d_out => d43_out1, en_out => open, sof_out => open);
CL44: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w44_in, w_num => w_num, w_en => w_en, d_out => d44_out1, en_out => open, sof_out => open);
CL45: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w45_in, w_num => w_num, w_en => w_en, d_out => d45_out1, en_out => open, sof_out => open);
CL46: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w46_in, w_num => w_num, w_en => w_en, d_out => d46_out1, en_out => open, sof_out => open);
CL47: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w47_in, w_num => w_num, w_en => w_en, d_out => d47_out1, en_out => open, sof_out => open);
CL48: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w48_in, w_num => w_num, w_en => w_en, d_out => d48_out1, en_out => open, sof_out => open);
CL49: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w49_in, w_num => w_num, w_en => w_en, d_out => d49_out1, en_out => open, sof_out => open);
CL50: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w50_in, w_num => w_num, w_en => w_en, d_out => d50_out1, en_out => open, sof_out => open);
CL51: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w51_in, w_num => w_num, w_en => w_en, d_out => d51_out1, en_out => open, sof_out => open);
CL52: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w52_in, w_num => w_num, w_en => w_en, d_out => d52_out1, en_out => open, sof_out => open);
CL53: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w53_in, w_num => w_num, w_en => w_en, d_out => d53_out1, en_out => open, sof_out => open);
CL54: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w54_in, w_num => w_num, w_en => w_en, d_out => d54_out1, en_out => open, sof_out => open);
CL55: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w55_in, w_num => w_num, w_en => w_en, d_out => d55_out1, en_out => open, sof_out => open);
CL56: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w56_in, w_num => w_num, w_en => w_en, d_out => d56_out1, en_out => open, sof_out => open);
CL57: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w57_in, w_num => w_num, w_en => w_en, d_out => d57_out1, en_out => open, sof_out => open);
CL58: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w58_in, w_num => w_num, w_en => w_en, d_out => d58_out1, en_out => open, sof_out => open);
CL59: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w59_in, w_num => w_num, w_en => w_en, d_out => d59_out1, en_out => open, sof_out => open);
CL60: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w60_in, w_num => w_num, w_en => w_en, d_out => d60_out1, en_out => open, sof_out => open);
CL61: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w61_in, w_num => w_num, w_en => w_en, d_out => d61_out1, en_out => open, sof_out => open);
CL62: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w62_in, w_num => w_num, w_en => w_en, d_out => d62_out1, en_out => open, sof_out => open);
CL63: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w63_in, w_num => w_num, w_en => w_en, d_out => d63_out1, en_out => open, sof_out => open);
CL64: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w64_in, w_num => w_num, w_en => w_en, d_out => d64_out1, en_out => open, sof_out => open);

CL65 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w65_in,  w_num => w_num, w_en => w_en, d_out => d65_out1 , en_out => open, sof_out => open);
CL66 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w66_in,  w_num => w_num, w_en => w_en, d_out => d66_out1 , en_out => open, sof_out => open);
CL67 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w67_in,  w_num => w_num, w_en => w_en, d_out => d67_out1 , en_out => open, sof_out => open);
CL68 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w68_in,  w_num => w_num, w_en => w_en, d_out => d68_out1 , en_out => open, sof_out => open);
CL69 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w69_in,  w_num => w_num, w_en => w_en, d_out => d69_out1 , en_out => open, sof_out => open);
CL70 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w70_in,  w_num => w_num, w_en => w_en, d_out => d70_out1 , en_out => open, sof_out => open);
CL71 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w71_in,  w_num => w_num, w_en => w_en, d_out => d71_out1 , en_out => open, sof_out => open);
CL72 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w72_in,  w_num => w_num, w_en => w_en, d_out => d72_out1 , en_out => open, sof_out => open);
CL73 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w73_in,  w_num => w_num, w_en => w_en, d_out => d73_out1 , en_out => open, sof_out => open);
CL74 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w74_in,  w_num => w_num, w_en => w_en, d_out => d74_out1 , en_out => open, sof_out => open);
CL75 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w75_in,  w_num => w_num, w_en => w_en, d_out => d75_out1 , en_out => open, sof_out => open);
CL76 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w76_in,  w_num => w_num, w_en => w_en, d_out => d76_out1 , en_out => open, sof_out => open);
CL77 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w77_in,  w_num => w_num, w_en => w_en, d_out => d77_out1 , en_out => open, sof_out => open);
CL78 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w78_in,  w_num => w_num, w_en => w_en, d_out => d78_out1 , en_out => open, sof_out => open);
CL79 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w79_in,  w_num => w_num, w_en => w_en, d_out => d79_out1 , en_out => open, sof_out => open);
CL80 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w80_in,  w_num => w_num, w_en => w_en, d_out => d80_out1 , en_out => open, sof_out => open);
CL81 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w81_in,  w_num => w_num, w_en => w_en, d_out => d81_out1 , en_out => open, sof_out => open);
CL82 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w82_in,  w_num => w_num, w_en => w_en, d_out => d82_out1 , en_out => open, sof_out => open);
CL83 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w83_in,  w_num => w_num, w_en => w_en, d_out => d83_out1 , en_out => open, sof_out => open);
CL84 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w84_in,  w_num => w_num, w_en => w_en, d_out => d84_out1 , en_out => open, sof_out => open);
CL85 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w85_in,  w_num => w_num, w_en => w_en, d_out => d85_out1 , en_out => open, sof_out => open);
CL86 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w86_in,  w_num => w_num, w_en => w_en, d_out => d86_out1 , en_out => open, sof_out => open);
CL87 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w87_in,  w_num => w_num, w_en => w_en, d_out => d87_out1 , en_out => open, sof_out => open);
CL88 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w88_in,  w_num => w_num, w_en => w_en, d_out => d88_out1 , en_out => open, sof_out => open);
CL89 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w89_in,  w_num => w_num, w_en => w_en, d_out => d89_out1 , en_out => open, sof_out => open);
CL90 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w90_in,  w_num => w_num, w_en => w_en, d_out => d90_out1 , en_out => open, sof_out => open);
CL91 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w91_in,  w_num => w_num, w_en => w_en, d_out => d91_out1 , en_out => open, sof_out => open);
CL92 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w92_in,  w_num => w_num, w_en => w_en, d_out => d92_out1 , en_out => open, sof_out => open);
CL93 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w93_in,  w_num => w_num, w_en => w_en, d_out => d93_out1 , en_out => open, sof_out => open);
CL94 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w94_in,  w_num => w_num, w_en => w_en, d_out => d94_out1 , en_out => open, sof_out => open);
CL95 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w95_in,  w_num => w_num, w_en => w_en, d_out => d95_out1 , en_out => open, sof_out => open);
CL96 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w96_in,  w_num => w_num, w_en => w_en, d_out => d96_out1 , en_out => open, sof_out => open);
CL97 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w97_in,  w_num => w_num, w_en => w_en, d_out => d97_out1 , en_out => open, sof_out => open);
CL98 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w98_in,  w_num => w_num, w_en => w_en, d_out => d98_out1 , en_out => open, sof_out => open);
CL99 : ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w99_in,  w_num => w_num, w_en => w_en, d_out => d99_out1 , en_out => open, sof_out => open);
CL100: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w100_in, w_num => w_num, w_en => w_en, d_out => d100_out1, en_out => open, sof_out => open);
CL101: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w101_in, w_num => w_num, w_en => w_en, d_out => d101_out1, en_out => open, sof_out => open);
CL102: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w102_in, w_num => w_num, w_en => w_en, d_out => d102_out1, en_out => open, sof_out => open);
CL103: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w103_in, w_num => w_num, w_en => w_en, d_out => d103_out1, en_out => open, sof_out => open);
CL104: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w104_in, w_num => w_num, w_en => w_en, d_out => d104_out1, en_out => open, sof_out => open);
CL105: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w105_in, w_num => w_num, w_en => w_en, d_out => d105_out1, en_out => open, sof_out => open);
CL106: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w106_in, w_num => w_num, w_en => w_en, d_out => d106_out1, en_out => open, sof_out => open);
CL107: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w107_in, w_num => w_num, w_en => w_en, d_out => d107_out1, en_out => open, sof_out => open);
CL108: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w108_in, w_num => w_num, w_en => w_en, d_out => d108_out1, en_out => open, sof_out => open);
CL109: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w109_in, w_num => w_num, w_en => w_en, d_out => d109_out1, en_out => open, sof_out => open);
CL110: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w110_in, w_num => w_num, w_en => w_en, d_out => d110_out1, en_out => open, sof_out => open);
CL111: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w111_in, w_num => w_num, w_en => w_en, d_out => d111_out1, en_out => open, sof_out => open);
CL112: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w112_in, w_num => w_num, w_en => w_en, d_out => d112_out1, en_out => open, sof_out => open);
CL113: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w113_in, w_num => w_num, w_en => w_en, d_out => d113_out1, en_out => open, sof_out => open);
CL114: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w114_in, w_num => w_num, w_en => w_en, d_out => d114_out1, en_out => open, sof_out => open);
CL115: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w115_in, w_num => w_num, w_en => w_en, d_out => d115_out1, en_out => open, sof_out => open);
CL116: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w116_in, w_num => w_num, w_en => w_en, d_out => d116_out1, en_out => open, sof_out => open);
CL117: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w117_in, w_num => w_num, w_en => w_en, d_out => d117_out1, en_out => open, sof_out => open);
CL118: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w118_in, w_num => w_num, w_en => w_en, d_out => d118_out1, en_out => open, sof_out => open);
CL119: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w119_in, w_num => w_num, w_en => w_en, d_out => d119_out1, en_out => open, sof_out => open);
CL120: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w120_in, w_num => w_num, w_en => w_en, d_out => d120_out1, en_out => open, sof_out => open);
CL121: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w121_in, w_num => w_num, w_en => w_en, d_out => d121_out1, en_out => open, sof_out => open);
CL122: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w122_in, w_num => w_num, w_en => w_en, d_out => d122_out1, en_out => open, sof_out => open);
CL123: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w123_in, w_num => w_num, w_en => w_en, d_out => d123_out1, en_out => open, sof_out => open);
CL124: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w124_in, w_num => w_num, w_en => w_en, d_out => d124_out1, en_out => open, sof_out => open);
CL125: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w125_in, w_num => w_num, w_en => w_en, d_out => d125_out1, en_out => open, sof_out => open);
CL126: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w126_in, w_num => w_num, w_en => w_en, d_out => d126_out1, en_out => open, sof_out => open);
CL127: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w127_in, w_num => w_num, w_en => w_en, d_out => d127_out1, en_out => open, sof_out => open);
CL128: ConvLayer128 generic map (mult_sum => mult_sum_CL,N => N,M => CL_w_width,W => CL_W,SR => CL_SR,in_row => in_row, in_col => in_col)port map ( clk => clk, rst => rst, d_in => d_in, en_in => en_in, sof_in => sof_in, w_in => w128_in, w_num => w_num, w_en => w_en, d_out => d128_out1, en_out => open, sof_out => open);


d01_out(7 downto 0) <= d01_out1(d01_out1'left downto d01_out1'left -7);
d02_out(7 downto 0) <= d02_out1(d02_out1'left downto d02_out1'left -7);
d03_out(7 downto 0) <= d03_out1(d03_out1'left downto d03_out1'left -7);
d04_out(7 downto 0) <= d04_out1(d04_out1'left downto d04_out1'left -7);
d05_out(7 downto 0) <= d05_out1(d05_out1'left downto d05_out1'left -7);
d06_out(7 downto 0) <= d06_out1(d06_out1'left downto d06_out1'left -7);
d07_out(7 downto 0) <= d07_out1(d07_out1'left downto d07_out1'left -7);
d08_out(7 downto 0) <= d08_out1(d08_out1'left downto d08_out1'left -7);
d09_out(7 downto 0) <= d09_out1(d09_out1'left downto d09_out1'left -7);
d10_out(7 downto 0) <= d10_out1(d10_out1'left downto d10_out1'left -7);
d11_out(7 downto 0) <= d11_out1(d11_out1'left downto d11_out1'left -7);
d12_out(7 downto 0) <= d12_out1(d12_out1'left downto d12_out1'left -7);
d13_out(7 downto 0) <= d13_out1(d13_out1'left downto d13_out1'left -7);
d14_out(7 downto 0) <= d14_out1(d14_out1'left downto d14_out1'left -7);
d15_out(7 downto 0) <= d15_out1(d15_out1'left downto d15_out1'left -7);
d16_out(7 downto 0) <= d16_out1(d16_out1'left downto d16_out1'left -7);
d17_out(7 downto 0) <= d17_out1(d17_out1'left downto d17_out1'left -7);
d18_out(7 downto 0) <= d18_out1(d18_out1'left downto d18_out1'left -7);
d19_out(7 downto 0) <= d19_out1(d19_out1'left downto d19_out1'left -7);
d20_out(7 downto 0) <= d20_out1(d20_out1'left downto d20_out1'left -7);
d21_out(7 downto 0) <= d21_out1(d21_out1'left downto d21_out1'left -7);
d22_out(7 downto 0) <= d22_out1(d22_out1'left downto d22_out1'left -7);
d23_out(7 downto 0) <= d23_out1(d23_out1'left downto d23_out1'left -7);
d24_out(7 downto 0) <= d24_out1(d24_out1'left downto d24_out1'left -7);
d25_out(7 downto 0) <= d25_out1(d25_out1'left downto d25_out1'left -7);
d26_out(7 downto 0) <= d26_out1(d26_out1'left downto d26_out1'left -7);
d27_out(7 downto 0) <= d27_out1(d27_out1'left downto d27_out1'left -7);
d28_out(7 downto 0) <= d28_out1(d28_out1'left downto d28_out1'left -7);
d29_out(7 downto 0) <= d29_out1(d29_out1'left downto d29_out1'left -7);
d30_out(7 downto 0) <= d30_out1(d30_out1'left downto d30_out1'left -7);
d31_out(7 downto 0) <= d31_out1(d31_out1'left downto d31_out1'left -7);
d32_out(7 downto 0) <= d32_out1(d32_out1'left downto d32_out1'left -7);
d33_out(7 downto 0) <= d33_out1(d33_out1'left downto d33_out1'left -7);
d34_out(7 downto 0) <= d34_out1(d34_out1'left downto d34_out1'left -7);
d35_out(7 downto 0) <= d35_out1(d35_out1'left downto d35_out1'left -7);
d36_out(7 downto 0) <= d36_out1(d36_out1'left downto d36_out1'left -7);
d37_out(7 downto 0) <= d37_out1(d37_out1'left downto d37_out1'left -7);
d38_out(7 downto 0) <= d38_out1(d38_out1'left downto d38_out1'left -7);
d39_out(7 downto 0) <= d39_out1(d39_out1'left downto d39_out1'left -7);
d40_out(7 downto 0) <= d40_out1(d40_out1'left downto d40_out1'left -7);
d41_out(7 downto 0) <= d41_out1(d41_out1'left downto d41_out1'left -7);
d42_out(7 downto 0) <= d42_out1(d42_out1'left downto d42_out1'left -7);
d43_out(7 downto 0) <= d43_out1(d43_out1'left downto d43_out1'left -7);
d44_out(7 downto 0) <= d44_out1(d44_out1'left downto d44_out1'left -7);
d45_out(7 downto 0) <= d45_out1(d45_out1'left downto d45_out1'left -7);
d46_out(7 downto 0) <= d46_out1(d46_out1'left downto d46_out1'left -7);
d47_out(7 downto 0) <= d47_out1(d47_out1'left downto d47_out1'left -7);
d48_out(7 downto 0) <= d48_out1(d48_out1'left downto d48_out1'left -7);
d49_out(7 downto 0) <= d49_out1(d49_out1'left downto d49_out1'left -7);
d50_out(7 downto 0) <= d50_out1(d50_out1'left downto d50_out1'left -7);
d51_out(7 downto 0) <= d51_out1(d51_out1'left downto d51_out1'left -7);
d52_out(7 downto 0) <= d52_out1(d52_out1'left downto d52_out1'left -7);
d53_out(7 downto 0) <= d53_out1(d53_out1'left downto d53_out1'left -7);
d54_out(7 downto 0) <= d54_out1(d54_out1'left downto d54_out1'left -7);
d55_out(7 downto 0) <= d55_out1(d55_out1'left downto d55_out1'left -7);
d56_out(7 downto 0) <= d56_out1(d56_out1'left downto d56_out1'left -7);
d57_out(7 downto 0) <= d57_out1(d57_out1'left downto d57_out1'left -7);
d58_out(7 downto 0) <= d58_out1(d58_out1'left downto d58_out1'left -7);
d59_out(7 downto 0) <= d59_out1(d59_out1'left downto d59_out1'left -7);
d60_out(7 downto 0) <= d60_out1(d60_out1'left downto d60_out1'left -7);
d61_out(7 downto 0) <= d61_out1(d61_out1'left downto d61_out1'left -7);
d62_out(7 downto 0) <= d62_out1(d62_out1'left downto d62_out1'left -7);
d63_out(7 downto 0) <= d63_out1(d63_out1'left downto d63_out1'left -7);
d64_out(7 downto 0) <= d64_out1(d64_out1'left downto d64_out1'left -7);

d65_out (7 downto 0) <= d65_out1 (d65_out1'left  downto d65_out1'left  -7);
d66_out (7 downto 0) <= d66_out1 (d66_out1'left  downto d66_out1'left  -7);
d67_out (7 downto 0) <= d67_out1 (d67_out1'left  downto d67_out1'left  -7);
d68_out (7 downto 0) <= d68_out1 (d68_out1'left  downto d68_out1'left  -7);
d69_out (7 downto 0) <= d69_out1 (d69_out1'left  downto d69_out1'left  -7);
d70_out (7 downto 0) <= d70_out1 (d70_out1'left  downto d70_out1'left  -7);
d71_out (7 downto 0) <= d71_out1 (d71_out1'left  downto d71_out1'left  -7);
d72_out (7 downto 0) <= d72_out1 (d72_out1'left  downto d72_out1'left  -7);
d73_out (7 downto 0) <= d73_out1 (d73_out1'left  downto d73_out1'left  -7);
d74_out (7 downto 0) <= d74_out1 (d74_out1'left  downto d74_out1'left  -7);
d75_out (7 downto 0) <= d75_out1 (d75_out1'left  downto d75_out1'left  -7);
d76_out (7 downto 0) <= d76_out1 (d76_out1'left  downto d76_out1'left  -7);
d77_out (7 downto 0) <= d77_out1 (d77_out1'left  downto d77_out1'left  -7);
d78_out (7 downto 0) <= d78_out1 (d78_out1'left  downto d78_out1'left  -7);
d79_out (7 downto 0) <= d79_out1 (d79_out1'left  downto d79_out1'left  -7);
d80_out (7 downto 0) <= d80_out1 (d80_out1'left  downto d80_out1'left  -7);
d81_out (7 downto 0) <= d81_out1 (d81_out1'left  downto d81_out1'left  -7);
d82_out (7 downto 0) <= d82_out1 (d82_out1'left  downto d82_out1'left  -7);
d83_out (7 downto 0) <= d83_out1 (d83_out1'left  downto d83_out1'left  -7);
d84_out (7 downto 0) <= d84_out1 (d84_out1'left  downto d84_out1'left  -7);
d85_out (7 downto 0) <= d85_out1 (d85_out1'left  downto d85_out1'left  -7);
d86_out (7 downto 0) <= d86_out1 (d86_out1'left  downto d86_out1'left  -7);
d87_out (7 downto 0) <= d87_out1 (d87_out1'left  downto d87_out1'left  -7);
d88_out (7 downto 0) <= d88_out1 (d88_out1'left  downto d88_out1'left  -7);
d89_out (7 downto 0) <= d89_out1 (d89_out1'left  downto d89_out1'left  -7);
d90_out (7 downto 0) <= d90_out1 (d90_out1'left  downto d90_out1'left  -7);
d91_out (7 downto 0) <= d91_out1 (d91_out1'left  downto d91_out1'left  -7);
d92_out (7 downto 0) <= d92_out1 (d92_out1'left  downto d92_out1'left  -7);
d93_out (7 downto 0) <= d93_out1 (d93_out1'left  downto d93_out1'left  -7);
d94_out (7 downto 0) <= d94_out1 (d94_out1'left  downto d94_out1'left  -7);
d95_out (7 downto 0) <= d95_out1 (d95_out1'left  downto d95_out1'left  -7);
d96_out (7 downto 0) <= d96_out1 (d96_out1'left  downto d96_out1'left  -7);
d97_out (7 downto 0) <= d97_out1 (d97_out1'left  downto d97_out1'left  -7);
d98_out (7 downto 0) <= d98_out1 (d98_out1'left  downto d98_out1'left  -7);
d99_out (7 downto 0) <= d99_out1 (d99_out1'left  downto d99_out1'left  -7);
d100_out(7 downto 0) <= d100_out1(d100_out1'left downto d100_out1'left -7);
d101_out(7 downto 0) <= d101_out1(d101_out1'left downto d101_out1'left -7);
d102_out(7 downto 0) <= d102_out1(d102_out1'left downto d102_out1'left -7);
d103_out(7 downto 0) <= d103_out1(d103_out1'left downto d103_out1'left -7);
d104_out(7 downto 0) <= d104_out1(d104_out1'left downto d104_out1'left -7);
d105_out(7 downto 0) <= d105_out1(d105_out1'left downto d105_out1'left -7);
d106_out(7 downto 0) <= d106_out1(d106_out1'left downto d106_out1'left -7);
d107_out(7 downto 0) <= d107_out1(d107_out1'left downto d107_out1'left -7);
d108_out(7 downto 0) <= d108_out1(d108_out1'left downto d108_out1'left -7);
d109_out(7 downto 0) <= d109_out1(d109_out1'left downto d109_out1'left -7);
d110_out(7 downto 0) <= d110_out1(d110_out1'left downto d110_out1'left -7);
d111_out(7 downto 0) <= d111_out1(d111_out1'left downto d111_out1'left -7);
d112_out(7 downto 0) <= d112_out1(d112_out1'left downto d112_out1'left -7);
d113_out(7 downto 0) <= d113_out1(d113_out1'left downto d113_out1'left -7);
d114_out(7 downto 0) <= d114_out1(d114_out1'left downto d114_out1'left -7);
d115_out(7 downto 0) <= d115_out1(d115_out1'left downto d115_out1'left -7);
d116_out(7 downto 0) <= d116_out1(d116_out1'left downto d116_out1'left -7);
d117_out(7 downto 0) <= d117_out1(d117_out1'left downto d117_out1'left -7);
d118_out(7 downto 0) <= d118_out1(d118_out1'left downto d118_out1'left -7);
d119_out(7 downto 0) <= d119_out1(d119_out1'left downto d119_out1'left -7);
d120_out(7 downto 0) <= d120_out1(d120_out1'left downto d120_out1'left -7);
d121_out(7 downto 0) <= d121_out1(d121_out1'left downto d121_out1'left -7);
d122_out(7 downto 0) <= d122_out1(d122_out1'left downto d122_out1'left -7);
d123_out(7 downto 0) <= d123_out1(d123_out1'left downto d123_out1'left -7);
d124_out(7 downto 0) <= d124_out1(d124_out1'left downto d124_out1'left -7);
d125_out(7 downto 0) <= d125_out1(d125_out1'left downto d125_out1'left -7);
d126_out(7 downto 0) <= d126_out1(d126_out1'left downto d126_out1'left -7);
d127_out(7 downto 0) <= d127_out1(d127_out1'left downto d127_out1'left -7);
d128_out(7 downto 0) <= d128_out1(d128_out1'left downto d128_out1'left -7);

  p_pca_weight : process (clk)
  begin
    if rising_edge(clk) then
       if pca_w_en = '1' then
          pca_mem(conv_integer('0' & pca_w_num)) <= pca_w_in;
       end if;
    end if;
  end process p_pca_weight;

pca_w01 <= pca_mem( 0);
pca_w02 <= pca_mem( 1);
pca_w03 <= pca_mem( 2);
pca_w04 <= pca_mem( 3);
pca_w05 <= pca_mem( 4);
pca_w06 <= pca_mem( 5);
pca_w07 <= pca_mem( 6);
pca_w08 <= pca_mem( 7);
pca_w09 <= pca_mem( 8);
pca_w10 <= pca_mem( 9);
pca_w11 <= pca_mem(10);
pca_w12 <= pca_mem(11);
pca_w13 <= pca_mem(12);
pca_w14 <= pca_mem(13);
pca_w15 <= pca_mem(14);
pca_w16 <= pca_mem(15);
pca_w17 <= pca_mem(16);
pca_w18 <= pca_mem(17);
pca_w19 <= pca_mem(18);
pca_w20 <= pca_mem(19);
pca_w21 <= pca_mem(20);
pca_w22 <= pca_mem(21);
pca_w23 <= pca_mem(22);
pca_w24 <= pca_mem(23);
pca_w25 <= pca_mem(24);
pca_w26 <= pca_mem(25);
pca_w27 <= pca_mem(26);
pca_w28 <= pca_mem(27);
pca_w29 <= pca_mem(28);
pca_w30 <= pca_mem(29);
pca_w31 <= pca_mem(30);
pca_w32 <= pca_mem(31);
pca_w33 <= pca_mem(32);
pca_w34 <= pca_mem(33);
pca_w35 <= pca_mem(34);
pca_w36 <= pca_mem(35);
pca_w37 <= pca_mem(36);
pca_w38 <= pca_mem(37);
pca_w39 <= pca_mem(38);
pca_w40 <= pca_mem(39);
pca_w41 <= pca_mem(40);
pca_w42 <= pca_mem(41);
pca_w43 <= pca_mem(42);
pca_w44 <= pca_mem(43);
pca_w45 <= pca_mem(44);
pca_w46 <= pca_mem(45);
pca_w47 <= pca_mem(46);
pca_w48 <= pca_mem(47);
pca_w49 <= pca_mem(48);
pca_w50 <= pca_mem(49);
pca_w51 <= pca_mem(50);
pca_w52 <= pca_mem(51);
pca_w53 <= pca_mem(52);
pca_w54 <= pca_mem(53);
pca_w55 <= pca_mem(54);
pca_w56 <= pca_mem(55);
pca_w57 <= pca_mem(56);
pca_w58 <= pca_mem(57);
pca_w59 <= pca_mem(58);
pca_w60 <= pca_mem(59);
pca_w61 <= pca_mem(60);
pca_w62 <= pca_mem(61);
pca_w63 <= pca_mem(62);
pca_w64 <= pca_mem(63);


pca_w65  <= pca_mem( 64);
pca_w66  <= pca_mem( 65);
pca_w67  <= pca_mem( 66);
pca_w68  <= pca_mem( 67);
pca_w69  <= pca_mem( 68);
pca_w70  <= pca_mem( 69);
pca_w71  <= pca_mem( 70);
pca_w72  <= pca_mem( 71);
pca_w73  <= pca_mem( 72);
pca_w74  <= pca_mem( 73);
pca_w75  <= pca_mem( 74);
pca_w76  <= pca_mem( 75);
pca_w77  <= pca_mem( 76);
pca_w78  <= pca_mem( 77);
pca_w79  <= pca_mem( 78);
pca_w80  <= pca_mem( 79);
pca_w81  <= pca_mem( 80);
pca_w82  <= pca_mem( 81);
pca_w83  <= pca_mem( 82);
pca_w84  <= pca_mem( 83);
pca_w85  <= pca_mem( 84);
pca_w86  <= pca_mem( 85);
pca_w87  <= pca_mem( 86);
pca_w88  <= pca_mem( 87);
pca_w89  <= pca_mem( 88);
pca_w90  <= pca_mem( 89);
pca_w91  <= pca_mem( 90);
pca_w92  <= pca_mem( 91);
pca_w93  <= pca_mem( 92);
pca_w94  <= pca_mem( 93);
pca_w95  <= pca_mem( 94);
pca_w96  <= pca_mem( 95);
pca_w97  <= pca_mem( 96);
pca_w98  <= pca_mem( 97);
pca_w99  <= pca_mem( 98);
pca_w100 <= pca_mem( 99);
pca_w101 <= pca_mem(100);
pca_w102 <= pca_mem(101);
pca_w103 <= pca_mem(102);
pca_w104 <= pca_mem(103);
pca_w105 <= pca_mem(104);
pca_w106 <= pca_mem(105);
pca_w107 <= pca_mem(106);
pca_w108 <= pca_mem(107);
pca_w109 <= pca_mem(108);
pca_w110 <= pca_mem(109);
pca_w111 <= pca_mem(110);
pca_w112 <= pca_mem(111);
pca_w113 <= pca_mem(112);
pca_w114 <= pca_mem(113);
pca_w115 <= pca_mem(114);
pca_w116 <= pca_mem(115);
pca_w117 <= pca_mem(116);
pca_w118 <= pca_mem(117);
pca_w119 <= pca_mem(118);
pca_w120 <= pca_mem(119);
pca_w121 <= pca_mem(120);
pca_w122 <= pca_mem(121);
pca_w123 <= pca_mem(122);
pca_w124 <= pca_mem(123);
pca_w125 <= pca_mem(124);
pca_w126 <= pca_mem(125);
pca_w127 <= pca_mem(126);
pca_w128 <= pca_mem(127);
g_PCA_en: if PCA_en = TRUE generate
--PCA32_1_inst: PCA_32 
--  generic map(
--           mult_sum => mult_sum,
--           N        => CL_W,
--           M        => PCAweightW,
--           in_row   => in_row,
--           in_col   => in_col
--           )
--  port map (
--           clk       => clk    ,
--           rst       => rst    ,
--d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, 
--d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
--d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, 
--d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
--
--           en_in     => cl_en_out,
--           sof_in    => cl_sof_out,
--
--           w01      => pca_w01, --x"d9", 
--           w02      => pca_w02, --x"66", 
--           w03      => pca_w03, --x"71", 
--           w04      => pca_w04, --x"f3", 
--           w05      => pca_w05, --x"12", 
--           w06      => pca_w06, --x"8e", 
--           w07      => pca_w07, --x"9c", 
--           w08      => pca_w08, --x"ab", 
--           w09      => pca_w09, --x"dc", 
--           w10      => pca_w10, --x"ec", 
--           w11      => pca_w11, --x"af", 
--           w12      => pca_w12, --x"b7", 
--           w13      => pca_w13, --x"67", 
--           w14      => pca_w14, --x"c9", 
--           w15      => pca_w15, --x"77", 
--           w16      => pca_w16, --x"5a", 
--           w17      => pca_w17, --x"45", 
--           w18      => pca_w18, --x"89", 
--           w19      => pca_w19, --x"a3", 
--           w20      => pca_w20, --x"0a", 
--           w21      => pca_w21, --x"9c", 
--           w22      => pca_w22, --x"c9", 
--           w23      => pca_w23, --x"65", 
--           w24      => pca_w24, --x"3d", 
--           w25      => pca_w25, --x"4c", 
--           w26      => pca_w26, --x"62", 
--           w27      => pca_w27, --x"2f", 
--           w28      => pca_w28, --x"66", 
--           w29      => pca_w29, --x"4b", 
--           w30      => pca_w30, --x"f3", 
--           w31      => pca_w31, --x"a1", 
--           w32      => pca_w32, --x"ba", 
--
--           d_out   => pca_d01_out   ,
--           en_out  => pca_en_out  ,
--           sof_out => pca_sof_out );


--PCA64_1_inst: PCA_128 
--  generic map(
--           mult_sum => mult_sum,
--           N        => CL_W,
--           M        => PCAweightW,
--           in_row   => in_row,
--           in_col   => in_col
--           )
--  port map (
--           clk       => clk    ,
--           rst       => rst    ,
--d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, 
--d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
--d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, 
--d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
--d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, 
--d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
--d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,
--d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
--           en_in     => cl_en_out,
--           sof_in    => cl_sof_out,
--
--           w01      => pca_w01, --x"d9", 
--           w02      => pca_w02, --x"66", 
--           w03      => pca_w03, --x"71", 
--           w04      => pca_w04, --x"f3", 
--           w05      => pca_w05, --x"12", 
--           w06      => pca_w06, --x"8e", 
--           w07      => pca_w07, --x"9c", 
--           w08      => pca_w08, --x"ab", 
--           w09      => pca_w09, --x"dc", 
--           w10      => pca_w10, --x"ec", 
--           w11      => pca_w11, --x"af", 
--           w12      => pca_w12, --x"b7", 
--           w13      => pca_w13, --x"67", 
--           w14      => pca_w14, --x"c9", 
--           w15      => pca_w15, --x"77", 
--           w16      => pca_w16, --x"5a", 
--           w17      => pca_w17, --x"45", 
--           w18      => pca_w18, --x"89", 
--           w19      => pca_w19, --x"a3", 
--           w20      => pca_w20, --x"0a", 
--           w21      => pca_w21, --x"9c", 
--           w22      => pca_w22, --x"c9", 
--           w23      => pca_w23, --x"65", 
--           w24      => pca_w24, --x"3d", 
--           w25      => pca_w25, --x"4c", 
--           w26      => pca_w26, --x"62", 
--           w27      => pca_w27, --x"2f", 
--           w28      => pca_w28, --x"66", 
--           w29      => pca_w29, --x"4b", 
--           w30      => pca_w30, --x"f3", 
--           w31      => pca_w31, --x"a1", 
--           w32      => pca_w32, --x"ba", 
--           w33      => pca_w33, --x"38", 
--           w34      => pca_w34, --x"89", 
--           w35      => pca_w35, --x"30", 
--           w36      => pca_w36, --x"e0", 
--           w37      => pca_w37, --x"91", 
--           w38      => pca_w38, --x"e0", 
--           w39      => pca_w39, --x"69", 
--           w40      => pca_w40, --x"f8", 
--           w41      => pca_w41, --x"2f", 
--           w42      => pca_w42, --x"10", 
--           w43      => pca_w43, --x"a2", 
--           w44      => pca_w44, --x"ab", 
--           w45      => pca_w45, --x"de", 
--           w46      => pca_w46, --x"6f", 
--           w47      => pca_w47, --x"25", 
--           w48      => pca_w48, --x"a8", 
--           w49      => pca_w49, --x"b4", 
--           w50      => pca_w50, --x"89", 
--           w51      => pca_w51, --x"de", 
--           w52      => pca_w52, --x"5f", 
--           w53      => pca_w53, --x"c2", 
--           w54      => pca_w54, --x"ad", 
--           w55      => pca_w55, --x"d7", 
--           w56      => pca_w56, --x"fc", 
--           w57      => pca_w57, --x"ce", 
--           w58      => pca_w58, --x"4a", 
--           w59      => pca_w59, --x"0b", 
--           w60      => pca_w60, --x"dd", 
--           w61      => pca_w61, --x"d3", 
--           w62      => pca_w62, --x"0f", 
--           w63      => pca_w63, --x"80", 
--           w64      => pca_w64, --x"90", 
--
--           d_out   => pca_d01_out   ,
--           en_out  => pca_en_out  ,
--           sof_out => pca_sof_out );


--PCA128_1_inst: PCA_128 
--  generic map(
--           mult_sum => mult_sum,
--           N        => CL_W,
--           M        => PCAweightW,
--           in_row   => in_row,
--           in_col   => in_col
--           )
--  port map (
--           clk       => clk    ,
--           rst       => rst    ,
--d01_in   => d01_out, d02_in    => d02_out, d03_in  => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in   => d08_out, 
--d09_in   => d09_out, d10_in    => d10_out, d11_in  => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in   => d16_out, 
--d17_in   => d17_out, d18_in    => d18_out, d19_in  => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in   => d24_out, 
--d25_in   => d25_out, d26_in    => d26_out, d27_in  => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in   => d32_out, 
--d33_in   => d33_out, d34_in    => d34_out, d35_in  => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in   => d40_out, 
--d41_in   => d41_out, d42_in    => d42_out, d43_in  => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in   => d48_out, 
--d49_in   => d49_out, d50_in    => d50_out, d51_in  => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in   => d56_out,
--d57_in   => d57_out, d58_in    => d58_out, d59_in  => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in   => d64_out, 
--
--d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, 
--d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
--d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, 
--d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
--d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,
--d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
--d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,
--d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
--           en_in     => cl_en_out,
--           sof_in    => cl_sof_out,
--
--w01 => Pw(59)(     7 downto    0), w02 => Pw(59)( 2*8-1 downto    8), w03 => Pw(59)( 3*8-1 downto  2*8), w04 => Pw(59)( 4*8-1 downto  3*8), w05 => Pw(59)( 5*8-1 downto  4*8), w06 => Pw(59)( 6*8-1 downto  5*8), w07 => Pw(59)( 7*8-1 downto  6*8), w08 => Pw(59)( 8*8-1 downto  7*8),  
--w09 => Pw(59)( 9*8-1 downto  8*8), w10 => Pw(59)(10*8-1 downto  9*8), w11 => Pw(59)(11*8-1 downto 10*8), w12 => Pw(59)(12*8-1 downto 11*8), w13 => Pw(59)(13*8-1 downto 12*8), w14 => Pw(59)(14*8-1 downto 13*8), w15 => Pw(59)(15*8-1 downto 14*8), w16 => Pw(59)(16*8-1 downto 15*8),  
--w17 => Pw(59)(17*8-1 downto 16*8), w18 => Pw(59)(18*8-1 downto 17*8), w19 => Pw(59)(19*8-1 downto 18*8), w20 => Pw(59)(20*8-1 downto 19*8), w21 => Pw(59)(21*8-1 downto 20*8), w22 => Pw(59)(22*8-1 downto 21*8), w23 => Pw(59)(23*8-1 downto 22*8), w24 => Pw(59)(24*8-1 downto 23*8),  
--w25 => Pw(59)(25*8-1 downto 24*8), w26 => Pw(59)(26*8-1 downto 25*8), w27 => Pw(59)(27*8-1 downto 26*8), w28 => Pw(59)(28*8-1 downto 27*8), w29 => Pw(59)(29*8-1 downto 28*8), w30 => Pw(59)(30*8-1 downto 29*8), w31 => Pw(59)(31*8-1 downto 30*8), w32 => Pw(59)(32*8-1 downto 31*8),  
--w33 => Pw(59)(33*8-1 downto 32*8), w34 => Pw(59)(34*8-1 downto 33*8), w35 => Pw(59)(35*8-1 downto 34*8), w36 => Pw(59)(36*8-1 downto 35*8), w37 => Pw(59)(37*8-1 downto 36*8), w38 => Pw(59)(38*8-1 downto 37*8), w39 => Pw(59)(39*8-1 downto 38*8), w40 => Pw(59)(40*8-1 downto 39*8),  
--w41 => Pw(59)(41*8-1 downto 40*8), w42 => Pw(59)(42*8-1 downto 41*8), w43 => Pw(59)(43*8-1 downto 42*8), w44 => Pw(59)(44*8-1 downto 43*8), w45 => Pw(59)(45*8-1 downto 44*8), w46 => Pw(59)(46*8-1 downto 45*8), w47 => Pw(59)(47*8-1 downto 46*8), w48 => Pw(59)(48*8-1 downto 47*8),  
--w49 => Pw(59)(49*8-1 downto 48*8), w50 => Pw(59)(50*8-1 downto 49*8), w51 => Pw(59)(51*8-1 downto 50*8), w52 => Pw(59)(52*8-1 downto 51*8), w53 => Pw(59)(53*8-1 downto 52*8), w54 => Pw(59)(54*8-1 downto 53*8), w55 => Pw(59)(55*8-1 downto 54*8), w56 => Pw(59)(56*8-1 downto 55*8),  
--w57 => Pw(59)(57*8-1 downto 56*8), w58 => Pw(59)(58*8-1 downto 57*8), w59 => Pw(59)(59*8-1 downto 58*8), w60 => Pw(59)(60*8-1 downto 59*8), w61 => Pw(59)(61*8-1 downto 60*8), w62 => Pw(59)(62*8-1 downto 61*8), w63 => Pw(59)(63*8-1 downto 62*8), w64 => Pw(59)(64*8-1 downto 63*8), 
--
--w65 => Pw()(*8-1 downto *8), w66 => Pw()(*8-1 downto *8), w67 => Pw()(*8-1 downto *8), w68 => Pw()(*8-1 downto *8), w69 => Pw()(*8-1 downto *8), w70 => Pw()(*8-1 downto *8), w71 => Pw()(*8-1 downto *8), w72 => Pw()(*8-1 downto *8), 
--w73 => Pw()(*8-1 downto *8), w74 => Pw()(*8-1 downto *8), w75 => Pw()(*8-1 downto *8), w76 => Pw()(*8-1 downto *8), w77 => Pw()(*8-1 downto *8), w78 => Pw()(*8-1 downto *8), w79 => Pw()(*8-1 downto *8), w80 => Pw()(*8-1 downto *8), 
--w81 => Pw()(*8-1 downto *8), w82 => Pw()(*8-1 downto *8), w83 => Pw()(*8-1 downto *8), w84 => Pw()(*8-1 downto *8), w85 => Pw()(*8-1 downto *8), w86 => Pw()(*8-1 downto *8), w87 => Pw()(*8-1 downto *8), w88 => Pw()(*8-1 downto *8), 
--w89 => Pw()(*8-1 downto *8), w90 => Pw()(*8-1 downto *8), w91 => Pw()(*8-1 downto *8), w92 => Pw()(*8-1 downto *8), w93 => Pw()(*8-1 downto *8), w94 => Pw()(*8-1 downto *8), w95 => Pw()(*8-1 downto *8), w96 => Pw()(*8-1 downto *8), 
--w97 => Pw()(*8-1 downto *8), w98 => Pw()(*8-1 downto *8), w99 => Pw()(*8-1 downto *8), w100=> Pw()(*8-1 downto *8), w101=> Pw()(*8-1 downto *8), w102=> Pw()(*8-1 downto *8), w103=> Pw()(*8-1 downto *8), w104=> Pw()(*8-1 downto *8), 
--w105=> Pw()(*8-1 downto *8), w106=> Pw()(*8-1 downto *8), w107=> Pw()(*8-1 downto *8), w108=> Pw()(*8-1 downto *8), w109=> Pw()(*8-1 downto *8), w110=> Pw()(*8-1 downto *8), w111=> Pw()(*8-1 downto *8), w112=> Pw()(*8-1 downto *8), 
--w113=> Pw()(*8-1 downto *8), w114=> Pw()(*8-1 downto *8), w115=> Pw()(*8-1 downto *8), w116=> Pw()(*8-1 downto *8), w117=> Pw()(*8-1 downto *8), w118=> Pw()(*8-1 downto *8), w119=> Pw()(*8-1 downto *8), w120=> Pw()(*8-1 downto *8), 
--w121=> Pw()(*8-1 downto *8), w122=> Pw()(*8-1 downto *8), w123=> Pw()(*8-1 downto *8), w124=> Pw()(*8-1 downto *8), w125=> Pw()(*8-1 downto *8), w126=> Pw()(*8-1 downto *8), w127=> Pw()(*8-1 downto *8), w128=> Pw()(*8-1 downto *8), 
--           d_out   => pca_d01_out   ,
--           en_out  => pca_en_out  ,
--           sof_out => pca_sof_out );


PCA128_1_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 

d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 1)(     7 downto    0), w02 => Pw( 1)( 2*8-1 downto    8), w03 => Pw( 1)( 3*8-1 downto  2*8), w04 => Pw( 1)( 4*8-1 downto  3*8), w05 => Pw( 1)( 5*8-1 downto  4*8), w06 => Pw( 1)( 6*8-1 downto  5*8), w07 => Pw( 1)( 7*8-1 downto  6*8), w08 => Pw( 1)( 8*8-1 downto  7*8),  w09 => Pw( 1)( 9*8-1 downto  8*8), w10 => Pw( 1)(10*8-1 downto  9*8), w11 => Pw( 1)(11*8-1 downto 10*8), w12 => Pw( 1)(12*8-1 downto 11*8), w13 => Pw( 1)(13*8-1 downto 12*8), w14 => Pw( 1)(14*8-1 downto 13*8), w15 => Pw( 1)(15*8-1 downto 14*8), w16 => Pw( 1)(16*8-1 downto 15*8),  
w17 => Pw( 1)(17*8-1 downto 16*8), w18 => Pw( 1)(18*8-1 downto 17*8), w19 => Pw( 1)(19*8-1 downto 18*8), w20 => Pw( 1)(20*8-1 downto 19*8), w21 => Pw( 1)(21*8-1 downto 20*8), w22 => Pw( 1)(22*8-1 downto 21*8), w23 => Pw( 1)(23*8-1 downto 22*8), w24 => Pw( 1)(24*8-1 downto 23*8),  w25 => Pw( 1)(25*8-1 downto 24*8), w26 => Pw( 1)(26*8-1 downto 25*8), w27 => Pw( 1)(27*8-1 downto 26*8), w28 => Pw( 1)(28*8-1 downto 27*8), w29 => Pw( 1)(29*8-1 downto 28*8), w30 => Pw( 1)(30*8-1 downto 29*8), w31 => Pw( 1)(31*8-1 downto 30*8), w32 => Pw( 1)(32*8-1 downto 31*8),  
w33 => Pw( 1)(33*8-1 downto 32*8), w34 => Pw( 1)(34*8-1 downto 33*8), w35 => Pw( 1)(35*8-1 downto 34*8), w36 => Pw( 1)(36*8-1 downto 35*8), w37 => Pw( 1)(37*8-1 downto 36*8), w38 => Pw( 1)(38*8-1 downto 37*8), w39 => Pw( 1)(39*8-1 downto 38*8), w40 => Pw( 1)(40*8-1 downto 39*8),  w41 => Pw( 1)(41*8-1 downto 40*8), w42 => Pw( 1)(42*8-1 downto 41*8), w43 => Pw( 1)(43*8-1 downto 42*8), w44 => Pw( 1)(44*8-1 downto 43*8), w45 => Pw( 1)(45*8-1 downto 44*8), w46 => Pw( 1)(46*8-1 downto 45*8), w47 => Pw( 1)(47*8-1 downto 46*8), w48 => Pw( 1)(48*8-1 downto 47*8),  
w49 => Pw( 1)(49*8-1 downto 48*8), w50 => Pw( 1)(50*8-1 downto 49*8), w51 => Pw( 1)(51*8-1 downto 50*8), w52 => Pw( 1)(52*8-1 downto 51*8), w53 => Pw( 1)(53*8-1 downto 52*8), w54 => Pw( 1)(54*8-1 downto 53*8), w55 => Pw( 1)(55*8-1 downto 54*8), w56 => Pw( 1)(56*8-1 downto 55*8),  w57 => Pw( 1)(57*8-1 downto 56*8), w58 => Pw( 1)(58*8-1 downto 57*8), w59 => Pw( 1)(59*8-1 downto 58*8), w60 => Pw( 1)(60*8-1 downto 59*8), w61 => Pw( 1)(61*8-1 downto 60*8), w62 => Pw( 1)(62*8-1 downto 61*8), w63 => Pw( 1)(63*8-1 downto 62*8), w64 => Pw( 1)(64*8-1 downto 63*8),  

w65 => Pw(1)( 65*8-1 downto  64*8), w66 => Pw(1)( 66*8-1 downto  65*8), w67 => Pw(1)( 67*8-1 downto  66*8), w68 => Pw(1)( 68*8-1 downto  67*8), w69 => Pw(1)( 69*8-1 downto  68*8), w70 => Pw(1)( 70*8-1 downto  69*8), w71 => Pw(1)( 71*8-1 downto  70*8), w72 => Pw(1)( 72*8-1 downto  71*8), w73 => Pw(1)( 73*8-1 downto  72*8), w74 => Pw(1)( 74*8-1 downto  73*8), w75 => Pw(1)( 75*8-1 downto  74*8), w76 => Pw(1)( 76*8-1 downto  75*8), w77 => Pw(1)( 77*8-1 downto  76*8), w78 => Pw(1)( 78*8-1 downto  77*8), w79 => Pw(1)( 79*8-1 downto  78*8), w80 => Pw(1)( 80*8-1 downto  79*8), 
w81 => Pw(1)( 81*8-1 downto  80*8), w82 => Pw(1)( 82*8-1 downto  81*8), w83 => Pw(1)( 83*8-1 downto  82*8), w84 => Pw(1)( 84*8-1 downto  83*8), w85 => Pw(1)( 85*8-1 downto  84*8), w86 => Pw(1)( 86*8-1 downto  85*8), w87 => Pw(1)( 87*8-1 downto  86*8), w88 => Pw(1)( 88*8-1 downto  87*8), w89 => Pw(1)( 89*8-1 downto  88*8), w90 => Pw(1)( 90*8-1 downto  89*8), w91 => Pw(1)( 91*8-1 downto  90*8), w92 => Pw(1)( 92*8-1 downto  91*8), w93 => Pw(1)( 93*8-1 downto  92*8), w94 => Pw(1)( 94*8-1 downto  93*8), w95 => Pw(1)( 95*8-1 downto  94*8), w96 => Pw(1)( 96*8-1 downto  95*8), 
w97 => Pw(1)( 97*8-1 downto  96*8), w98 => Pw(1)( 98*8-1 downto  97*8), w99 => Pw(1)( 99*8-1 downto  98*8), w100=> Pw(1)(100*8-1 downto  99*8), w101=> Pw(1)(101*8-1 downto 100*8), w102=> Pw(1)(102*8-1 downto 101*8), w103=> Pw(1)(103*8-1 downto 102*8), w104=> Pw(1)(104*8-1 downto 103*8), w105=> Pw(1)(105*8-1 downto 104*8), w106=> Pw(1)(106*8-1 downto 105*8), w107=> Pw(1)(107*8-1 downto 106*8), w108=> Pw(1)(108*8-1 downto 107*8), w109=> Pw(1)(109*8-1 downto 108*8), w110=> Pw(1)(110*8-1 downto 109*8), w111=> Pw(1)(111*8-1 downto 110*8), w112=> Pw(1)(112*8-1 downto 111*8), 
w113=> Pw(1)(113*8-1 downto 112*8), w114=> Pw(1)(114*8-1 downto 113*8), w115=> Pw(1)(115*8-1 downto 114*8), w116=> Pw(1)(116*8-1 downto 115*8), w117=> Pw(1)(117*8-1 downto 116*8), w118=> Pw(1)(118*8-1 downto 117*8), w119=> Pw(1)(119*8-1 downto 118*8), w120=> Pw(1)(120*8-1 downto 119*8), w121=> Pw(1)(121*8-1 downto 120*8), w122=> Pw(1)(122*8-1 downto 121*8), w123=> Pw(1)(123*8-1 downto 122*8), w124=> Pw(1)(124*8-1 downto 123*8), w125=> Pw(1)(125*8-1 downto 124*8), w126=> Pw(1)(126*8-1 downto 125*8), w127=> Pw(1)(127*8-1 downto 126*8), w128=> Pw(1)(128*8-1 downto 127*8), 

--w65 => Pw()( 65*8-1 downto  64*8), w66 => Pw()( 66*8-1 downto  65*8), w67 => Pw()( 67*8-1 downto  66*8), w68 => Pw()( 68*8-1 downto  67*8), w69 => Pw()( 69*8-1 downto  68*8), w70 => Pw()( 70*8-1 downto  69*8), w71 => Pw()( 71*8-1 downto  70*8), w72 => Pw()( 72*8-1 downto  71*8), 
--w73 => Pw()( 73*8-1 downto  72*8), w74 => Pw()( 74*8-1 downto  73*8), w75 => Pw()( 75*8-1 downto  74*8), w76 => Pw()( 76*8-1 downto  75*8), w77 => Pw()( 77*8-1 downto  76*8), w78 => Pw()( 78*8-1 downto  77*8), w79 => Pw()( 79*8-1 downto  78*8), w80 => Pw()( 80*8-1 downto  79*8), 
--w81 => Pw()( 81*8-1 downto  80*8), w82 => Pw()( 82*8-1 downto  81*8), w83 => Pw()( 83*8-1 downto  82*8), w84 => Pw()( 84*8-1 downto  83*8), w85 => Pw()( 85*8-1 downto  84*8), w86 => Pw()( 86*8-1 downto  85*8), w87 => Pw()( 87*8-1 downto  86*8), w88 => Pw()( 88*8-1 downto  87*8), 
--w89 => Pw()( 89*8-1 downto  88*8), w90 => Pw()( 90*8-1 downto  89*8), w91 => Pw()( 91*8-1 downto  90*8), w92 => Pw()( 92*8-1 downto  91*8), w93 => Pw()( 93*8-1 downto  92*8), w94 => Pw()( 94*8-1 downto  93*8), w95 => Pw()( 95*8-1 downto  94*8), w96 => Pw()( 96*8-1 downto  95*8), 
--w97 => Pw()( 97*8-1 downto  96*8), w98 => Pw()( 98*8-1 downto  97*8), w99 => Pw()( 99*8-1 downto  98*8), w100=> Pw()(100*8-1 downto  99*8), w101=> Pw()(101*8-1 downto 100*8), w102=> Pw()(102*8-1 downto 101*8), w103=> Pw()(103*8-1 downto 102*8), w104=> Pw()(104*8-1 downto 103*8), 
--w105=> Pw()(105*8-1 downto 104*8), w106=> Pw()(106*8-1 downto 105*8), w107=> Pw()(107*8-1 downto 106*8), w108=> Pw()(108*8-1 downto 107*8), w109=> Pw()(109*8-1 downto 108*8), w110=> Pw()(110*8-1 downto 109*8), w111=> Pw()(111*8-1 downto 110*8), w112=> Pw()(112*8-1 downto 111*8), 
--w113=> Pw()(113*8-1 downto 112*8), w114=> Pw()(114*8-1 downto 113*8), w115=> Pw()(115*8-1 downto 114*8), w116=> Pw()(116*8-1 downto 115*8), w117=> Pw()(117*8-1 downto 116*8), w118=> Pw()(118*8-1 downto 117*8), w119=> Pw()(119*8-1 downto 118*8), w120=> Pw()(120*8-1 downto 119*8), 
--w121=> Pw()(121*8-1 downto 120*8), w122=> Pw()(122*8-1 downto 121*8), w123=> Pw()(123*8-1 downto 122*8), w124=> Pw()(124*8-1 downto 123*8), w125=> Pw()(125*8-1 downto 124*8), w126=> Pw()(126*8-1 downto 125*8), w127=> Pw()(127*8-1 downto 126*8), w128=> Pw()(128*8-1 downto 127*8), 
           d_out   => pca_d01_out   ,
           en_out  => pca_en_out  ,
           sof_out => open );


PCA128_2_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 2)(     7 downto    0), w02 => Pw( 2)( 2*8-1 downto    8), w03 => Pw( 2)( 3*8-1 downto  2*8), w04 => Pw( 2)( 4*8-1 downto  3*8), w05 => Pw( 2)( 5*8-1 downto  4*8), w06 => Pw( 2)( 6*8-1 downto  5*8), w07 => Pw( 2)( 7*8-1 downto  6*8), w08 => Pw( 2)( 8*8-1 downto  7*8),  
w09 => Pw( 2)( 9*8-1 downto  8*8), w10 => Pw( 2)(10*8-1 downto  9*8), w11 => Pw( 2)(11*8-1 downto 10*8), w12 => Pw( 2)(12*8-1 downto 11*8), w13 => Pw( 2)(13*8-1 downto 12*8), w14 => Pw( 2)(14*8-1 downto 13*8), w15 => Pw( 2)(15*8-1 downto 14*8), w16 => Pw( 2)(16*8-1 downto 15*8),  
w17 => Pw( 2)(17*8-1 downto 16*8), w18 => Pw( 2)(18*8-1 downto 17*8), w19 => Pw( 2)(19*8-1 downto 18*8), w20 => Pw( 2)(20*8-1 downto 19*8), w21 => Pw( 2)(21*8-1 downto 20*8), w22 => Pw( 2)(22*8-1 downto 21*8), w23 => Pw( 2)(23*8-1 downto 22*8), w24 => Pw( 2)(24*8-1 downto 23*8),  
w25 => Pw( 2)(25*8-1 downto 24*8), w26 => Pw( 2)(26*8-1 downto 25*8), w27 => Pw( 2)(27*8-1 downto 26*8), w28 => Pw( 2)(28*8-1 downto 27*8), w29 => Pw( 2)(29*8-1 downto 28*8), w30 => Pw( 2)(30*8-1 downto 29*8), w31 => Pw( 2)(31*8-1 downto 30*8), w32 => Pw( 2)(32*8-1 downto 31*8),  
w33 => Pw( 2)(33*8-1 downto 32*8), w34 => Pw( 2)(34*8-1 downto 33*8), w35 => Pw( 2)(35*8-1 downto 34*8), w36 => Pw( 2)(36*8-1 downto 35*8), w37 => Pw( 2)(37*8-1 downto 36*8), w38 => Pw( 2)(38*8-1 downto 37*8), w39 => Pw( 2)(39*8-1 downto 38*8), w40 => Pw( 2)(40*8-1 downto 39*8),  
w41 => Pw( 2)(41*8-1 downto 40*8), w42 => Pw( 2)(42*8-1 downto 41*8), w43 => Pw( 2)(43*8-1 downto 42*8), w44 => Pw( 2)(44*8-1 downto 43*8), w45 => Pw( 2)(45*8-1 downto 44*8), w46 => Pw( 2)(46*8-1 downto 45*8), w47 => Pw( 2)(47*8-1 downto 46*8), w48 => Pw( 2)(48*8-1 downto 47*8),  
w49 => Pw( 2)(49*8-1 downto 48*8), w50 => Pw( 2)(50*8-1 downto 49*8), w51 => Pw( 2)(51*8-1 downto 50*8), w52 => Pw( 2)(52*8-1 downto 51*8), w53 => Pw( 2)(53*8-1 downto 52*8), w54 => Pw( 2)(54*8-1 downto 53*8), w55 => Pw( 2)(55*8-1 downto 54*8), w56 => Pw( 2)(56*8-1 downto 55*8),  
w57 => Pw( 2)(57*8-1 downto 56*8), w58 => Pw( 2)(58*8-1 downto 57*8), w59 => Pw( 2)(59*8-1 downto 58*8), w60 => Pw( 2)(60*8-1 downto 59*8), w61 => Pw( 2)(61*8-1 downto 60*8), w62 => Pw( 2)(62*8-1 downto 61*8), w63 => Pw( 2)(63*8-1 downto 62*8), w64 => Pw( 2)(64*8-1 downto 63*8), 
w65 => Pw(2)( 65*8-1 downto  64*8), w66 => Pw(2)( 66*8-1 downto  65*8), w67 => Pw(2)( 67*8-1 downto  66*8), w68 => Pw(2)( 68*8-1 downto  67*8), w69 => Pw(2)( 69*8-1 downto  68*8), w70 => Pw(2)( 70*8-1 downto  69*8), w71 => Pw(2)( 71*8-1 downto  70*8), w72 => Pw(2)( 72*8-1 downto  71*8), 
w73 => Pw(2)( 73*8-1 downto  72*8), w74 => Pw(2)( 74*8-1 downto  73*8), w75 => Pw(2)( 75*8-1 downto  74*8), w76 => Pw(2)( 76*8-1 downto  75*8), w77 => Pw(2)( 77*8-1 downto  76*8), w78 => Pw(2)( 78*8-1 downto  77*8), w79 => Pw(2)( 79*8-1 downto  78*8), w80 => Pw(2)( 80*8-1 downto  79*8), 
w81 => Pw(2)( 81*8-1 downto  80*8), w82 => Pw(2)( 82*8-1 downto  81*8), w83 => Pw(2)( 83*8-1 downto  82*8), w84 => Pw(2)( 84*8-1 downto  83*8), w85 => Pw(2)( 85*8-1 downto  84*8), w86 => Pw(2)( 86*8-1 downto  85*8), w87 => Pw(2)( 87*8-1 downto  86*8), w88 => Pw(2)( 88*8-1 downto  87*8), 
w89 => Pw(2)( 89*8-1 downto  88*8), w90 => Pw(2)( 90*8-1 downto  89*8), w91 => Pw(2)( 91*8-1 downto  90*8), w92 => Pw(2)( 92*8-1 downto  91*8), w93 => Pw(2)( 93*8-1 downto  92*8), w94 => Pw(2)( 94*8-1 downto  93*8), w95 => Pw(2)( 95*8-1 downto  94*8), w96 => Pw(2)( 96*8-1 downto  95*8), 
w97 => Pw(2)( 97*8-1 downto  96*8), w98 => Pw(2)( 98*8-1 downto  97*8), w99 => Pw(2)( 99*8-1 downto  98*8), w100=> Pw(2)(100*8-1 downto  99*8), w101=> Pw(2)(101*8-1 downto 100*8), w102=> Pw(2)(102*8-1 downto 101*8), w103=> Pw(2)(103*8-1 downto 102*8), w104=> Pw(2)(104*8-1 downto 103*8), 
w105=> Pw(2)(105*8-1 downto 104*8), w106=> Pw(2)(106*8-1 downto 105*8), w107=> Pw(2)(107*8-1 downto 106*8), w108=> Pw(2)(108*8-1 downto 107*8), w109=> Pw(2)(109*8-1 downto 108*8), w110=> Pw(2)(110*8-1 downto 109*8), w111=> Pw(2)(111*8-1 downto 110*8), w112=> Pw(2)(112*8-1 downto 111*8), 
w113=> Pw(2)(113*8-1 downto 112*8), w114=> Pw(2)(114*8-1 downto 113*8), w115=> Pw(2)(115*8-1 downto 114*8), w116=> Pw(2)(116*8-1 downto 115*8), w117=> Pw(2)(117*8-1 downto 116*8), w118=> Pw(2)(118*8-1 downto 117*8), w119=> Pw(2)(119*8-1 downto 118*8), w120=> Pw(2)(120*8-1 downto 119*8), 
w121=> Pw(2)(121*8-1 downto 120*8), w122=> Pw(2)(122*8-1 downto 121*8), w123=> Pw(2)(123*8-1 downto 122*8), w124=> Pw(2)(124*8-1 downto 123*8), w125=> Pw(2)(125*8-1 downto 124*8), w126=> Pw(2)(126*8-1 downto 125*8), w127=> Pw(2)(127*8-1 downto 126*8), w128=> Pw(2)(128*8-1 downto 127*8), 

           d_out   => pca_d02_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_3_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 3)(     7 downto    0), w02 => Pw( 3)( 2*8-1 downto    8), w03 => Pw( 3)( 3*8-1 downto  2*8), w04 => Pw( 3)( 4*8-1 downto  3*8), w05 => Pw( 3)( 5*8-1 downto  4*8), w06 => Pw( 3)( 6*8-1 downto  5*8), w07 => Pw( 3)( 7*8-1 downto  6*8), w08 => Pw( 3)( 8*8-1 downto  7*8),  
w09 => Pw( 3)( 9*8-1 downto  8*8), w10 => Pw( 3)(10*8-1 downto  9*8), w11 => Pw( 3)(11*8-1 downto 10*8), w12 => Pw( 3)(12*8-1 downto 11*8), w13 => Pw( 3)(13*8-1 downto 12*8), w14 => Pw( 3)(14*8-1 downto 13*8), w15 => Pw( 3)(15*8-1 downto 14*8), w16 => Pw( 3)(16*8-1 downto 15*8),  
w17 => Pw( 3)(17*8-1 downto 16*8), w18 => Pw( 3)(18*8-1 downto 17*8), w19 => Pw( 3)(19*8-1 downto 18*8), w20 => Pw( 3)(20*8-1 downto 19*8), w21 => Pw( 3)(21*8-1 downto 20*8), w22 => Pw( 3)(22*8-1 downto 21*8), w23 => Pw( 3)(23*8-1 downto 22*8), w24 => Pw( 3)(24*8-1 downto 23*8),  
w25 => Pw( 3)(25*8-1 downto 24*8), w26 => Pw( 3)(26*8-1 downto 25*8), w27 => Pw( 3)(27*8-1 downto 26*8), w28 => Pw( 3)(28*8-1 downto 27*8), w29 => Pw( 3)(29*8-1 downto 28*8), w30 => Pw( 3)(30*8-1 downto 29*8), w31 => Pw( 3)(31*8-1 downto 30*8), w32 => Pw( 3)(32*8-1 downto 31*8),  
w33 => Pw( 3)(33*8-1 downto 32*8), w34 => Pw( 3)(34*8-1 downto 33*8), w35 => Pw( 3)(35*8-1 downto 34*8), w36 => Pw( 3)(36*8-1 downto 35*8), w37 => Pw( 3)(37*8-1 downto 36*8), w38 => Pw( 3)(38*8-1 downto 37*8), w39 => Pw( 3)(39*8-1 downto 38*8), w40 => Pw( 3)(40*8-1 downto 39*8),  
w41 => Pw( 3)(41*8-1 downto 40*8), w42 => Pw( 3)(42*8-1 downto 41*8), w43 => Pw( 3)(43*8-1 downto 42*8), w44 => Pw( 3)(44*8-1 downto 43*8), w45 => Pw( 3)(45*8-1 downto 44*8), w46 => Pw( 3)(46*8-1 downto 45*8), w47 => Pw( 3)(47*8-1 downto 46*8), w48 => Pw( 3)(48*8-1 downto 47*8),  
w49 => Pw( 3)(49*8-1 downto 48*8), w50 => Pw( 3)(50*8-1 downto 49*8), w51 => Pw( 3)(51*8-1 downto 50*8), w52 => Pw( 3)(52*8-1 downto 51*8), w53 => Pw( 3)(53*8-1 downto 52*8), w54 => Pw( 3)(54*8-1 downto 53*8), w55 => Pw( 3)(55*8-1 downto 54*8), w56 => Pw( 3)(56*8-1 downto 55*8),  
w57 => Pw( 3)(57*8-1 downto 56*8), w58 => Pw( 3)(58*8-1 downto 57*8), w59 => Pw( 3)(59*8-1 downto 58*8), w60 => Pw( 3)(60*8-1 downto 59*8), w61 => Pw( 3)(61*8-1 downto 60*8), w62 => Pw( 3)(62*8-1 downto 61*8), w63 => Pw( 3)(63*8-1 downto 62*8), w64 => Pw( 3)(64*8-1 downto 63*8), 
w65 => Pw(3)( 65*8-1 downto  64*8), w66 => Pw(3)( 66*8-1 downto  65*8), w67 => Pw(3)( 67*8-1 downto  66*8), w68 => Pw(3)( 68*8-1 downto  67*8), w69 => Pw(3)( 69*8-1 downto  68*8), w70 => Pw(3)( 70*8-1 downto  69*8), w71 => Pw(3)( 71*8-1 downto  70*8), w72 => Pw(3)( 72*8-1 downto  71*8), 
w73 => Pw(3)( 73*8-1 downto  72*8), w74 => Pw(3)( 74*8-1 downto  73*8), w75 => Pw(3)( 75*8-1 downto  74*8), w76 => Pw(3)( 76*8-1 downto  75*8), w77 => Pw(3)( 77*8-1 downto  76*8), w78 => Pw(3)( 78*8-1 downto  77*8), w79 => Pw(3)( 79*8-1 downto  78*8), w80 => Pw(3)( 80*8-1 downto  79*8), 
w81 => Pw(3)( 81*8-1 downto  80*8), w82 => Pw(3)( 82*8-1 downto  81*8), w83 => Pw(3)( 83*8-1 downto  82*8), w84 => Pw(3)( 84*8-1 downto  83*8), w85 => Pw(3)( 85*8-1 downto  84*8), w86 => Pw(3)( 86*8-1 downto  85*8), w87 => Pw(3)( 87*8-1 downto  86*8), w88 => Pw(3)( 88*8-1 downto  87*8), 
w89 => Pw(3)( 89*8-1 downto  88*8), w90 => Pw(3)( 90*8-1 downto  89*8), w91 => Pw(3)( 91*8-1 downto  90*8), w92 => Pw(3)( 92*8-1 downto  91*8), w93 => Pw(3)( 93*8-1 downto  92*8), w94 => Pw(3)( 94*8-1 downto  93*8), w95 => Pw(3)( 95*8-1 downto  94*8), w96 => Pw(3)( 96*8-1 downto  95*8), 
w97 => Pw(3)( 97*8-1 downto  96*8), w98 => Pw(3)( 98*8-1 downto  97*8), w99 => Pw(3)( 99*8-1 downto  98*8), w100=> Pw(3)(100*8-1 downto  99*8), w101=> Pw(3)(101*8-1 downto 100*8), w102=> Pw(3)(102*8-1 downto 101*8), w103=> Pw(3)(103*8-1 downto 102*8), w104=> Pw(3)(104*8-1 downto 103*8), 
w105=> Pw(3)(105*8-1 downto 104*8), w106=> Pw(3)(106*8-1 downto 105*8), w107=> Pw(3)(107*8-1 downto 106*8), w108=> Pw(3)(108*8-1 downto 107*8), w109=> Pw(3)(109*8-1 downto 108*8), w110=> Pw(3)(110*8-1 downto 109*8), w111=> Pw(3)(111*8-1 downto 110*8), w112=> Pw(3)(112*8-1 downto 111*8), 
w113=> Pw(3)(113*8-1 downto 112*8), w114=> Pw(3)(114*8-1 downto 113*8), w115=> Pw(3)(115*8-1 downto 114*8), w116=> Pw(3)(116*8-1 downto 115*8), w117=> Pw(3)(117*8-1 downto 116*8), w118=> Pw(3)(118*8-1 downto 117*8), w119=> Pw(3)(119*8-1 downto 118*8), w120=> Pw(3)(120*8-1 downto 119*8), 
w121=> Pw(3)(121*8-1 downto 120*8), w122=> Pw(3)(122*8-1 downto 121*8), w123=> Pw(3)(123*8-1 downto 122*8), w124=> Pw(3)(124*8-1 downto 123*8), w125=> Pw(3)(125*8-1 downto 124*8), w126=> Pw(3)(126*8-1 downto 125*8), w127=> Pw(3)(127*8-1 downto 126*8), w128=> Pw(3)(128*8-1 downto 127*8), 

           d_out   => pca_d03_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_4_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,
  
w01 => Pw( 4)(     7 downto    0), w02 => Pw( 4)( 2*8-1 downto    8), w03 => Pw( 4)( 3*8-1 downto  2*8), w04 => Pw( 4)( 4*8-1 downto  3*8), w05 => Pw( 4)( 5*8-1 downto  4*8), w06 => Pw( 4)( 6*8-1 downto  5*8), w07 => Pw( 4)( 7*8-1 downto  6*8), w08 => Pw( 4)( 8*8-1 downto  7*8),  
w09 => Pw( 4)( 9*8-1 downto  8*8), w10 => Pw( 4)(10*8-1 downto  9*8), w11 => Pw( 4)(11*8-1 downto 10*8), w12 => Pw( 4)(12*8-1 downto 11*8), w13 => Pw( 4)(13*8-1 downto 12*8), w14 => Pw( 4)(14*8-1 downto 13*8), w15 => Pw( 4)(15*8-1 downto 14*8), w16 => Pw( 4)(16*8-1 downto 15*8),  
w17 => Pw( 4)(17*8-1 downto 16*8), w18 => Pw( 4)(18*8-1 downto 17*8), w19 => Pw( 4)(19*8-1 downto 18*8), w20 => Pw( 4)(20*8-1 downto 19*8), w21 => Pw( 4)(21*8-1 downto 20*8), w22 => Pw( 4)(22*8-1 downto 21*8), w23 => Pw( 4)(23*8-1 downto 22*8), w24 => Pw( 4)(24*8-1 downto 23*8),  
w25 => Pw( 4)(25*8-1 downto 24*8), w26 => Pw( 4)(26*8-1 downto 25*8), w27 => Pw( 4)(27*8-1 downto 26*8), w28 => Pw( 4)(28*8-1 downto 27*8), w29 => Pw( 4)(29*8-1 downto 28*8), w30 => Pw( 4)(30*8-1 downto 29*8), w31 => Pw( 4)(31*8-1 downto 30*8), w32 => Pw( 4)(32*8-1 downto 31*8),  
w33 => Pw( 4)(33*8-1 downto 32*8), w34 => Pw( 4)(34*8-1 downto 33*8), w35 => Pw( 4)(35*8-1 downto 34*8), w36 => Pw( 4)(36*8-1 downto 35*8), w37 => Pw( 4)(37*8-1 downto 36*8), w38 => Pw( 4)(38*8-1 downto 37*8), w39 => Pw( 4)(39*8-1 downto 38*8), w40 => Pw( 4)(40*8-1 downto 39*8),  
w41 => Pw( 4)(41*8-1 downto 40*8), w42 => Pw( 4)(42*8-1 downto 41*8), w43 => Pw( 4)(43*8-1 downto 42*8), w44 => Pw( 4)(44*8-1 downto 43*8), w45 => Pw( 4)(45*8-1 downto 44*8), w46 => Pw( 4)(46*8-1 downto 45*8), w47 => Pw( 4)(47*8-1 downto 46*8), w48 => Pw( 4)(48*8-1 downto 47*8),  
w49 => Pw( 4)(49*8-1 downto 48*8), w50 => Pw( 4)(50*8-1 downto 49*8), w51 => Pw( 4)(51*8-1 downto 50*8), w52 => Pw( 4)(52*8-1 downto 51*8), w53 => Pw( 4)(53*8-1 downto 52*8), w54 => Pw( 4)(54*8-1 downto 53*8), w55 => Pw( 4)(55*8-1 downto 54*8), w56 => Pw( 4)(56*8-1 downto 55*8),  
w57 => Pw( 4)(57*8-1 downto 56*8), w58 => Pw( 4)(58*8-1 downto 57*8), w59 => Pw( 4)(59*8-1 downto 58*8), w60 => Pw( 4)(60*8-1 downto 59*8), w61 => Pw( 4)(61*8-1 downto 60*8), w62 => Pw( 4)(62*8-1 downto 61*8), w63 => Pw( 4)(63*8-1 downto 62*8), w64 => Pw( 4)(64*8-1 downto 63*8), 
w65 => Pw(4)( 65*8-1 downto  64*8), w66 => Pw(4)( 66*8-1 downto  65*8), w67 => Pw(4)( 67*8-1 downto  66*8), w68 => Pw(4)( 68*8-1 downto  67*8), w69 => Pw(4)( 69*8-1 downto  68*8), w70 => Pw(4)( 70*8-1 downto  69*8), w71 => Pw(4)( 71*8-1 downto  70*8), w72 => Pw(4)( 72*8-1 downto  71*8), 
w73 => Pw(4)( 73*8-1 downto  72*8), w74 => Pw(4)( 74*8-1 downto  73*8), w75 => Pw(4)( 75*8-1 downto  74*8), w76 => Pw(4)( 76*8-1 downto  75*8), w77 => Pw(4)( 77*8-1 downto  76*8), w78 => Pw(4)( 78*8-1 downto  77*8), w79 => Pw(4)( 79*8-1 downto  78*8), w80 => Pw(4)( 80*8-1 downto  79*8), 
w81 => Pw(4)( 81*8-1 downto  80*8), w82 => Pw(4)( 82*8-1 downto  81*8), w83 => Pw(4)( 83*8-1 downto  82*8), w84 => Pw(4)( 84*8-1 downto  83*8), w85 => Pw(4)( 85*8-1 downto  84*8), w86 => Pw(4)( 86*8-1 downto  85*8), w87 => Pw(4)( 87*8-1 downto  86*8), w88 => Pw(4)( 88*8-1 downto  87*8), 
w89 => Pw(4)( 89*8-1 downto  88*8), w90 => Pw(4)( 90*8-1 downto  89*8), w91 => Pw(4)( 91*8-1 downto  90*8), w92 => Pw(4)( 92*8-1 downto  91*8), w93 => Pw(4)( 93*8-1 downto  92*8), w94 => Pw(4)( 94*8-1 downto  93*8), w95 => Pw(4)( 95*8-1 downto  94*8), w96 => Pw(4)( 96*8-1 downto  95*8), 
w97 => Pw(4)( 97*8-1 downto  96*8), w98 => Pw(4)( 98*8-1 downto  97*8), w99 => Pw(4)( 99*8-1 downto  98*8), w100=> Pw(4)(100*8-1 downto  99*8), w101=> Pw(4)(101*8-1 downto 100*8), w102=> Pw(4)(102*8-1 downto 101*8), w103=> Pw(4)(103*8-1 downto 102*8), w104=> Pw(4)(104*8-1 downto 103*8), 
w105=> Pw(4)(105*8-1 downto 104*8), w106=> Pw(4)(106*8-1 downto 105*8), w107=> Pw(4)(107*8-1 downto 106*8), w108=> Pw(4)(108*8-1 downto 107*8), w109=> Pw(4)(109*8-1 downto 108*8), w110=> Pw(4)(110*8-1 downto 109*8), w111=> Pw(4)(111*8-1 downto 110*8), w112=> Pw(4)(112*8-1 downto 111*8), 
w113=> Pw(4)(113*8-1 downto 112*8), w114=> Pw(4)(114*8-1 downto 113*8), w115=> Pw(4)(115*8-1 downto 114*8), w116=> Pw(4)(116*8-1 downto 115*8), w117=> Pw(4)(117*8-1 downto 116*8), w118=> Pw(4)(118*8-1 downto 117*8), w119=> Pw(4)(119*8-1 downto 118*8), w120=> Pw(4)(120*8-1 downto 119*8), 
w121=> Pw(4)(121*8-1 downto 120*8), w122=> Pw(4)(122*8-1 downto 121*8), w123=> Pw(4)(123*8-1 downto 122*8), w124=> Pw(4)(124*8-1 downto 123*8), w125=> Pw(4)(125*8-1 downto 124*8), w126=> Pw(4)(126*8-1 downto 125*8), w127=> Pw(4)(127*8-1 downto 126*8), w128=> Pw(4)(128*8-1 downto 127*8), 

           d_out   => pca_d04_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_5_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 5)(     7 downto    0), w02 => Pw( 5)( 2*8-1 downto    8), w03 => Pw( 5)( 3*8-1 downto  2*8), w04 => Pw( 5)( 4*8-1 downto  3*8), w05 => Pw( 5)( 5*8-1 downto  4*8), w06 => Pw( 5)( 6*8-1 downto  5*8), w07 => Pw( 5)( 7*8-1 downto  6*8), w08 => Pw( 5)( 8*8-1 downto  7*8),  
w09 => Pw( 5)( 9*8-1 downto  8*8), w10 => Pw( 5)(10*8-1 downto  9*8), w11 => Pw( 5)(11*8-1 downto 10*8), w12 => Pw( 5)(12*8-1 downto 11*8), w13 => Pw( 5)(13*8-1 downto 12*8), w14 => Pw( 5)(14*8-1 downto 13*8), w15 => Pw( 5)(15*8-1 downto 14*8), w16 => Pw( 5)(16*8-1 downto 15*8),  
w17 => Pw( 5)(17*8-1 downto 16*8), w18 => Pw( 5)(18*8-1 downto 17*8), w19 => Pw( 5)(19*8-1 downto 18*8), w20 => Pw( 5)(20*8-1 downto 19*8), w21 => Pw( 5)(21*8-1 downto 20*8), w22 => Pw( 5)(22*8-1 downto 21*8), w23 => Pw( 5)(23*8-1 downto 22*8), w24 => Pw( 5)(24*8-1 downto 23*8),  
w25 => Pw( 5)(25*8-1 downto 24*8), w26 => Pw( 5)(26*8-1 downto 25*8), w27 => Pw( 5)(27*8-1 downto 26*8), w28 => Pw( 5)(28*8-1 downto 27*8), w29 => Pw( 5)(29*8-1 downto 28*8), w30 => Pw( 5)(30*8-1 downto 29*8), w31 => Pw( 5)(31*8-1 downto 30*8), w32 => Pw( 5)(32*8-1 downto 31*8),  
w33 => Pw( 5)(33*8-1 downto 32*8), w34 => Pw( 5)(34*8-1 downto 33*8), w35 => Pw( 5)(35*8-1 downto 34*8), w36 => Pw( 5)(36*8-1 downto 35*8), w37 => Pw( 5)(37*8-1 downto 36*8), w38 => Pw( 5)(38*8-1 downto 37*8), w39 => Pw( 5)(39*8-1 downto 38*8), w40 => Pw( 5)(40*8-1 downto 39*8),  
w41 => Pw( 5)(41*8-1 downto 40*8), w42 => Pw( 5)(42*8-1 downto 41*8), w43 => Pw( 5)(43*8-1 downto 42*8), w44 => Pw( 5)(44*8-1 downto 43*8), w45 => Pw( 5)(45*8-1 downto 44*8), w46 => Pw( 5)(46*8-1 downto 45*8), w47 => Pw( 5)(47*8-1 downto 46*8), w48 => Pw( 5)(48*8-1 downto 47*8),  
w49 => Pw( 5)(49*8-1 downto 48*8), w50 => Pw( 5)(50*8-1 downto 49*8), w51 => Pw( 5)(51*8-1 downto 50*8), w52 => Pw( 5)(52*8-1 downto 51*8), w53 => Pw( 5)(53*8-1 downto 52*8), w54 => Pw( 5)(54*8-1 downto 53*8), w55 => Pw( 5)(55*8-1 downto 54*8), w56 => Pw( 5)(56*8-1 downto 55*8),  
w57 => Pw( 5)(57*8-1 downto 56*8), w58 => Pw( 5)(58*8-1 downto 57*8), w59 => Pw( 5)(59*8-1 downto 58*8), w60 => Pw( 5)(60*8-1 downto 59*8), w61 => Pw( 5)(61*8-1 downto 60*8), w62 => Pw( 5)(62*8-1 downto 61*8), w63 => Pw( 5)(63*8-1 downto 62*8), w64 => Pw( 5)(64*8-1 downto 63*8), 
w65 => Pw(5)( 65*8-1 downto  64*8), w66 => Pw(5)( 66*8-1 downto  65*8), w67 => Pw(5)( 67*8-1 downto  66*8), w68 => Pw(5)( 68*8-1 downto  67*8), w69 => Pw(5)( 69*8-1 downto  68*8), w70 => Pw(5)( 70*8-1 downto  69*8), w71 => Pw(5)( 71*8-1 downto  70*8), w72 => Pw(5)( 72*8-1 downto  71*8), 
w73 => Pw(5)( 73*8-1 downto  72*8), w74 => Pw(5)( 74*8-1 downto  73*8), w75 => Pw(5)( 75*8-1 downto  74*8), w76 => Pw(5)( 76*8-1 downto  75*8), w77 => Pw(5)( 77*8-1 downto  76*8), w78 => Pw(5)( 78*8-1 downto  77*8), w79 => Pw(5)( 79*8-1 downto  78*8), w80 => Pw(5)( 80*8-1 downto  79*8), 
w81 => Pw(5)( 81*8-1 downto  80*8), w82 => Pw(5)( 82*8-1 downto  81*8), w83 => Pw(5)( 83*8-1 downto  82*8), w84 => Pw(5)( 84*8-1 downto  83*8), w85 => Pw(5)( 85*8-1 downto  84*8), w86 => Pw(5)( 86*8-1 downto  85*8), w87 => Pw(5)( 87*8-1 downto  86*8), w88 => Pw(5)( 88*8-1 downto  87*8), 
w89 => Pw(5)( 89*8-1 downto  88*8), w90 => Pw(5)( 90*8-1 downto  89*8), w91 => Pw(5)( 91*8-1 downto  90*8), w92 => Pw(5)( 92*8-1 downto  91*8), w93 => Pw(5)( 93*8-1 downto  92*8), w94 => Pw(5)( 94*8-1 downto  93*8), w95 => Pw(5)( 95*8-1 downto  94*8), w96 => Pw(5)( 96*8-1 downto  95*8), 
w97 => Pw(5)( 97*8-1 downto  96*8), w98 => Pw(5)( 98*8-1 downto  97*8), w99 => Pw(5)( 99*8-1 downto  98*8), w100=> Pw(5)(100*8-1 downto  99*8), w101=> Pw(5)(101*8-1 downto 100*8), w102=> Pw(5)(102*8-1 downto 101*8), w103=> Pw(5)(103*8-1 downto 102*8), w104=> Pw(5)(104*8-1 downto 103*8), 
w105=> Pw(5)(105*8-1 downto 104*8), w106=> Pw(5)(106*8-1 downto 105*8), w107=> Pw(5)(107*8-1 downto 106*8), w108=> Pw(5)(108*8-1 downto 107*8), w109=> Pw(5)(109*8-1 downto 108*8), w110=> Pw(5)(110*8-1 downto 109*8), w111=> Pw(5)(111*8-1 downto 110*8), w112=> Pw(5)(112*8-1 downto 111*8), 
w113=> Pw(5)(113*8-1 downto 112*8), w114=> Pw(5)(114*8-1 downto 113*8), w115=> Pw(5)(115*8-1 downto 114*8), w116=> Pw(5)(116*8-1 downto 115*8), w117=> Pw(5)(117*8-1 downto 116*8), w118=> Pw(5)(118*8-1 downto 117*8), w119=> Pw(5)(119*8-1 downto 118*8), w120=> Pw(5)(120*8-1 downto 119*8), 
w121=> Pw(5)(121*8-1 downto 120*8), w122=> Pw(5)(122*8-1 downto 121*8), w123=> Pw(5)(123*8-1 downto 122*8), w124=> Pw(5)(124*8-1 downto 123*8), w125=> Pw(5)(125*8-1 downto 124*8), w126=> Pw(5)(126*8-1 downto 125*8), w127=> Pw(5)(127*8-1 downto 126*8), w128=> Pw(5)(128*8-1 downto 127*8), 

           d_out   => pca_d05_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_6_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 6)(     7 downto    0), w02 => Pw( 6)( 2*8-1 downto    8), w03 => Pw( 6)( 3*8-1 downto  2*8), w04 => Pw( 6)( 4*8-1 downto  3*8), w05 => Pw( 6)( 5*8-1 downto  4*8), w06 => Pw( 6)( 6*8-1 downto  5*8), w07 => Pw( 6)( 7*8-1 downto  6*8), w08 => Pw( 6)( 8*8-1 downto  7*8),  
w09 => Pw( 6)( 9*8-1 downto  8*8), w10 => Pw( 6)(10*8-1 downto  9*8), w11 => Pw( 6)(11*8-1 downto 10*8), w12 => Pw( 6)(12*8-1 downto 11*8), w13 => Pw( 6)(13*8-1 downto 12*8), w14 => Pw( 6)(14*8-1 downto 13*8), w15 => Pw( 6)(15*8-1 downto 14*8), w16 => Pw( 6)(16*8-1 downto 15*8),  
w17 => Pw( 6)(17*8-1 downto 16*8), w18 => Pw( 6)(18*8-1 downto 17*8), w19 => Pw( 6)(19*8-1 downto 18*8), w20 => Pw( 6)(20*8-1 downto 19*8), w21 => Pw( 6)(21*8-1 downto 20*8), w22 => Pw( 6)(22*8-1 downto 21*8), w23 => Pw( 6)(23*8-1 downto 22*8), w24 => Pw( 6)(24*8-1 downto 23*8),  
w25 => Pw( 6)(25*8-1 downto 24*8), w26 => Pw( 6)(26*8-1 downto 25*8), w27 => Pw( 6)(27*8-1 downto 26*8), w28 => Pw( 6)(28*8-1 downto 27*8), w29 => Pw( 6)(29*8-1 downto 28*8), w30 => Pw( 6)(30*8-1 downto 29*8), w31 => Pw( 6)(31*8-1 downto 30*8), w32 => Pw( 6)(32*8-1 downto 31*8),  
w33 => Pw( 6)(33*8-1 downto 32*8), w34 => Pw( 6)(34*8-1 downto 33*8), w35 => Pw( 6)(35*8-1 downto 34*8), w36 => Pw( 6)(36*8-1 downto 35*8), w37 => Pw( 6)(37*8-1 downto 36*8), w38 => Pw( 6)(38*8-1 downto 37*8), w39 => Pw( 6)(39*8-1 downto 38*8), w40 => Pw( 6)(40*8-1 downto 39*8),  
w41 => Pw( 6)(41*8-1 downto 40*8), w42 => Pw( 6)(42*8-1 downto 41*8), w43 => Pw( 6)(43*8-1 downto 42*8), w44 => Pw( 6)(44*8-1 downto 43*8), w45 => Pw( 6)(45*8-1 downto 44*8), w46 => Pw( 6)(46*8-1 downto 45*8), w47 => Pw( 6)(47*8-1 downto 46*8), w48 => Pw( 6)(48*8-1 downto 47*8),  
w49 => Pw( 6)(49*8-1 downto 48*8), w50 => Pw( 6)(50*8-1 downto 49*8), w51 => Pw( 6)(51*8-1 downto 50*8), w52 => Pw( 6)(52*8-1 downto 51*8), w53 => Pw( 6)(53*8-1 downto 52*8), w54 => Pw( 6)(54*8-1 downto 53*8), w55 => Pw( 6)(55*8-1 downto 54*8), w56 => Pw( 6)(56*8-1 downto 55*8),  
w57 => Pw( 6)(57*8-1 downto 56*8), w58 => Pw( 6)(58*8-1 downto 57*8), w59 => Pw( 6)(59*8-1 downto 58*8), w60 => Pw( 6)(60*8-1 downto 59*8), w61 => Pw( 6)(61*8-1 downto 60*8), w62 => Pw( 6)(62*8-1 downto 61*8), w63 => Pw( 6)(63*8-1 downto 62*8), w64 => Pw( 6)(64*8-1 downto 63*8), 
w65 => Pw(6)( 65*8-1 downto  64*8), w66 => Pw(6)( 66*8-1 downto  65*8), w67 => Pw(6)( 67*8-1 downto  66*8), w68 => Pw(6)( 68*8-1 downto  67*8), w69 => Pw(6)( 69*8-1 downto  68*8), w70 => Pw(6)( 70*8-1 downto  69*8), w71 => Pw(6)( 71*8-1 downto  70*8), w72 => Pw(6)( 72*8-1 downto  71*8), 
w73 => Pw(6)( 73*8-1 downto  72*8), w74 => Pw(6)( 74*8-1 downto  73*8), w75 => Pw(6)( 75*8-1 downto  74*8), w76 => Pw(6)( 76*8-1 downto  75*8), w77 => Pw(6)( 77*8-1 downto  76*8), w78 => Pw(6)( 78*8-1 downto  77*8), w79 => Pw(6)( 79*8-1 downto  78*8), w80 => Pw(6)( 80*8-1 downto  79*8), 
w81 => Pw(6)( 81*8-1 downto  80*8), w82 => Pw(6)( 82*8-1 downto  81*8), w83 => Pw(6)( 83*8-1 downto  82*8), w84 => Pw(6)( 84*8-1 downto  83*8), w85 => Pw(6)( 85*8-1 downto  84*8), w86 => Pw(6)( 86*8-1 downto  85*8), w87 => Pw(6)( 87*8-1 downto  86*8), w88 => Pw(6)( 88*8-1 downto  87*8), 
w89 => Pw(6)( 89*8-1 downto  88*8), w90 => Pw(6)( 90*8-1 downto  89*8), w91 => Pw(6)( 91*8-1 downto  90*8), w92 => Pw(6)( 92*8-1 downto  91*8), w93 => Pw(6)( 93*8-1 downto  92*8), w94 => Pw(6)( 94*8-1 downto  93*8), w95 => Pw(6)( 95*8-1 downto  94*8), w96 => Pw(6)( 96*8-1 downto  95*8), 
w97 => Pw(6)( 97*8-1 downto  96*8), w98 => Pw(6)( 98*8-1 downto  97*8), w99 => Pw(6)( 99*8-1 downto  98*8), w100=> Pw(6)(100*8-1 downto  99*8), w101=> Pw(6)(101*8-1 downto 100*8), w102=> Pw(6)(102*8-1 downto 101*8), w103=> Pw(6)(103*8-1 downto 102*8), w104=> Pw(6)(104*8-1 downto 103*8), 
w105=> Pw(6)(105*8-1 downto 104*8), w106=> Pw(6)(106*8-1 downto 105*8), w107=> Pw(6)(107*8-1 downto 106*8), w108=> Pw(6)(108*8-1 downto 107*8), w109=> Pw(6)(109*8-1 downto 108*8), w110=> Pw(6)(110*8-1 downto 109*8), w111=> Pw(6)(111*8-1 downto 110*8), w112=> Pw(6)(112*8-1 downto 111*8), 
w113=> Pw(6)(113*8-1 downto 112*8), w114=> Pw(6)(114*8-1 downto 113*8), w115=> Pw(6)(115*8-1 downto 114*8), w116=> Pw(6)(116*8-1 downto 115*8), w117=> Pw(6)(117*8-1 downto 116*8), w118=> Pw(6)(118*8-1 downto 117*8), w119=> Pw(6)(119*8-1 downto 118*8), w120=> Pw(6)(120*8-1 downto 119*8), 
w121=> Pw(6)(121*8-1 downto 120*8), w122=> Pw(6)(122*8-1 downto 121*8), w123=> Pw(6)(123*8-1 downto 122*8), w124=> Pw(6)(124*8-1 downto 123*8), w125=> Pw(6)(125*8-1 downto 124*8), w126=> Pw(6)(126*8-1 downto 125*8), w127=> Pw(6)(127*8-1 downto 126*8), w128=> Pw(6)(128*8-1 downto 127*8), 

           d_out   => pca_d06_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_7_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 7)(     7 downto    0), w02 => Pw( 7)( 2*8-1 downto    8), w03 => Pw( 7)( 3*8-1 downto  2*8), w04 => Pw( 7)( 4*8-1 downto  3*8), w05 => Pw( 7)( 5*8-1 downto  4*8), w06 => Pw( 7)( 6*8-1 downto  5*8), w07 => Pw( 7)( 7*8-1 downto  6*8), w08 => Pw( 7)( 8*8-1 downto  7*8),  
w09 => Pw( 7)( 9*8-1 downto  8*8), w10 => Pw( 7)(10*8-1 downto  9*8), w11 => Pw( 7)(11*8-1 downto 10*8), w12 => Pw( 7)(12*8-1 downto 11*8), w13 => Pw( 7)(13*8-1 downto 12*8), w14 => Pw( 7)(14*8-1 downto 13*8), w15 => Pw( 7)(15*8-1 downto 14*8), w16 => Pw( 7)(16*8-1 downto 15*8),  
w17 => Pw( 7)(17*8-1 downto 16*8), w18 => Pw( 7)(18*8-1 downto 17*8), w19 => Pw( 7)(19*8-1 downto 18*8), w20 => Pw( 7)(20*8-1 downto 19*8), w21 => Pw( 7)(21*8-1 downto 20*8), w22 => Pw( 7)(22*8-1 downto 21*8), w23 => Pw( 7)(23*8-1 downto 22*8), w24 => Pw( 7)(24*8-1 downto 23*8),  
w25 => Pw( 7)(25*8-1 downto 24*8), w26 => Pw( 7)(26*8-1 downto 25*8), w27 => Pw( 7)(27*8-1 downto 26*8), w28 => Pw( 7)(28*8-1 downto 27*8), w29 => Pw( 7)(29*8-1 downto 28*8), w30 => Pw( 7)(30*8-1 downto 29*8), w31 => Pw( 7)(31*8-1 downto 30*8), w32 => Pw( 7)(32*8-1 downto 31*8),  
w33 => Pw( 7)(33*8-1 downto 32*8), w34 => Pw( 7)(34*8-1 downto 33*8), w35 => Pw( 7)(35*8-1 downto 34*8), w36 => Pw( 7)(36*8-1 downto 35*8), w37 => Pw( 7)(37*8-1 downto 36*8), w38 => Pw( 7)(38*8-1 downto 37*8), w39 => Pw( 7)(39*8-1 downto 38*8), w40 => Pw( 7)(40*8-1 downto 39*8),  
w41 => Pw( 7)(41*8-1 downto 40*8), w42 => Pw( 7)(42*8-1 downto 41*8), w43 => Pw( 7)(43*8-1 downto 42*8), w44 => Pw( 7)(44*8-1 downto 43*8), w45 => Pw( 7)(45*8-1 downto 44*8), w46 => Pw( 7)(46*8-1 downto 45*8), w47 => Pw( 7)(47*8-1 downto 46*8), w48 => Pw( 7)(48*8-1 downto 47*8),  
w49 => Pw( 7)(49*8-1 downto 48*8), w50 => Pw( 7)(50*8-1 downto 49*8), w51 => Pw( 7)(51*8-1 downto 50*8), w52 => Pw( 7)(52*8-1 downto 51*8), w53 => Pw( 7)(53*8-1 downto 52*8), w54 => Pw( 7)(54*8-1 downto 53*8), w55 => Pw( 7)(55*8-1 downto 54*8), w56 => Pw( 7)(56*8-1 downto 55*8),  
w57 => Pw( 7)(57*8-1 downto 56*8), w58 => Pw( 7)(58*8-1 downto 57*8), w59 => Pw( 7)(59*8-1 downto 58*8), w60 => Pw( 7)(60*8-1 downto 59*8), w61 => Pw( 7)(61*8-1 downto 60*8), w62 => Pw( 7)(62*8-1 downto 61*8), w63 => Pw( 7)(63*8-1 downto 62*8), w64 => Pw( 7)(64*8-1 downto 63*8), 
w65 => Pw(7)( 65*8-1 downto  64*8), w66 => Pw(7)( 66*8-1 downto  65*8), w67 => Pw(7)( 67*8-1 downto  66*8), w68 => Pw(7)( 68*8-1 downto  67*8), w69 => Pw(7)( 69*8-1 downto  68*8), w70 => Pw(7)( 70*8-1 downto  69*8), w71 => Pw(7)( 71*8-1 downto  70*8), w72 => Pw(7)( 72*8-1 downto  71*8), 
w73 => Pw(7)( 73*8-1 downto  72*8), w74 => Pw(7)( 74*8-1 downto  73*8), w75 => Pw(7)( 75*8-1 downto  74*8), w76 => Pw(7)( 76*8-1 downto  75*8), w77 => Pw(7)( 77*8-1 downto  76*8), w78 => Pw(7)( 78*8-1 downto  77*8), w79 => Pw(7)( 79*8-1 downto  78*8), w80 => Pw(7)( 80*8-1 downto  79*8), 
w81 => Pw(7)( 81*8-1 downto  80*8), w82 => Pw(7)( 82*8-1 downto  81*8), w83 => Pw(7)( 83*8-1 downto  82*8), w84 => Pw(7)( 84*8-1 downto  83*8), w85 => Pw(7)( 85*8-1 downto  84*8), w86 => Pw(7)( 86*8-1 downto  85*8), w87 => Pw(7)( 87*8-1 downto  86*8), w88 => Pw(7)( 88*8-1 downto  87*8), 
w89 => Pw(7)( 89*8-1 downto  88*8), w90 => Pw(7)( 90*8-1 downto  89*8), w91 => Pw(7)( 91*8-1 downto  90*8), w92 => Pw(7)( 92*8-1 downto  91*8), w93 => Pw(7)( 93*8-1 downto  92*8), w94 => Pw(7)( 94*8-1 downto  93*8), w95 => Pw(7)( 95*8-1 downto  94*8), w96 => Pw(7)( 96*8-1 downto  95*8), 
w97 => Pw(7)( 97*8-1 downto  96*8), w98 => Pw(7)( 98*8-1 downto  97*8), w99 => Pw(7)( 99*8-1 downto  98*8), w100=> Pw(7)(100*8-1 downto  99*8), w101=> Pw(7)(101*8-1 downto 100*8), w102=> Pw(7)(102*8-1 downto 101*8), w103=> Pw(7)(103*8-1 downto 102*8), w104=> Pw(7)(104*8-1 downto 103*8), 
w105=> Pw(7)(105*8-1 downto 104*8), w106=> Pw(7)(106*8-1 downto 105*8), w107=> Pw(7)(107*8-1 downto 106*8), w108=> Pw(7)(108*8-1 downto 107*8), w109=> Pw(7)(109*8-1 downto 108*8), w110=> Pw(7)(110*8-1 downto 109*8), w111=> Pw(7)(111*8-1 downto 110*8), w112=> Pw(7)(112*8-1 downto 111*8), 
w113=> Pw(7)(113*8-1 downto 112*8), w114=> Pw(7)(114*8-1 downto 113*8), w115=> Pw(7)(115*8-1 downto 114*8), w116=> Pw(7)(116*8-1 downto 115*8), w117=> Pw(7)(117*8-1 downto 116*8), w118=> Pw(7)(118*8-1 downto 117*8), w119=> Pw(7)(119*8-1 downto 118*8), w120=> Pw(7)(120*8-1 downto 119*8), 
w121=> Pw(7)(121*8-1 downto 120*8), w122=> Pw(7)(122*8-1 downto 121*8), w123=> Pw(7)(123*8-1 downto 122*8), w124=> Pw(7)(124*8-1 downto 123*8), w125=> Pw(7)(125*8-1 downto 124*8), w126=> Pw(7)(126*8-1 downto 125*8), w127=> Pw(7)(127*8-1 downto 126*8), w128=> Pw(7)(128*8-1 downto 127*8), 

           d_out   => pca_d07_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_8_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 8)(     7 downto    0), w02 => Pw( 8)( 2*8-1 downto    8), w03 => Pw( 8)( 3*8-1 downto  2*8), w04 => Pw( 8)( 4*8-1 downto  3*8), w05 => Pw( 8)( 5*8-1 downto  4*8), w06 => Pw( 8)( 6*8-1 downto  5*8), w07 => Pw( 8)( 7*8-1 downto  6*8), w08 => Pw( 8)( 8*8-1 downto  7*8),  
w09 => Pw( 8)( 9*8-1 downto  8*8), w10 => Pw( 8)(10*8-1 downto  9*8), w11 => Pw( 8)(11*8-1 downto 10*8), w12 => Pw( 8)(12*8-1 downto 11*8), w13 => Pw( 8)(13*8-1 downto 12*8), w14 => Pw( 8)(14*8-1 downto 13*8), w15 => Pw( 8)(15*8-1 downto 14*8), w16 => Pw( 8)(16*8-1 downto 15*8),  
w17 => Pw( 8)(17*8-1 downto 16*8), w18 => Pw( 8)(18*8-1 downto 17*8), w19 => Pw( 8)(19*8-1 downto 18*8), w20 => Pw( 8)(20*8-1 downto 19*8), w21 => Pw( 8)(21*8-1 downto 20*8), w22 => Pw( 8)(22*8-1 downto 21*8), w23 => Pw( 8)(23*8-1 downto 22*8), w24 => Pw( 8)(24*8-1 downto 23*8),  
w25 => Pw( 8)(25*8-1 downto 24*8), w26 => Pw( 8)(26*8-1 downto 25*8), w27 => Pw( 8)(27*8-1 downto 26*8), w28 => Pw( 8)(28*8-1 downto 27*8), w29 => Pw( 8)(29*8-1 downto 28*8), w30 => Pw( 8)(30*8-1 downto 29*8), w31 => Pw( 8)(31*8-1 downto 30*8), w32 => Pw( 8)(32*8-1 downto 31*8),  
w33 => Pw( 8)(33*8-1 downto 32*8), w34 => Pw( 8)(34*8-1 downto 33*8), w35 => Pw( 8)(35*8-1 downto 34*8), w36 => Pw( 8)(36*8-1 downto 35*8), w37 => Pw( 8)(37*8-1 downto 36*8), w38 => Pw( 8)(38*8-1 downto 37*8), w39 => Pw( 8)(39*8-1 downto 38*8), w40 => Pw( 8)(40*8-1 downto 39*8),  
w41 => Pw( 8)(41*8-1 downto 40*8), w42 => Pw( 8)(42*8-1 downto 41*8), w43 => Pw( 8)(43*8-1 downto 42*8), w44 => Pw( 8)(44*8-1 downto 43*8), w45 => Pw( 8)(45*8-1 downto 44*8), w46 => Pw( 8)(46*8-1 downto 45*8), w47 => Pw( 8)(47*8-1 downto 46*8), w48 => Pw( 8)(48*8-1 downto 47*8),  
w49 => Pw( 8)(49*8-1 downto 48*8), w50 => Pw( 8)(50*8-1 downto 49*8), w51 => Pw( 8)(51*8-1 downto 50*8), w52 => Pw( 8)(52*8-1 downto 51*8), w53 => Pw( 8)(53*8-1 downto 52*8), w54 => Pw( 8)(54*8-1 downto 53*8), w55 => Pw( 8)(55*8-1 downto 54*8), w56 => Pw( 8)(56*8-1 downto 55*8),  
w57 => Pw( 8)(57*8-1 downto 56*8), w58 => Pw( 8)(58*8-1 downto 57*8), w59 => Pw( 8)(59*8-1 downto 58*8), w60 => Pw( 8)(60*8-1 downto 59*8), w61 => Pw( 8)(61*8-1 downto 60*8), w62 => Pw( 8)(62*8-1 downto 61*8), w63 => Pw( 8)(63*8-1 downto 62*8), w64 => Pw( 8)(64*8-1 downto 63*8), 
w65 => Pw(8)( 65*8-1 downto  64*8), w66 => Pw(8)( 66*8-1 downto  65*8), w67 => Pw(8)( 67*8-1 downto  66*8), w68 => Pw(8)( 68*8-1 downto  67*8), w69 => Pw(8)( 69*8-1 downto  68*8), w70 => Pw(8)( 70*8-1 downto  69*8), w71 => Pw(8)( 71*8-1 downto  70*8), w72 => Pw(8)( 72*8-1 downto  71*8), 
w73 => Pw(8)( 73*8-1 downto  72*8), w74 => Pw(8)( 74*8-1 downto  73*8), w75 => Pw(8)( 75*8-1 downto  74*8), w76 => Pw(8)( 76*8-1 downto  75*8), w77 => Pw(8)( 77*8-1 downto  76*8), w78 => Pw(8)( 78*8-1 downto  77*8), w79 => Pw(8)( 79*8-1 downto  78*8), w80 => Pw(8)( 80*8-1 downto  79*8), 
w81 => Pw(8)( 81*8-1 downto  80*8), w82 => Pw(8)( 82*8-1 downto  81*8), w83 => Pw(8)( 83*8-1 downto  82*8), w84 => Pw(8)( 84*8-1 downto  83*8), w85 => Pw(8)( 85*8-1 downto  84*8), w86 => Pw(8)( 86*8-1 downto  85*8), w87 => Pw(8)( 87*8-1 downto  86*8), w88 => Pw(8)( 88*8-1 downto  87*8), 
w89 => Pw(8)( 89*8-1 downto  88*8), w90 => Pw(8)( 90*8-1 downto  89*8), w91 => Pw(8)( 91*8-1 downto  90*8), w92 => Pw(8)( 92*8-1 downto  91*8), w93 => Pw(8)( 93*8-1 downto  92*8), w94 => Pw(8)( 94*8-1 downto  93*8), w95 => Pw(8)( 95*8-1 downto  94*8), w96 => Pw(8)( 96*8-1 downto  95*8), 
w97 => Pw(8)( 97*8-1 downto  96*8), w98 => Pw(8)( 98*8-1 downto  97*8), w99 => Pw(8)( 99*8-1 downto  98*8), w100=> Pw(8)(100*8-1 downto  99*8), w101=> Pw(8)(101*8-1 downto 100*8), w102=> Pw(8)(102*8-1 downto 101*8), w103=> Pw(8)(103*8-1 downto 102*8), w104=> Pw(8)(104*8-1 downto 103*8), 
w105=> Pw(8)(105*8-1 downto 104*8), w106=> Pw(8)(106*8-1 downto 105*8), w107=> Pw(8)(107*8-1 downto 106*8), w108=> Pw(8)(108*8-1 downto 107*8), w109=> Pw(8)(109*8-1 downto 108*8), w110=> Pw(8)(110*8-1 downto 109*8), w111=> Pw(8)(111*8-1 downto 110*8), w112=> Pw(8)(112*8-1 downto 111*8), 
w113=> Pw(8)(113*8-1 downto 112*8), w114=> Pw(8)(114*8-1 downto 113*8), w115=> Pw(8)(115*8-1 downto 114*8), w116=> Pw(8)(116*8-1 downto 115*8), w117=> Pw(8)(117*8-1 downto 116*8), w118=> Pw(8)(118*8-1 downto 117*8), w119=> Pw(8)(119*8-1 downto 118*8), w120=> Pw(8)(120*8-1 downto 119*8), 
w121=> Pw(8)(121*8-1 downto 120*8), w122=> Pw(8)(122*8-1 downto 121*8), w123=> Pw(8)(123*8-1 downto 122*8), w124=> Pw(8)(124*8-1 downto 123*8), w125=> Pw(8)(125*8-1 downto 124*8), w126=> Pw(8)(126*8-1 downto 125*8), w127=> Pw(8)(127*8-1 downto 126*8), w128=> Pw(8)(128*8-1 downto 127*8), 

           d_out   => pca_d08_out   ,
           en_out  => open  ,
           sof_out => open );

  
  PCA128_9_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw( 9)(     7 downto    0), w02 => Pw( 9)( 2*8-1 downto    8), w03 => Pw( 9)( 3*8-1 downto  2*8), w04 => Pw( 9)( 4*8-1 downto  3*8), w05 => Pw( 9)( 5*8-1 downto  4*8), w06 => Pw( 9)( 6*8-1 downto  5*8), w07 => Pw( 9)( 7*8-1 downto  6*8), w08 => Pw( 9)( 8*8-1 downto  7*8),  
w09 => Pw( 9)( 9*8-1 downto  8*8), w10 => Pw( 9)(10*8-1 downto  9*8), w11 => Pw( 9)(11*8-1 downto 10*8), w12 => Pw( 9)(12*8-1 downto 11*8), w13 => Pw( 9)(13*8-1 downto 12*8), w14 => Pw( 9)(14*8-1 downto 13*8), w15 => Pw( 9)(15*8-1 downto 14*8), w16 => Pw( 9)(16*8-1 downto 15*8),  
w17 => Pw( 9)(17*8-1 downto 16*8), w18 => Pw( 9)(18*8-1 downto 17*8), w19 => Pw( 9)(19*8-1 downto 18*8), w20 => Pw( 9)(20*8-1 downto 19*8), w21 => Pw( 9)(21*8-1 downto 20*8), w22 => Pw( 9)(22*8-1 downto 21*8), w23 => Pw( 9)(23*8-1 downto 22*8), w24 => Pw( 9)(24*8-1 downto 23*8),  
w25 => Pw( 9)(25*8-1 downto 24*8), w26 => Pw( 9)(26*8-1 downto 25*8), w27 => Pw( 9)(27*8-1 downto 26*8), w28 => Pw( 9)(28*8-1 downto 27*8), w29 => Pw( 9)(29*8-1 downto 28*8), w30 => Pw( 9)(30*8-1 downto 29*8), w31 => Pw( 9)(31*8-1 downto 30*8), w32 => Pw( 9)(32*8-1 downto 31*8),  
w33 => Pw( 9)(33*8-1 downto 32*8), w34 => Pw( 9)(34*8-1 downto 33*8), w35 => Pw( 9)(35*8-1 downto 34*8), w36 => Pw( 9)(36*8-1 downto 35*8), w37 => Pw( 9)(37*8-1 downto 36*8), w38 => Pw( 9)(38*8-1 downto 37*8), w39 => Pw( 9)(39*8-1 downto 38*8), w40 => Pw( 9)(40*8-1 downto 39*8),  
w41 => Pw( 9)(41*8-1 downto 40*8), w42 => Pw( 9)(42*8-1 downto 41*8), w43 => Pw( 9)(43*8-1 downto 42*8), w44 => Pw( 9)(44*8-1 downto 43*8), w45 => Pw( 9)(45*8-1 downto 44*8), w46 => Pw( 9)(46*8-1 downto 45*8), w47 => Pw( 9)(47*8-1 downto 46*8), w48 => Pw( 9)(48*8-1 downto 47*8),  
w49 => Pw( 9)(49*8-1 downto 48*8), w50 => Pw( 9)(50*8-1 downto 49*8), w51 => Pw( 9)(51*8-1 downto 50*8), w52 => Pw( 9)(52*8-1 downto 51*8), w53 => Pw( 9)(53*8-1 downto 52*8), w54 => Pw( 9)(54*8-1 downto 53*8), w55 => Pw( 9)(55*8-1 downto 54*8), w56 => Pw( 9)(56*8-1 downto 55*8),  
w57 => Pw( 9)(57*8-1 downto 56*8), w58 => Pw( 9)(58*8-1 downto 57*8), w59 => Pw( 9)(59*8-1 downto 58*8), w60 => Pw( 9)(60*8-1 downto 59*8), w61 => Pw( 9)(61*8-1 downto 60*8), w62 => Pw( 9)(62*8-1 downto 61*8), w63 => Pw( 9)(63*8-1 downto 62*8), w64 => Pw( 9)(64*8-1 downto 63*8), 
w65 => Pw(9)( 65*8-1 downto  64*8), w66 => Pw(9)( 66*8-1 downto  65*8), w67 => Pw(9)( 67*8-1 downto  66*8), w68 => Pw(9)( 68*8-1 downto  67*8), w69 => Pw(9)( 69*8-1 downto  68*8), w70 => Pw(9)( 70*8-1 downto  69*8), w71 => Pw(9)( 71*8-1 downto  70*8), w72 => Pw(9)( 72*8-1 downto  71*8), 
w73 => Pw(9)( 73*8-1 downto  72*8), w74 => Pw(9)( 74*8-1 downto  73*8), w75 => Pw(9)( 75*8-1 downto  74*8), w76 => Pw(9)( 76*8-1 downto  75*8), w77 => Pw(9)( 77*8-1 downto  76*8), w78 => Pw(9)( 78*8-1 downto  77*8), w79 => Pw(9)( 79*8-1 downto  78*8), w80 => Pw(9)( 80*8-1 downto  79*8), 
w81 => Pw(9)( 81*8-1 downto  80*8), w82 => Pw(9)( 82*8-1 downto  81*8), w83 => Pw(9)( 83*8-1 downto  82*8), w84 => Pw(9)( 84*8-1 downto  83*8), w85 => Pw(9)( 85*8-1 downto  84*8), w86 => Pw(9)( 86*8-1 downto  85*8), w87 => Pw(9)( 87*8-1 downto  86*8), w88 => Pw(9)( 88*8-1 downto  87*8), 
w89 => Pw(9)( 89*8-1 downto  88*8), w90 => Pw(9)( 90*8-1 downto  89*8), w91 => Pw(9)( 91*8-1 downto  90*8), w92 => Pw(9)( 92*8-1 downto  91*8), w93 => Pw(9)( 93*8-1 downto  92*8), w94 => Pw(9)( 94*8-1 downto  93*8), w95 => Pw(9)( 95*8-1 downto  94*8), w96 => Pw(9)( 96*8-1 downto  95*8), 
w97 => Pw(9)( 97*8-1 downto  96*8), w98 => Pw(9)( 98*8-1 downto  97*8), w99 => Pw(9)( 99*8-1 downto  98*8), w100=> Pw(9)(100*8-1 downto  99*8), w101=> Pw(9)(101*8-1 downto 100*8), w102=> Pw(9)(102*8-1 downto 101*8), w103=> Pw(9)(103*8-1 downto 102*8), w104=> Pw(9)(104*8-1 downto 103*8), 
w105=> Pw(9)(105*8-1 downto 104*8), w106=> Pw(9)(106*8-1 downto 105*8), w107=> Pw(9)(107*8-1 downto 106*8), w108=> Pw(9)(108*8-1 downto 107*8), w109=> Pw(9)(109*8-1 downto 108*8), w110=> Pw(9)(110*8-1 downto 109*8), w111=> Pw(9)(111*8-1 downto 110*8), w112=> Pw(9)(112*8-1 downto 111*8), 
w113=> Pw(9)(113*8-1 downto 112*8), w114=> Pw(9)(114*8-1 downto 113*8), w115=> Pw(9)(115*8-1 downto 114*8), w116=> Pw(9)(116*8-1 downto 115*8), w117=> Pw(9)(117*8-1 downto 116*8), w118=> Pw(9)(118*8-1 downto 117*8), w119=> Pw(9)(119*8-1 downto 118*8), w120=> Pw(9)(120*8-1 downto 119*8), 
w121=> Pw(9)(121*8-1 downto 120*8), w122=> Pw(9)(122*8-1 downto 121*8), w123=> Pw(9)(123*8-1 downto 122*8), w124=> Pw(9)(124*8-1 downto 123*8), w125=> Pw(9)(125*8-1 downto 124*8), w126=> Pw(9)(126*8-1 downto 125*8), w127=> Pw(9)(127*8-1 downto 126*8), w128=> Pw(9)(128*8-1 downto 127*8), 

           d_out   => pca_d09_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_10_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(10)(     7 downto    0), w02 => Pw(10)( 2*8-1 downto    8), w03 => Pw(10)( 3*8-1 downto  2*8), w04 => Pw(10)( 4*8-1 downto  3*8), w05 => Pw(10)( 5*8-1 downto  4*8), w06 => Pw(10)( 6*8-1 downto  5*8), w07 => Pw(10)( 7*8-1 downto  6*8), w08 => Pw(10)( 8*8-1 downto  7*8),  
w09 => Pw(10)( 9*8-1 downto  8*8), w10 => Pw(10)(10*8-1 downto  9*8), w11 => Pw(10)(11*8-1 downto 10*8), w12 => Pw(10)(12*8-1 downto 11*8), w13 => Pw(10)(13*8-1 downto 12*8), w14 => Pw(10)(14*8-1 downto 13*8), w15 => Pw(10)(15*8-1 downto 14*8), w16 => Pw(10)(16*8-1 downto 15*8),  
w17 => Pw(10)(17*8-1 downto 16*8), w18 => Pw(10)(18*8-1 downto 17*8), w19 => Pw(10)(19*8-1 downto 18*8), w20 => Pw(10)(20*8-1 downto 19*8), w21 => Pw(10)(21*8-1 downto 20*8), w22 => Pw(10)(22*8-1 downto 21*8), w23 => Pw(10)(23*8-1 downto 22*8), w24 => Pw(10)(24*8-1 downto 23*8),  
w25 => Pw(10)(25*8-1 downto 24*8), w26 => Pw(10)(26*8-1 downto 25*8), w27 => Pw(10)(27*8-1 downto 26*8), w28 => Pw(10)(28*8-1 downto 27*8), w29 => Pw(10)(29*8-1 downto 28*8), w30 => Pw(10)(30*8-1 downto 29*8), w31 => Pw(10)(31*8-1 downto 30*8), w32 => Pw(10)(32*8-1 downto 31*8),  
w33 => Pw(10)(33*8-1 downto 32*8), w34 => Pw(10)(34*8-1 downto 33*8), w35 => Pw(10)(35*8-1 downto 34*8), w36 => Pw(10)(36*8-1 downto 35*8), w37 => Pw(10)(37*8-1 downto 36*8), w38 => Pw(10)(38*8-1 downto 37*8), w39 => Pw(10)(39*8-1 downto 38*8), w40 => Pw(10)(40*8-1 downto 39*8),  
w41 => Pw(10)(41*8-1 downto 40*8), w42 => Pw(10)(42*8-1 downto 41*8), w43 => Pw(10)(43*8-1 downto 42*8), w44 => Pw(10)(44*8-1 downto 43*8), w45 => Pw(10)(45*8-1 downto 44*8), w46 => Pw(10)(46*8-1 downto 45*8), w47 => Pw(10)(47*8-1 downto 46*8), w48 => Pw(10)(48*8-1 downto 47*8),  
w49 => Pw(10)(49*8-1 downto 48*8), w50 => Pw(10)(50*8-1 downto 49*8), w51 => Pw(10)(51*8-1 downto 50*8), w52 => Pw(10)(52*8-1 downto 51*8), w53 => Pw(10)(53*8-1 downto 52*8), w54 => Pw(10)(54*8-1 downto 53*8), w55 => Pw(10)(55*8-1 downto 54*8), w56 => Pw(10)(56*8-1 downto 55*8),  
w57 => Pw(10)(57*8-1 downto 56*8), w58 => Pw(10)(58*8-1 downto 57*8), w59 => Pw(10)(59*8-1 downto 58*8), w60 => Pw(10)(60*8-1 downto 59*8), w61 => Pw(10)(61*8-1 downto 60*8), w62 => Pw(10)(62*8-1 downto 61*8), w63 => Pw(10)(63*8-1 downto 62*8), w64 => Pw(10)(64*8-1 downto 63*8), 
w65 => Pw(10)( 65*8-1 downto  64*8), w66 => Pw(10)( 66*8-1 downto  65*8), w67 => Pw(10)( 67*8-1 downto  66*8), w68 => Pw(10)( 68*8-1 downto  67*8), w69 => Pw(10)( 69*8-1 downto  68*8), w70 => Pw(10)( 70*8-1 downto  69*8), w71 => Pw(10)( 71*8-1 downto  70*8), w72 => Pw(10)( 72*8-1 downto  71*8), 
w73 => Pw(10)( 73*8-1 downto  72*8), w74 => Pw(10)( 74*8-1 downto  73*8), w75 => Pw(10)( 75*8-1 downto  74*8), w76 => Pw(10)( 76*8-1 downto  75*8), w77 => Pw(10)( 77*8-1 downto  76*8), w78 => Pw(10)( 78*8-1 downto  77*8), w79 => Pw(10)( 79*8-1 downto  78*8), w80 => Pw(10)( 80*8-1 downto  79*8), 
w81 => Pw(10)( 81*8-1 downto  80*8), w82 => Pw(10)( 82*8-1 downto  81*8), w83 => Pw(10)( 83*8-1 downto  82*8), w84 => Pw(10)( 84*8-1 downto  83*8), w85 => Pw(10)( 85*8-1 downto  84*8), w86 => Pw(10)( 86*8-1 downto  85*8), w87 => Pw(10)( 87*8-1 downto  86*8), w88 => Pw(10)( 88*8-1 downto  87*8), 
w89 => Pw(10)( 89*8-1 downto  88*8), w90 => Pw(10)( 90*8-1 downto  89*8), w91 => Pw(10)( 91*8-1 downto  90*8), w92 => Pw(10)( 92*8-1 downto  91*8), w93 => Pw(10)( 93*8-1 downto  92*8), w94 => Pw(10)( 94*8-1 downto  93*8), w95 => Pw(10)( 95*8-1 downto  94*8), w96 => Pw(10)( 96*8-1 downto  95*8), 
w97 => Pw(10)( 97*8-1 downto  96*8), w98 => Pw(10)( 98*8-1 downto  97*8), w99 => Pw(10)( 99*8-1 downto  98*8), w100=> Pw(10)(100*8-1 downto  99*8), w101=> Pw(10)(101*8-1 downto 100*8), w102=> Pw(10)(102*8-1 downto 101*8), w103=> Pw(10)(103*8-1 downto 102*8), w104=> Pw(10)(104*8-1 downto 103*8), 
w105=> Pw(10)(105*8-1 downto 104*8), w106=> Pw(10)(106*8-1 downto 105*8), w107=> Pw(10)(107*8-1 downto 106*8), w108=> Pw(10)(108*8-1 downto 107*8), w109=> Pw(10)(109*8-1 downto 108*8), w110=> Pw(10)(110*8-1 downto 109*8), w111=> Pw(10)(111*8-1 downto 110*8), w112=> Pw(10)(112*8-1 downto 111*8), 
w113=> Pw(10)(113*8-1 downto 112*8), w114=> Pw(10)(114*8-1 downto 113*8), w115=> Pw(10)(115*8-1 downto 114*8), w116=> Pw(10)(116*8-1 downto 115*8), w117=> Pw(10)(117*8-1 downto 116*8), w118=> Pw(10)(118*8-1 downto 117*8), w119=> Pw(10)(119*8-1 downto 118*8), w120=> Pw(10)(120*8-1 downto 119*8), 
w121=> Pw(10)(121*8-1 downto 120*8), w122=> Pw(10)(122*8-1 downto 121*8), w123=> Pw(10)(123*8-1 downto 122*8), w124=> Pw(10)(124*8-1 downto 123*8), w125=> Pw(10)(125*8-1 downto 124*8), w126=> Pw(10)(126*8-1 downto 125*8), w127=> Pw(10)(127*8-1 downto 126*8), w128=> Pw(10)(128*8-1 downto 127*8), 

           d_out   => pca_d10_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_11_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(11)(     7 downto    0), w02 => Pw(11)( 2*8-1 downto    8), w03 => Pw(11)( 3*8-1 downto  2*8), w04 => Pw(11)( 4*8-1 downto  3*8), w05 => Pw(11)( 5*8-1 downto  4*8), w06 => Pw(11)( 6*8-1 downto  5*8), w07 => Pw(11)( 7*8-1 downto  6*8), w08 => Pw(11)( 8*8-1 downto  7*8),  
w09 => Pw(11)( 9*8-1 downto  8*8), w10 => Pw(11)(10*8-1 downto  9*8), w11 => Pw(11)(11*8-1 downto 10*8), w12 => Pw(11)(12*8-1 downto 11*8), w13 => Pw(11)(13*8-1 downto 12*8), w14 => Pw(11)(14*8-1 downto 13*8), w15 => Pw(11)(15*8-1 downto 14*8), w16 => Pw(11)(16*8-1 downto 15*8),  
w17 => Pw(11)(17*8-1 downto 16*8), w18 => Pw(11)(18*8-1 downto 17*8), w19 => Pw(11)(19*8-1 downto 18*8), w20 => Pw(11)(20*8-1 downto 19*8), w21 => Pw(11)(21*8-1 downto 20*8), w22 => Pw(11)(22*8-1 downto 21*8), w23 => Pw(11)(23*8-1 downto 22*8), w24 => Pw(11)(24*8-1 downto 23*8),  
w25 => Pw(11)(25*8-1 downto 24*8), w26 => Pw(11)(26*8-1 downto 25*8), w27 => Pw(11)(27*8-1 downto 26*8), w28 => Pw(11)(28*8-1 downto 27*8), w29 => Pw(11)(29*8-1 downto 28*8), w30 => Pw(11)(30*8-1 downto 29*8), w31 => Pw(11)(31*8-1 downto 30*8), w32 => Pw(11)(32*8-1 downto 31*8),  
w33 => Pw(11)(33*8-1 downto 32*8), w34 => Pw(11)(34*8-1 downto 33*8), w35 => Pw(11)(35*8-1 downto 34*8), w36 => Pw(11)(36*8-1 downto 35*8), w37 => Pw(11)(37*8-1 downto 36*8), w38 => Pw(11)(38*8-1 downto 37*8), w39 => Pw(11)(39*8-1 downto 38*8), w40 => Pw(11)(40*8-1 downto 39*8),  
w41 => Pw(11)(41*8-1 downto 40*8), w42 => Pw(11)(42*8-1 downto 41*8), w43 => Pw(11)(43*8-1 downto 42*8), w44 => Pw(11)(44*8-1 downto 43*8), w45 => Pw(11)(45*8-1 downto 44*8), w46 => Pw(11)(46*8-1 downto 45*8), w47 => Pw(11)(47*8-1 downto 46*8), w48 => Pw(11)(48*8-1 downto 47*8),  
w49 => Pw(11)(49*8-1 downto 48*8), w50 => Pw(11)(50*8-1 downto 49*8), w51 => Pw(11)(51*8-1 downto 50*8), w52 => Pw(11)(52*8-1 downto 51*8), w53 => Pw(11)(53*8-1 downto 52*8), w54 => Pw(11)(54*8-1 downto 53*8), w55 => Pw(11)(55*8-1 downto 54*8), w56 => Pw(11)(56*8-1 downto 55*8),  
w57 => Pw(11)(57*8-1 downto 56*8), w58 => Pw(11)(58*8-1 downto 57*8), w59 => Pw(11)(59*8-1 downto 58*8), w60 => Pw(11)(60*8-1 downto 59*8), w61 => Pw(11)(61*8-1 downto 60*8), w62 => Pw(11)(62*8-1 downto 61*8), w63 => Pw(11)(63*8-1 downto 62*8), w64 => Pw(11)(64*8-1 downto 63*8), 
w65 => Pw(11)( 65*8-1 downto  64*8), w66 => Pw(11)( 66*8-1 downto  65*8), w67 => Pw(11)( 67*8-1 downto  66*8), w68 => Pw(11)( 68*8-1 downto  67*8), w69 => Pw(11)( 69*8-1 downto  68*8), w70 => Pw(11)( 70*8-1 downto  69*8), w71 => Pw(11)( 71*8-1 downto  70*8), w72 => Pw(11)( 72*8-1 downto  71*8), 
w73 => Pw(11)( 73*8-1 downto  72*8), w74 => Pw(11)( 74*8-1 downto  73*8), w75 => Pw(11)( 75*8-1 downto  74*8), w76 => Pw(11)( 76*8-1 downto  75*8), w77 => Pw(11)( 77*8-1 downto  76*8), w78 => Pw(11)( 78*8-1 downto  77*8), w79 => Pw(11)( 79*8-1 downto  78*8), w80 => Pw(11)( 80*8-1 downto  79*8), 
w81 => Pw(11)( 81*8-1 downto  80*8), w82 => Pw(11)( 82*8-1 downto  81*8), w83 => Pw(11)( 83*8-1 downto  82*8), w84 => Pw(11)( 84*8-1 downto  83*8), w85 => Pw(11)( 85*8-1 downto  84*8), w86 => Pw(11)( 86*8-1 downto  85*8), w87 => Pw(11)( 87*8-1 downto  86*8), w88 => Pw(11)( 88*8-1 downto  87*8), 
w89 => Pw(11)( 89*8-1 downto  88*8), w90 => Pw(11)( 90*8-1 downto  89*8), w91 => Pw(11)( 91*8-1 downto  90*8), w92 => Pw(11)( 92*8-1 downto  91*8), w93 => Pw(11)( 93*8-1 downto  92*8), w94 => Pw(11)( 94*8-1 downto  93*8), w95 => Pw(11)( 95*8-1 downto  94*8), w96 => Pw(11)( 96*8-1 downto  95*8), 
w97 => Pw(11)( 97*8-1 downto  96*8), w98 => Pw(11)( 98*8-1 downto  97*8), w99 => Pw(11)( 99*8-1 downto  98*8), w100=> Pw(11)(100*8-1 downto  99*8), w101=> Pw(11)(101*8-1 downto 100*8), w102=> Pw(11)(102*8-1 downto 101*8), w103=> Pw(11)(103*8-1 downto 102*8), w104=> Pw(11)(104*8-1 downto 103*8), 
w105=> Pw(11)(105*8-1 downto 104*8), w106=> Pw(11)(106*8-1 downto 105*8), w107=> Pw(11)(107*8-1 downto 106*8), w108=> Pw(11)(108*8-1 downto 107*8), w109=> Pw(11)(109*8-1 downto 108*8), w110=> Pw(11)(110*8-1 downto 109*8), w111=> Pw(11)(111*8-1 downto 110*8), w112=> Pw(11)(112*8-1 downto 111*8), 
w113=> Pw(11)(113*8-1 downto 112*8), w114=> Pw(11)(114*8-1 downto 113*8), w115=> Pw(11)(115*8-1 downto 114*8), w116=> Pw(11)(116*8-1 downto 115*8), w117=> Pw(11)(117*8-1 downto 116*8), w118=> Pw(11)(118*8-1 downto 117*8), w119=> Pw(11)(119*8-1 downto 118*8), w120=> Pw(11)(120*8-1 downto 119*8), 
w121=> Pw(11)(121*8-1 downto 120*8), w122=> Pw(11)(122*8-1 downto 121*8), w123=> Pw(11)(123*8-1 downto 122*8), w124=> Pw(11)(124*8-1 downto 123*8), w125=> Pw(11)(125*8-1 downto 124*8), w126=> Pw(11)(126*8-1 downto 125*8), w127=> Pw(11)(127*8-1 downto 126*8), w128=> Pw(11)(128*8-1 downto 127*8), 

           d_out   => pca_d11_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_12_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(12)(     7 downto    0), w02 => Pw(12)( 2*8-1 downto    8), w03 => Pw(12)( 3*8-1 downto  2*8), w04 => Pw(12)( 4*8-1 downto  3*8), w05 => Pw(12)( 5*8-1 downto  4*8), w06 => Pw(12)( 6*8-1 downto  5*8), w07 => Pw(12)( 7*8-1 downto  6*8), w08 => Pw(12)( 8*8-1 downto  7*8),  
w09 => Pw(12)( 9*8-1 downto  8*8), w10 => Pw(12)(10*8-1 downto  9*8), w11 => Pw(12)(11*8-1 downto 10*8), w12 => Pw(12)(12*8-1 downto 11*8), w13 => Pw(12)(13*8-1 downto 12*8), w14 => Pw(12)(14*8-1 downto 13*8), w15 => Pw(12)(15*8-1 downto 14*8), w16 => Pw(12)(16*8-1 downto 15*8),  
w17 => Pw(12)(17*8-1 downto 16*8), w18 => Pw(12)(18*8-1 downto 17*8), w19 => Pw(12)(19*8-1 downto 18*8), w20 => Pw(12)(20*8-1 downto 19*8), w21 => Pw(12)(21*8-1 downto 20*8), w22 => Pw(12)(22*8-1 downto 21*8), w23 => Pw(12)(23*8-1 downto 22*8), w24 => Pw(12)(24*8-1 downto 23*8),  
w25 => Pw(12)(25*8-1 downto 24*8), w26 => Pw(12)(26*8-1 downto 25*8), w27 => Pw(12)(27*8-1 downto 26*8), w28 => Pw(12)(28*8-1 downto 27*8), w29 => Pw(12)(29*8-1 downto 28*8), w30 => Pw(12)(30*8-1 downto 29*8), w31 => Pw(12)(31*8-1 downto 30*8), w32 => Pw(12)(32*8-1 downto 31*8),  
w33 => Pw(12)(33*8-1 downto 32*8), w34 => Pw(12)(34*8-1 downto 33*8), w35 => Pw(12)(35*8-1 downto 34*8), w36 => Pw(12)(36*8-1 downto 35*8), w37 => Pw(12)(37*8-1 downto 36*8), w38 => Pw(12)(38*8-1 downto 37*8), w39 => Pw(12)(39*8-1 downto 38*8), w40 => Pw(12)(40*8-1 downto 39*8),  
w41 => Pw(12)(41*8-1 downto 40*8), w42 => Pw(12)(42*8-1 downto 41*8), w43 => Pw(12)(43*8-1 downto 42*8), w44 => Pw(12)(44*8-1 downto 43*8), w45 => Pw(12)(45*8-1 downto 44*8), w46 => Pw(12)(46*8-1 downto 45*8), w47 => Pw(12)(47*8-1 downto 46*8), w48 => Pw(12)(48*8-1 downto 47*8),  
w49 => Pw(12)(49*8-1 downto 48*8), w50 => Pw(12)(50*8-1 downto 49*8), w51 => Pw(12)(51*8-1 downto 50*8), w52 => Pw(12)(52*8-1 downto 51*8), w53 => Pw(12)(53*8-1 downto 52*8), w54 => Pw(12)(54*8-1 downto 53*8), w55 => Pw(12)(55*8-1 downto 54*8), w56 => Pw(12)(56*8-1 downto 55*8),  
w57 => Pw(12)(57*8-1 downto 56*8), w58 => Pw(12)(58*8-1 downto 57*8), w59 => Pw(12)(59*8-1 downto 58*8), w60 => Pw(12)(60*8-1 downto 59*8), w61 => Pw(12)(61*8-1 downto 60*8), w62 => Pw(12)(62*8-1 downto 61*8), w63 => Pw(12)(63*8-1 downto 62*8), w64 => Pw(12)(64*8-1 downto 63*8), 
w65 => Pw(12)( 65*8-1 downto  64*8), w66 => Pw(12)( 66*8-1 downto  65*8), w67 => Pw(12)( 67*8-1 downto  66*8), w68 => Pw(12)( 68*8-1 downto  67*8), w69 => Pw(12)( 69*8-1 downto  68*8), w70 => Pw(12)( 70*8-1 downto  69*8), w71 => Pw(12)( 71*8-1 downto  70*8), w72 => Pw(12)( 72*8-1 downto  71*8), 
w73 => Pw(12)( 73*8-1 downto  72*8), w74 => Pw(12)( 74*8-1 downto  73*8), w75 => Pw(12)( 75*8-1 downto  74*8), w76 => Pw(12)( 76*8-1 downto  75*8), w77 => Pw(12)( 77*8-1 downto  76*8), w78 => Pw(12)( 78*8-1 downto  77*8), w79 => Pw(12)( 79*8-1 downto  78*8), w80 => Pw(12)( 80*8-1 downto  79*8), 
w81 => Pw(12)( 81*8-1 downto  80*8), w82 => Pw(12)( 82*8-1 downto  81*8), w83 => Pw(12)( 83*8-1 downto  82*8), w84 => Pw(12)( 84*8-1 downto  83*8), w85 => Pw(12)( 85*8-1 downto  84*8), w86 => Pw(12)( 86*8-1 downto  85*8), w87 => Pw(12)( 87*8-1 downto  86*8), w88 => Pw(12)( 88*8-1 downto  87*8), 
w89 => Pw(12)( 89*8-1 downto  88*8), w90 => Pw(12)( 90*8-1 downto  89*8), w91 => Pw(12)( 91*8-1 downto  90*8), w92 => Pw(12)( 92*8-1 downto  91*8), w93 => Pw(12)( 93*8-1 downto  92*8), w94 => Pw(12)( 94*8-1 downto  93*8), w95 => Pw(12)( 95*8-1 downto  94*8), w96 => Pw(12)( 96*8-1 downto  95*8), 
w97 => Pw(12)( 97*8-1 downto  96*8), w98 => Pw(12)( 98*8-1 downto  97*8), w99 => Pw(12)( 99*8-1 downto  98*8), w100=> Pw(12)(100*8-1 downto  99*8), w101=> Pw(12)(101*8-1 downto 100*8), w102=> Pw(12)(102*8-1 downto 101*8), w103=> Pw(12)(103*8-1 downto 102*8), w104=> Pw(12)(104*8-1 downto 103*8), 
w105=> Pw(12)(105*8-1 downto 104*8), w106=> Pw(12)(106*8-1 downto 105*8), w107=> Pw(12)(107*8-1 downto 106*8), w108=> Pw(12)(108*8-1 downto 107*8), w109=> Pw(12)(109*8-1 downto 108*8), w110=> Pw(12)(110*8-1 downto 109*8), w111=> Pw(12)(111*8-1 downto 110*8), w112=> Pw(12)(112*8-1 downto 111*8), 
w113=> Pw(12)(113*8-1 downto 112*8), w114=> Pw(12)(114*8-1 downto 113*8), w115=> Pw(12)(115*8-1 downto 114*8), w116=> Pw(12)(116*8-1 downto 115*8), w117=> Pw(12)(117*8-1 downto 116*8), w118=> Pw(12)(118*8-1 downto 117*8), w119=> Pw(12)(119*8-1 downto 118*8), w120=> Pw(12)(120*8-1 downto 119*8), 
w121=> Pw(12)(121*8-1 downto 120*8), w122=> Pw(12)(122*8-1 downto 121*8), w123=> Pw(12)(123*8-1 downto 122*8), w124=> Pw(12)(124*8-1 downto 123*8), w125=> Pw(12)(125*8-1 downto 124*8), w126=> Pw(12)(126*8-1 downto 125*8), w127=> Pw(12)(127*8-1 downto 126*8), w128=> Pw(12)(128*8-1 downto 127*8), 

           d_out   => pca_d12_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_13_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(13)(     7 downto    0), w02 => Pw(13)( 2*8-1 downto    8), w03 => Pw(13)( 3*8-1 downto  2*8), w04 => Pw(13)( 4*8-1 downto  3*8), w05 => Pw(13)( 5*8-1 downto  4*8), w06 => Pw(13)( 6*8-1 downto  5*8), w07 => Pw(13)( 7*8-1 downto  6*8), w08 => Pw(13)( 8*8-1 downto  7*8),  
w09 => Pw(13)( 9*8-1 downto  8*8), w10 => Pw(13)(10*8-1 downto  9*8), w11 => Pw(13)(11*8-1 downto 10*8), w12 => Pw(13)(12*8-1 downto 11*8), w13 => Pw(13)(13*8-1 downto 12*8), w14 => Pw(13)(14*8-1 downto 13*8), w15 => Pw(13)(15*8-1 downto 14*8), w16 => Pw(13)(16*8-1 downto 15*8),  
w17 => Pw(13)(17*8-1 downto 16*8), w18 => Pw(13)(18*8-1 downto 17*8), w19 => Pw(13)(19*8-1 downto 18*8), w20 => Pw(13)(20*8-1 downto 19*8), w21 => Pw(13)(21*8-1 downto 20*8), w22 => Pw(13)(22*8-1 downto 21*8), w23 => Pw(13)(23*8-1 downto 22*8), w24 => Pw(13)(24*8-1 downto 23*8),  
w25 => Pw(13)(25*8-1 downto 24*8), w26 => Pw(13)(26*8-1 downto 25*8), w27 => Pw(13)(27*8-1 downto 26*8), w28 => Pw(13)(28*8-1 downto 27*8), w29 => Pw(13)(29*8-1 downto 28*8), w30 => Pw(13)(30*8-1 downto 29*8), w31 => Pw(13)(31*8-1 downto 30*8), w32 => Pw(13)(32*8-1 downto 31*8),  
w33 => Pw(13)(33*8-1 downto 32*8), w34 => Pw(13)(34*8-1 downto 33*8), w35 => Pw(13)(35*8-1 downto 34*8), w36 => Pw(13)(36*8-1 downto 35*8), w37 => Pw(13)(37*8-1 downto 36*8), w38 => Pw(13)(38*8-1 downto 37*8), w39 => Pw(13)(39*8-1 downto 38*8), w40 => Pw(13)(40*8-1 downto 39*8),  
w41 => Pw(13)(41*8-1 downto 40*8), w42 => Pw(13)(42*8-1 downto 41*8), w43 => Pw(13)(43*8-1 downto 42*8), w44 => Pw(13)(44*8-1 downto 43*8), w45 => Pw(13)(45*8-1 downto 44*8), w46 => Pw(13)(46*8-1 downto 45*8), w47 => Pw(13)(47*8-1 downto 46*8), w48 => Pw(13)(48*8-1 downto 47*8),  
w49 => Pw(13)(49*8-1 downto 48*8), w50 => Pw(13)(50*8-1 downto 49*8), w51 => Pw(13)(51*8-1 downto 50*8), w52 => Pw(13)(52*8-1 downto 51*8), w53 => Pw(13)(53*8-1 downto 52*8), w54 => Pw(13)(54*8-1 downto 53*8), w55 => Pw(13)(55*8-1 downto 54*8), w56 => Pw(13)(56*8-1 downto 55*8),  
w57 => Pw(13)(57*8-1 downto 56*8), w58 => Pw(13)(58*8-1 downto 57*8), w59 => Pw(13)(59*8-1 downto 58*8), w60 => Pw(13)(60*8-1 downto 59*8), w61 => Pw(13)(61*8-1 downto 60*8), w62 => Pw(13)(62*8-1 downto 61*8), w63 => Pw(13)(63*8-1 downto 62*8), w64 => Pw(13)(64*8-1 downto 63*8), 
w65 => Pw(13)( 65*8-1 downto  64*8), w66 => Pw(13)( 66*8-1 downto  65*8), w67 => Pw(13)( 67*8-1 downto  66*8), w68 => Pw(13)( 68*8-1 downto  67*8), w69 => Pw(13)( 69*8-1 downto  68*8), w70 => Pw(13)( 70*8-1 downto  69*8), w71 => Pw(13)( 71*8-1 downto  70*8), w72 => Pw(13)( 72*8-1 downto  71*8), 
w73 => Pw(13)( 73*8-1 downto  72*8), w74 => Pw(13)( 74*8-1 downto  73*8), w75 => Pw(13)( 75*8-1 downto  74*8), w76 => Pw(13)( 76*8-1 downto  75*8), w77 => Pw(13)( 77*8-1 downto  76*8), w78 => Pw(13)( 78*8-1 downto  77*8), w79 => Pw(13)( 79*8-1 downto  78*8), w80 => Pw(13)( 80*8-1 downto  79*8), 
w81 => Pw(13)( 81*8-1 downto  80*8), w82 => Pw(13)( 82*8-1 downto  81*8), w83 => Pw(13)( 83*8-1 downto  82*8), w84 => Pw(13)( 84*8-1 downto  83*8), w85 => Pw(13)( 85*8-1 downto  84*8), w86 => Pw(13)( 86*8-1 downto  85*8), w87 => Pw(13)( 87*8-1 downto  86*8), w88 => Pw(13)( 88*8-1 downto  87*8), 
w89 => Pw(13)( 89*8-1 downto  88*8), w90 => Pw(13)( 90*8-1 downto  89*8), w91 => Pw(13)( 91*8-1 downto  90*8), w92 => Pw(13)( 92*8-1 downto  91*8), w93 => Pw(13)( 93*8-1 downto  92*8), w94 => Pw(13)( 94*8-1 downto  93*8), w95 => Pw(13)( 95*8-1 downto  94*8), w96 => Pw(13)( 96*8-1 downto  95*8), 
w97 => Pw(13)( 97*8-1 downto  96*8), w98 => Pw(13)( 98*8-1 downto  97*8), w99 => Pw(13)( 99*8-1 downto  98*8), w100=> Pw(13)(100*8-1 downto  99*8), w101=> Pw(13)(101*8-1 downto 100*8), w102=> Pw(13)(102*8-1 downto 101*8), w103=> Pw(13)(103*8-1 downto 102*8), w104=> Pw(13)(104*8-1 downto 103*8), 
w105=> Pw(13)(105*8-1 downto 104*8), w106=> Pw(13)(106*8-1 downto 105*8), w107=> Pw(13)(107*8-1 downto 106*8), w108=> Pw(13)(108*8-1 downto 107*8), w109=> Pw(13)(109*8-1 downto 108*8), w110=> Pw(13)(110*8-1 downto 109*8), w111=> Pw(13)(111*8-1 downto 110*8), w112=> Pw(13)(112*8-1 downto 111*8), 
w113=> Pw(13)(113*8-1 downto 112*8), w114=> Pw(13)(114*8-1 downto 113*8), w115=> Pw(13)(115*8-1 downto 114*8), w116=> Pw(13)(116*8-1 downto 115*8), w117=> Pw(13)(117*8-1 downto 116*8), w118=> Pw(13)(118*8-1 downto 117*8), w119=> Pw(13)(119*8-1 downto 118*8), w120=> Pw(13)(120*8-1 downto 119*8), 
w121=> Pw(13)(121*8-1 downto 120*8), w122=> Pw(13)(122*8-1 downto 121*8), w123=> Pw(13)(123*8-1 downto 122*8), w124=> Pw(13)(124*8-1 downto 123*8), w125=> Pw(13)(125*8-1 downto 124*8), w126=> Pw(13)(126*8-1 downto 125*8), w127=> Pw(13)(127*8-1 downto 126*8), w128=> Pw(13)(128*8-1 downto 127*8), 

           d_out   => pca_d13_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_14_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(14)(     7 downto    0), w02 => Pw(14)( 2*8-1 downto    8), w03 => Pw(14)( 3*8-1 downto  2*8), w04 => Pw(14)( 4*8-1 downto  3*8), w05 => Pw(14)( 5*8-1 downto  4*8), w06 => Pw(14)( 6*8-1 downto  5*8), w07 => Pw(14)( 7*8-1 downto  6*8), w08 => Pw(14)( 8*8-1 downto  7*8),  
w09 => Pw(14)( 9*8-1 downto  8*8), w10 => Pw(14)(10*8-1 downto  9*8), w11 => Pw(14)(11*8-1 downto 10*8), w12 => Pw(14)(12*8-1 downto 11*8), w13 => Pw(14)(13*8-1 downto 12*8), w14 => Pw(14)(14*8-1 downto 13*8), w15 => Pw(14)(15*8-1 downto 14*8), w16 => Pw(14)(16*8-1 downto 15*8),  
w17 => Pw(14)(17*8-1 downto 16*8), w18 => Pw(14)(18*8-1 downto 17*8), w19 => Pw(14)(19*8-1 downto 18*8), w20 => Pw(14)(20*8-1 downto 19*8), w21 => Pw(14)(21*8-1 downto 20*8), w22 => Pw(14)(22*8-1 downto 21*8), w23 => Pw(14)(23*8-1 downto 22*8), w24 => Pw(14)(24*8-1 downto 23*8),  
w25 => Pw(14)(25*8-1 downto 24*8), w26 => Pw(14)(26*8-1 downto 25*8), w27 => Pw(14)(27*8-1 downto 26*8), w28 => Pw(14)(28*8-1 downto 27*8), w29 => Pw(14)(29*8-1 downto 28*8), w30 => Pw(14)(30*8-1 downto 29*8), w31 => Pw(14)(31*8-1 downto 30*8), w32 => Pw(14)(32*8-1 downto 31*8),  
w33 => Pw(14)(33*8-1 downto 32*8), w34 => Pw(14)(34*8-1 downto 33*8), w35 => Pw(14)(35*8-1 downto 34*8), w36 => Pw(14)(36*8-1 downto 35*8), w37 => Pw(14)(37*8-1 downto 36*8), w38 => Pw(14)(38*8-1 downto 37*8), w39 => Pw(14)(39*8-1 downto 38*8), w40 => Pw(14)(40*8-1 downto 39*8),  
w41 => Pw(14)(41*8-1 downto 40*8), w42 => Pw(14)(42*8-1 downto 41*8), w43 => Pw(14)(43*8-1 downto 42*8), w44 => Pw(14)(44*8-1 downto 43*8), w45 => Pw(14)(45*8-1 downto 44*8), w46 => Pw(14)(46*8-1 downto 45*8), w47 => Pw(14)(47*8-1 downto 46*8), w48 => Pw(14)(48*8-1 downto 47*8),  
w49 => Pw(14)(49*8-1 downto 48*8), w50 => Pw(14)(50*8-1 downto 49*8), w51 => Pw(14)(51*8-1 downto 50*8), w52 => Pw(14)(52*8-1 downto 51*8), w53 => Pw(14)(53*8-1 downto 52*8), w54 => Pw(14)(54*8-1 downto 53*8), w55 => Pw(14)(55*8-1 downto 54*8), w56 => Pw(14)(56*8-1 downto 55*8),  
w57 => Pw(14)(57*8-1 downto 56*8), w58 => Pw(14)(58*8-1 downto 57*8), w59 => Pw(14)(59*8-1 downto 58*8), w60 => Pw(14)(60*8-1 downto 59*8), w61 => Pw(14)(61*8-1 downto 60*8), w62 => Pw(14)(62*8-1 downto 61*8), w63 => Pw(14)(63*8-1 downto 62*8), w64 => Pw(14)(64*8-1 downto 63*8), 
w65 => Pw(14)( 65*8-1 downto  64*8), w66 => Pw(14)( 66*8-1 downto  65*8), w67 => Pw(14)( 67*8-1 downto  66*8), w68 => Pw(14)( 68*8-1 downto  67*8), w69 => Pw(14)( 69*8-1 downto  68*8), w70 => Pw(14)( 70*8-1 downto  69*8), w71 => Pw(14)( 71*8-1 downto  70*8), w72 => Pw(14)( 72*8-1 downto  71*8), 
w73 => Pw(14)( 73*8-1 downto  72*8), w74 => Pw(14)( 74*8-1 downto  73*8), w75 => Pw(14)( 75*8-1 downto  74*8), w76 => Pw(14)( 76*8-1 downto  75*8), w77 => Pw(14)( 77*8-1 downto  76*8), w78 => Pw(14)( 78*8-1 downto  77*8), w79 => Pw(14)( 79*8-1 downto  78*8), w80 => Pw(14)( 80*8-1 downto  79*8), 
w81 => Pw(14)( 81*8-1 downto  80*8), w82 => Pw(14)( 82*8-1 downto  81*8), w83 => Pw(14)( 83*8-1 downto  82*8), w84 => Pw(14)( 84*8-1 downto  83*8), w85 => Pw(14)( 85*8-1 downto  84*8), w86 => Pw(14)( 86*8-1 downto  85*8), w87 => Pw(14)( 87*8-1 downto  86*8), w88 => Pw(14)( 88*8-1 downto  87*8), 
w89 => Pw(14)( 89*8-1 downto  88*8), w90 => Pw(14)( 90*8-1 downto  89*8), w91 => Pw(14)( 91*8-1 downto  90*8), w92 => Pw(14)( 92*8-1 downto  91*8), w93 => Pw(14)( 93*8-1 downto  92*8), w94 => Pw(14)( 94*8-1 downto  93*8), w95 => Pw(14)( 95*8-1 downto  94*8), w96 => Pw(14)( 96*8-1 downto  95*8), 
w97 => Pw(14)( 97*8-1 downto  96*8), w98 => Pw(14)( 98*8-1 downto  97*8), w99 => Pw(14)( 99*8-1 downto  98*8), w100=> Pw(14)(100*8-1 downto  99*8), w101=> Pw(14)(101*8-1 downto 100*8), w102=> Pw(14)(102*8-1 downto 101*8), w103=> Pw(14)(103*8-1 downto 102*8), w104=> Pw(14)(104*8-1 downto 103*8), 
w105=> Pw(14)(105*8-1 downto 104*8), w106=> Pw(14)(106*8-1 downto 105*8), w107=> Pw(14)(107*8-1 downto 106*8), w108=> Pw(14)(108*8-1 downto 107*8), w109=> Pw(14)(109*8-1 downto 108*8), w110=> Pw(14)(110*8-1 downto 109*8), w111=> Pw(14)(111*8-1 downto 110*8), w112=> Pw(14)(112*8-1 downto 111*8), 
w113=> Pw(14)(113*8-1 downto 112*8), w114=> Pw(14)(114*8-1 downto 113*8), w115=> Pw(14)(115*8-1 downto 114*8), w116=> Pw(14)(116*8-1 downto 115*8), w117=> Pw(14)(117*8-1 downto 116*8), w118=> Pw(14)(118*8-1 downto 117*8), w119=> Pw(14)(119*8-1 downto 118*8), w120=> Pw(14)(120*8-1 downto 119*8), 
w121=> Pw(14)(121*8-1 downto 120*8), w122=> Pw(14)(122*8-1 downto 121*8), w123=> Pw(14)(123*8-1 downto 122*8), w124=> Pw(14)(124*8-1 downto 123*8), w125=> Pw(14)(125*8-1 downto 124*8), w126=> Pw(14)(126*8-1 downto 125*8), w127=> Pw(14)(127*8-1 downto 126*8), w128=> Pw(14)(128*8-1 downto 127*8), 

           d_out   => pca_d14_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_15_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(15)(     7 downto    0), w02 => Pw(15)( 2*8-1 downto    8), w03 => Pw(15)( 3*8-1 downto  2*8), w04 => Pw(15)( 4*8-1 downto  3*8), w05 => Pw(15)( 5*8-1 downto  4*8), w06 => Pw(15)( 6*8-1 downto  5*8), w07 => Pw(15)( 7*8-1 downto  6*8), w08 => Pw(15)( 8*8-1 downto  7*8),  
w09 => Pw(15)( 9*8-1 downto  8*8), w10 => Pw(15)(10*8-1 downto  9*8), w11 => Pw(15)(11*8-1 downto 10*8), w12 => Pw(15)(12*8-1 downto 11*8), w13 => Pw(15)(13*8-1 downto 12*8), w14 => Pw(15)(14*8-1 downto 13*8), w15 => Pw(15)(15*8-1 downto 14*8), w16 => Pw(15)(16*8-1 downto 15*8),  
w17 => Pw(15)(17*8-1 downto 16*8), w18 => Pw(15)(18*8-1 downto 17*8), w19 => Pw(15)(19*8-1 downto 18*8), w20 => Pw(15)(20*8-1 downto 19*8), w21 => Pw(15)(21*8-1 downto 20*8), w22 => Pw(15)(22*8-1 downto 21*8), w23 => Pw(15)(23*8-1 downto 22*8), w24 => Pw(15)(24*8-1 downto 23*8),  
w25 => Pw(15)(25*8-1 downto 24*8), w26 => Pw(15)(26*8-1 downto 25*8), w27 => Pw(15)(27*8-1 downto 26*8), w28 => Pw(15)(28*8-1 downto 27*8), w29 => Pw(15)(29*8-1 downto 28*8), w30 => Pw(15)(30*8-1 downto 29*8), w31 => Pw(15)(31*8-1 downto 30*8), w32 => Pw(15)(32*8-1 downto 31*8),  
w33 => Pw(15)(33*8-1 downto 32*8), w34 => Pw(15)(34*8-1 downto 33*8), w35 => Pw(15)(35*8-1 downto 34*8), w36 => Pw(15)(36*8-1 downto 35*8), w37 => Pw(15)(37*8-1 downto 36*8), w38 => Pw(15)(38*8-1 downto 37*8), w39 => Pw(15)(39*8-1 downto 38*8), w40 => Pw(15)(40*8-1 downto 39*8),  
w41 => Pw(15)(41*8-1 downto 40*8), w42 => Pw(15)(42*8-1 downto 41*8), w43 => Pw(15)(43*8-1 downto 42*8), w44 => Pw(15)(44*8-1 downto 43*8), w45 => Pw(15)(45*8-1 downto 44*8), w46 => Pw(15)(46*8-1 downto 45*8), w47 => Pw(15)(47*8-1 downto 46*8), w48 => Pw(15)(48*8-1 downto 47*8),  
w49 => Pw(15)(49*8-1 downto 48*8), w50 => Pw(15)(50*8-1 downto 49*8), w51 => Pw(15)(51*8-1 downto 50*8), w52 => Pw(15)(52*8-1 downto 51*8), w53 => Pw(15)(53*8-1 downto 52*8), w54 => Pw(15)(54*8-1 downto 53*8), w55 => Pw(15)(55*8-1 downto 54*8), w56 => Pw(15)(56*8-1 downto 55*8),  
w57 => Pw(15)(57*8-1 downto 56*8), w58 => Pw(15)(58*8-1 downto 57*8), w59 => Pw(15)(59*8-1 downto 58*8), w60 => Pw(15)(60*8-1 downto 59*8), w61 => Pw(15)(61*8-1 downto 60*8), w62 => Pw(15)(62*8-1 downto 61*8), w63 => Pw(15)(63*8-1 downto 62*8), w64 => Pw(15)(64*8-1 downto 63*8), 
w65 => Pw(15)( 65*8-1 downto  64*8), w66 => Pw(15)( 66*8-1 downto  65*8), w67 => Pw(15)( 67*8-1 downto  66*8), w68 => Pw(15)( 68*8-1 downto  67*8), w69 => Pw(15)( 69*8-1 downto  68*8), w70 => Pw(15)( 70*8-1 downto  69*8), w71 => Pw(15)( 71*8-1 downto  70*8), w72 => Pw(15)( 72*8-1 downto  71*8), 
w73 => Pw(15)( 73*8-1 downto  72*8), w74 => Pw(15)( 74*8-1 downto  73*8), w75 => Pw(15)( 75*8-1 downto  74*8), w76 => Pw(15)( 76*8-1 downto  75*8), w77 => Pw(15)( 77*8-1 downto  76*8), w78 => Pw(15)( 78*8-1 downto  77*8), w79 => Pw(15)( 79*8-1 downto  78*8), w80 => Pw(15)( 80*8-1 downto  79*8), 
w81 => Pw(15)( 81*8-1 downto  80*8), w82 => Pw(15)( 82*8-1 downto  81*8), w83 => Pw(15)( 83*8-1 downto  82*8), w84 => Pw(15)( 84*8-1 downto  83*8), w85 => Pw(15)( 85*8-1 downto  84*8), w86 => Pw(15)( 86*8-1 downto  85*8), w87 => Pw(15)( 87*8-1 downto  86*8), w88 => Pw(15)( 88*8-1 downto  87*8), 
w89 => Pw(15)( 89*8-1 downto  88*8), w90 => Pw(15)( 90*8-1 downto  89*8), w91 => Pw(15)( 91*8-1 downto  90*8), w92 => Pw(15)( 92*8-1 downto  91*8), w93 => Pw(15)( 93*8-1 downto  92*8), w94 => Pw(15)( 94*8-1 downto  93*8), w95 => Pw(15)( 95*8-1 downto  94*8), w96 => Pw(15)( 96*8-1 downto  95*8), 
w97 => Pw(15)( 97*8-1 downto  96*8), w98 => Pw(15)( 98*8-1 downto  97*8), w99 => Pw(15)( 99*8-1 downto  98*8), w100=> Pw(15)(100*8-1 downto  99*8), w101=> Pw(15)(101*8-1 downto 100*8), w102=> Pw(15)(102*8-1 downto 101*8), w103=> Pw(15)(103*8-1 downto 102*8), w104=> Pw(15)(104*8-1 downto 103*8), 
w105=> Pw(15)(105*8-1 downto 104*8), w106=> Pw(15)(106*8-1 downto 105*8), w107=> Pw(15)(107*8-1 downto 106*8), w108=> Pw(15)(108*8-1 downto 107*8), w109=> Pw(15)(109*8-1 downto 108*8), w110=> Pw(15)(110*8-1 downto 109*8), w111=> Pw(15)(111*8-1 downto 110*8), w112=> Pw(15)(112*8-1 downto 111*8), 
w113=> Pw(15)(113*8-1 downto 112*8), w114=> Pw(15)(114*8-1 downto 113*8), w115=> Pw(15)(115*8-1 downto 114*8), w116=> Pw(15)(116*8-1 downto 115*8), w117=> Pw(15)(117*8-1 downto 116*8), w118=> Pw(15)(118*8-1 downto 117*8), w119=> Pw(15)(119*8-1 downto 118*8), w120=> Pw(15)(120*8-1 downto 119*8), 
w121=> Pw(15)(121*8-1 downto 120*8), w122=> Pw(15)(122*8-1 downto 121*8), w123=> Pw(15)(123*8-1 downto 122*8), w124=> Pw(15)(124*8-1 downto 123*8), w125=> Pw(15)(125*8-1 downto 124*8), w126=> Pw(15)(126*8-1 downto 125*8), w127=> Pw(15)(127*8-1 downto 126*8), w128=> Pw(15)(128*8-1 downto 127*8), 

           d_out   => pca_d15_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_16_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(16)(     7 downto    0), w02 => Pw(16)( 2*8-1 downto    8), w03 => Pw(16)( 3*8-1 downto  2*8), w04 => Pw(16)( 4*8-1 downto  3*8), w05 => Pw(16)( 5*8-1 downto  4*8), w06 => Pw(16)( 6*8-1 downto  5*8), w07 => Pw(16)( 7*8-1 downto  6*8), w08 => Pw(16)( 8*8-1 downto  7*8),  
w09 => Pw(16)( 9*8-1 downto  8*8), w10 => Pw(16)(10*8-1 downto  9*8), w11 => Pw(16)(11*8-1 downto 10*8), w12 => Pw(16)(12*8-1 downto 11*8), w13 => Pw(16)(13*8-1 downto 12*8), w14 => Pw(16)(14*8-1 downto 13*8), w15 => Pw(16)(15*8-1 downto 14*8), w16 => Pw(16)(16*8-1 downto 15*8),  
w17 => Pw(16)(17*8-1 downto 16*8), w18 => Pw(16)(18*8-1 downto 17*8), w19 => Pw(16)(19*8-1 downto 18*8), w20 => Pw(16)(20*8-1 downto 19*8), w21 => Pw(16)(21*8-1 downto 20*8), w22 => Pw(16)(22*8-1 downto 21*8), w23 => Pw(16)(23*8-1 downto 22*8), w24 => Pw(16)(24*8-1 downto 23*8),  
w25 => Pw(16)(25*8-1 downto 24*8), w26 => Pw(16)(26*8-1 downto 25*8), w27 => Pw(16)(27*8-1 downto 26*8), w28 => Pw(16)(28*8-1 downto 27*8), w29 => Pw(16)(29*8-1 downto 28*8), w30 => Pw(16)(30*8-1 downto 29*8), w31 => Pw(16)(31*8-1 downto 30*8), w32 => Pw(16)(32*8-1 downto 31*8),  
w33 => Pw(16)(33*8-1 downto 32*8), w34 => Pw(16)(34*8-1 downto 33*8), w35 => Pw(16)(35*8-1 downto 34*8), w36 => Pw(16)(36*8-1 downto 35*8), w37 => Pw(16)(37*8-1 downto 36*8), w38 => Pw(16)(38*8-1 downto 37*8), w39 => Pw(16)(39*8-1 downto 38*8), w40 => Pw(16)(40*8-1 downto 39*8),  
w41 => Pw(16)(41*8-1 downto 40*8), w42 => Pw(16)(42*8-1 downto 41*8), w43 => Pw(16)(43*8-1 downto 42*8), w44 => Pw(16)(44*8-1 downto 43*8), w45 => Pw(16)(45*8-1 downto 44*8), w46 => Pw(16)(46*8-1 downto 45*8), w47 => Pw(16)(47*8-1 downto 46*8), w48 => Pw(16)(48*8-1 downto 47*8),  
w49 => Pw(16)(49*8-1 downto 48*8), w50 => Pw(16)(50*8-1 downto 49*8), w51 => Pw(16)(51*8-1 downto 50*8), w52 => Pw(16)(52*8-1 downto 51*8), w53 => Pw(16)(53*8-1 downto 52*8), w54 => Pw(16)(54*8-1 downto 53*8), w55 => Pw(16)(55*8-1 downto 54*8), w56 => Pw(16)(56*8-1 downto 55*8),  
w57 => Pw(16)(57*8-1 downto 56*8), w58 => Pw(16)(58*8-1 downto 57*8), w59 => Pw(16)(59*8-1 downto 58*8), w60 => Pw(16)(60*8-1 downto 59*8), w61 => Pw(16)(61*8-1 downto 60*8), w62 => Pw(16)(62*8-1 downto 61*8), w63 => Pw(16)(63*8-1 downto 62*8), w64 => Pw(16)(64*8-1 downto 63*8), 
w65 => Pw(16)( 65*8-1 downto  64*8), w66 => Pw(16)( 66*8-1 downto  65*8), w67 => Pw(16)( 67*8-1 downto  66*8), w68 => Pw(16)( 68*8-1 downto  67*8), w69 => Pw(16)( 69*8-1 downto  68*8), w70 => Pw(16)( 70*8-1 downto  69*8), w71 => Pw(16)( 71*8-1 downto  70*8), w72 => Pw(16)( 72*8-1 downto  71*8), 
w73 => Pw(16)( 73*8-1 downto  72*8), w74 => Pw(16)( 74*8-1 downto  73*8), w75 => Pw(16)( 75*8-1 downto  74*8), w76 => Pw(16)( 76*8-1 downto  75*8), w77 => Pw(16)( 77*8-1 downto  76*8), w78 => Pw(16)( 78*8-1 downto  77*8), w79 => Pw(16)( 79*8-1 downto  78*8), w80 => Pw(16)( 80*8-1 downto  79*8), 
w81 => Pw(16)( 81*8-1 downto  80*8), w82 => Pw(16)( 82*8-1 downto  81*8), w83 => Pw(16)( 83*8-1 downto  82*8), w84 => Pw(16)( 84*8-1 downto  83*8), w85 => Pw(16)( 85*8-1 downto  84*8), w86 => Pw(16)( 86*8-1 downto  85*8), w87 => Pw(16)( 87*8-1 downto  86*8), w88 => Pw(16)( 88*8-1 downto  87*8), 
w89 => Pw(16)( 89*8-1 downto  88*8), w90 => Pw(16)( 90*8-1 downto  89*8), w91 => Pw(16)( 91*8-1 downto  90*8), w92 => Pw(16)( 92*8-1 downto  91*8), w93 => Pw(16)( 93*8-1 downto  92*8), w94 => Pw(16)( 94*8-1 downto  93*8), w95 => Pw(16)( 95*8-1 downto  94*8), w96 => Pw(16)( 96*8-1 downto  95*8), 
w97 => Pw(16)( 97*8-1 downto  96*8), w98 => Pw(16)( 98*8-1 downto  97*8), w99 => Pw(16)( 99*8-1 downto  98*8), w100=> Pw(16)(100*8-1 downto  99*8), w101=> Pw(16)(101*8-1 downto 100*8), w102=> Pw(16)(102*8-1 downto 101*8), w103=> Pw(16)(103*8-1 downto 102*8), w104=> Pw(16)(104*8-1 downto 103*8), 
w105=> Pw(16)(105*8-1 downto 104*8), w106=> Pw(16)(106*8-1 downto 105*8), w107=> Pw(16)(107*8-1 downto 106*8), w108=> Pw(16)(108*8-1 downto 107*8), w109=> Pw(16)(109*8-1 downto 108*8), w110=> Pw(16)(110*8-1 downto 109*8), w111=> Pw(16)(111*8-1 downto 110*8), w112=> Pw(16)(112*8-1 downto 111*8), 
w113=> Pw(16)(113*8-1 downto 112*8), w114=> Pw(16)(114*8-1 downto 113*8), w115=> Pw(16)(115*8-1 downto 114*8), w116=> Pw(16)(116*8-1 downto 115*8), w117=> Pw(16)(117*8-1 downto 116*8), w118=> Pw(16)(118*8-1 downto 117*8), w119=> Pw(16)(119*8-1 downto 118*8), w120=> Pw(16)(120*8-1 downto 119*8), 
w121=> Pw(16)(121*8-1 downto 120*8), w122=> Pw(16)(122*8-1 downto 121*8), w123=> Pw(16)(123*8-1 downto 122*8), w124=> Pw(16)(124*8-1 downto 123*8), w125=> Pw(16)(125*8-1 downto 124*8), w126=> Pw(16)(126*8-1 downto 125*8), w127=> Pw(16)(127*8-1 downto 126*8), w128=> Pw(16)(128*8-1 downto 127*8), 

           d_out   => pca_d16_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_17_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out, 

w01 => Pw(17)(     7 downto    0), w02 => Pw(17)( 2*8-1 downto    8), w03 => Pw(17)( 3*8-1 downto  2*8), w04 => Pw(17)( 4*8-1 downto  3*8), w05 => Pw(17)( 5*8-1 downto  4*8), w06 => Pw(17)( 6*8-1 downto  5*8), w07 => Pw(17)( 7*8-1 downto  6*8), w08 => Pw(17)( 8*8-1 downto  7*8),  
w09 => Pw(17)( 9*8-1 downto  8*8), w10 => Pw(17)(10*8-1 downto  9*8), w11 => Pw(17)(11*8-1 downto 10*8), w12 => Pw(17)(12*8-1 downto 11*8), w13 => Pw(17)(13*8-1 downto 12*8), w14 => Pw(17)(14*8-1 downto 13*8), w15 => Pw(17)(15*8-1 downto 14*8), w16 => Pw(17)(16*8-1 downto 15*8),  
w17 => Pw(17)(17*8-1 downto 16*8), w18 => Pw(17)(18*8-1 downto 17*8), w19 => Pw(17)(19*8-1 downto 18*8), w20 => Pw(17)(20*8-1 downto 19*8), w21 => Pw(17)(21*8-1 downto 20*8), w22 => Pw(17)(22*8-1 downto 21*8), w23 => Pw(17)(23*8-1 downto 22*8), w24 => Pw(17)(24*8-1 downto 23*8),  
w25 => Pw(17)(25*8-1 downto 24*8), w26 => Pw(17)(26*8-1 downto 25*8), w27 => Pw(17)(27*8-1 downto 26*8), w28 => Pw(17)(28*8-1 downto 27*8), w29 => Pw(17)(29*8-1 downto 28*8), w30 => Pw(17)(30*8-1 downto 29*8), w31 => Pw(17)(31*8-1 downto 30*8), w32 => Pw(17)(32*8-1 downto 31*8),  
w33 => Pw(17)(33*8-1 downto 32*8), w34 => Pw(17)(34*8-1 downto 33*8), w35 => Pw(17)(35*8-1 downto 34*8), w36 => Pw(17)(36*8-1 downto 35*8), w37 => Pw(17)(37*8-1 downto 36*8), w38 => Pw(17)(38*8-1 downto 37*8), w39 => Pw(17)(39*8-1 downto 38*8), w40 => Pw(17)(40*8-1 downto 39*8),  
w41 => Pw(17)(41*8-1 downto 40*8), w42 => Pw(17)(42*8-1 downto 41*8), w43 => Pw(17)(43*8-1 downto 42*8), w44 => Pw(17)(44*8-1 downto 43*8), w45 => Pw(17)(45*8-1 downto 44*8), w46 => Pw(17)(46*8-1 downto 45*8), w47 => Pw(17)(47*8-1 downto 46*8), w48 => Pw(17)(48*8-1 downto 47*8),  
w49 => Pw(17)(49*8-1 downto 48*8), w50 => Pw(17)(50*8-1 downto 49*8), w51 => Pw(17)(51*8-1 downto 50*8), w52 => Pw(17)(52*8-1 downto 51*8), w53 => Pw(17)(53*8-1 downto 52*8), w54 => Pw(17)(54*8-1 downto 53*8), w55 => Pw(17)(55*8-1 downto 54*8), w56 => Pw(17)(56*8-1 downto 55*8),  
w57 => Pw(17)(57*8-1 downto 56*8), w58 => Pw(17)(58*8-1 downto 57*8), w59 => Pw(17)(59*8-1 downto 58*8), w60 => Pw(17)(60*8-1 downto 59*8), w61 => Pw(17)(61*8-1 downto 60*8), w62 => Pw(17)(62*8-1 downto 61*8), w63 => Pw(17)(63*8-1 downto 62*8), w64 => Pw(17)(64*8-1 downto 63*8), 
w65 => Pw(17)( 65*8-1 downto  64*8), w66 => Pw(17)( 66*8-1 downto  65*8), w67 => Pw(17)( 67*8-1 downto  66*8), w68 => Pw(17)( 68*8-1 downto  67*8), w69 => Pw(17)( 69*8-1 downto  68*8), w70 => Pw(17)( 70*8-1 downto  69*8), w71 => Pw(17)( 71*8-1 downto  70*8), w72 => Pw(17)( 72*8-1 downto  71*8), 
w73 => Pw(17)( 73*8-1 downto  72*8), w74 => Pw(17)( 74*8-1 downto  73*8), w75 => Pw(17)( 75*8-1 downto  74*8), w76 => Pw(17)( 76*8-1 downto  75*8), w77 => Pw(17)( 77*8-1 downto  76*8), w78 => Pw(17)( 78*8-1 downto  77*8), w79 => Pw(17)( 79*8-1 downto  78*8), w80 => Pw(17)( 80*8-1 downto  79*8), 
w81 => Pw(17)( 81*8-1 downto  80*8), w82 => Pw(17)( 82*8-1 downto  81*8), w83 => Pw(17)( 83*8-1 downto  82*8), w84 => Pw(17)( 84*8-1 downto  83*8), w85 => Pw(17)( 85*8-1 downto  84*8), w86 => Pw(17)( 86*8-1 downto  85*8), w87 => Pw(17)( 87*8-1 downto  86*8), w88 => Pw(17)( 88*8-1 downto  87*8), 
w89 => Pw(17)( 89*8-1 downto  88*8), w90 => Pw(17)( 90*8-1 downto  89*8), w91 => Pw(17)( 91*8-1 downto  90*8), w92 => Pw(17)( 92*8-1 downto  91*8), w93 => Pw(17)( 93*8-1 downto  92*8), w94 => Pw(17)( 94*8-1 downto  93*8), w95 => Pw(17)( 95*8-1 downto  94*8), w96 => Pw(17)( 96*8-1 downto  95*8), 
w97 => Pw(17)( 97*8-1 downto  96*8), w98 => Pw(17)( 98*8-1 downto  97*8), w99 => Pw(17)( 99*8-1 downto  98*8), w100=> Pw(17)(100*8-1 downto  99*8), w101=> Pw(17)(101*8-1 downto 100*8), w102=> Pw(17)(102*8-1 downto 101*8), w103=> Pw(17)(103*8-1 downto 102*8), w104=> Pw(17)(104*8-1 downto 103*8), 
w105=> Pw(17)(105*8-1 downto 104*8), w106=> Pw(17)(106*8-1 downto 105*8), w107=> Pw(17)(107*8-1 downto 106*8), w108=> Pw(17)(108*8-1 downto 107*8), w109=> Pw(17)(109*8-1 downto 108*8), w110=> Pw(17)(110*8-1 downto 109*8), w111=> Pw(17)(111*8-1 downto 110*8), w112=> Pw(17)(112*8-1 downto 111*8), 
w113=> Pw(17)(113*8-1 downto 112*8), w114=> Pw(17)(114*8-1 downto 113*8), w115=> Pw(17)(115*8-1 downto 114*8), w116=> Pw(17)(116*8-1 downto 115*8), w117=> Pw(17)(117*8-1 downto 116*8), w118=> Pw(17)(118*8-1 downto 117*8), w119=> Pw(17)(119*8-1 downto 118*8), w120=> Pw(17)(120*8-1 downto 119*8), 
w121=> Pw(17)(121*8-1 downto 120*8), w122=> Pw(17)(122*8-1 downto 121*8), w123=> Pw(17)(123*8-1 downto 122*8), w124=> Pw(17)(124*8-1 downto 123*8), w125=> Pw(17)(125*8-1 downto 124*8), w126=> Pw(17)(126*8-1 downto 125*8), w127=> Pw(17)(127*8-1 downto 126*8), w128=> Pw(17)(128*8-1 downto 127*8), 

           d_out   => pca_d17_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_18_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(18)(     7 downto    0), w02 => Pw(18)( 2*8-1 downto    8), w03 => Pw(18)( 3*8-1 downto  2*8), w04 => Pw(18)( 4*8-1 downto  3*8), w05 => Pw(18)( 5*8-1 downto  4*8), w06 => Pw(18)( 6*8-1 downto  5*8), w07 => Pw(18)( 7*8-1 downto  6*8), w08 => Pw(18)( 8*8-1 downto  7*8),  
w09 => Pw(18)( 9*8-1 downto  8*8), w10 => Pw(18)(10*8-1 downto  9*8), w11 => Pw(18)(11*8-1 downto 10*8), w12 => Pw(18)(12*8-1 downto 11*8), w13 => Pw(18)(13*8-1 downto 12*8), w14 => Pw(18)(14*8-1 downto 13*8), w15 => Pw(18)(15*8-1 downto 14*8), w16 => Pw(18)(16*8-1 downto 15*8),  
w17 => Pw(18)(17*8-1 downto 16*8), w18 => Pw(18)(18*8-1 downto 17*8), w19 => Pw(18)(19*8-1 downto 18*8), w20 => Pw(18)(20*8-1 downto 19*8), w21 => Pw(18)(21*8-1 downto 20*8), w22 => Pw(18)(22*8-1 downto 21*8), w23 => Pw(18)(23*8-1 downto 22*8), w24 => Pw(18)(24*8-1 downto 23*8),  
w25 => Pw(18)(25*8-1 downto 24*8), w26 => Pw(18)(26*8-1 downto 25*8), w27 => Pw(18)(27*8-1 downto 26*8), w28 => Pw(18)(28*8-1 downto 27*8), w29 => Pw(18)(29*8-1 downto 28*8), w30 => Pw(18)(30*8-1 downto 29*8), w31 => Pw(18)(31*8-1 downto 30*8), w32 => Pw(18)(32*8-1 downto 31*8),  
w33 => Pw(18)(33*8-1 downto 32*8), w34 => Pw(18)(34*8-1 downto 33*8), w35 => Pw(18)(35*8-1 downto 34*8), w36 => Pw(18)(36*8-1 downto 35*8), w37 => Pw(18)(37*8-1 downto 36*8), w38 => Pw(18)(38*8-1 downto 37*8), w39 => Pw(18)(39*8-1 downto 38*8), w40 => Pw(18)(40*8-1 downto 39*8),  
w41 => Pw(18)(41*8-1 downto 40*8), w42 => Pw(18)(42*8-1 downto 41*8), w43 => Pw(18)(43*8-1 downto 42*8), w44 => Pw(18)(44*8-1 downto 43*8), w45 => Pw(18)(45*8-1 downto 44*8), w46 => Pw(18)(46*8-1 downto 45*8), w47 => Pw(18)(47*8-1 downto 46*8), w48 => Pw(18)(48*8-1 downto 47*8),  
w49 => Pw(18)(49*8-1 downto 48*8), w50 => Pw(18)(50*8-1 downto 49*8), w51 => Pw(18)(51*8-1 downto 50*8), w52 => Pw(18)(52*8-1 downto 51*8), w53 => Pw(18)(53*8-1 downto 52*8), w54 => Pw(18)(54*8-1 downto 53*8), w55 => Pw(18)(55*8-1 downto 54*8), w56 => Pw(18)(56*8-1 downto 55*8),  
w57 => Pw(18)(57*8-1 downto 56*8), w58 => Pw(18)(58*8-1 downto 57*8), w59 => Pw(18)(59*8-1 downto 58*8), w60 => Pw(18)(60*8-1 downto 59*8), w61 => Pw(18)(61*8-1 downto 60*8), w62 => Pw(18)(62*8-1 downto 61*8), w63 => Pw(18)(63*8-1 downto 62*8), w64 => Pw(18)(64*8-1 downto 63*8), 
w65 => Pw(18)( 65*8-1 downto  64*8), w66 => Pw(18)( 66*8-1 downto  65*8), w67 => Pw(18)( 67*8-1 downto  66*8), w68 => Pw(18)( 68*8-1 downto  67*8), w69 => Pw(18)( 69*8-1 downto  68*8), w70 => Pw(18)( 70*8-1 downto  69*8), w71 => Pw(18)( 71*8-1 downto  70*8), w72 => Pw(18)( 72*8-1 downto  71*8), 
w73 => Pw(18)( 73*8-1 downto  72*8), w74 => Pw(18)( 74*8-1 downto  73*8), w75 => Pw(18)( 75*8-1 downto  74*8), w76 => Pw(18)( 76*8-1 downto  75*8), w77 => Pw(18)( 77*8-1 downto  76*8), w78 => Pw(18)( 78*8-1 downto  77*8), w79 => Pw(18)( 79*8-1 downto  78*8), w80 => Pw(18)( 80*8-1 downto  79*8), 
w81 => Pw(18)( 81*8-1 downto  80*8), w82 => Pw(18)( 82*8-1 downto  81*8), w83 => Pw(18)( 83*8-1 downto  82*8), w84 => Pw(18)( 84*8-1 downto  83*8), w85 => Pw(18)( 85*8-1 downto  84*8), w86 => Pw(18)( 86*8-1 downto  85*8), w87 => Pw(18)( 87*8-1 downto  86*8), w88 => Pw(18)( 88*8-1 downto  87*8), 
w89 => Pw(18)( 89*8-1 downto  88*8), w90 => Pw(18)( 90*8-1 downto  89*8), w91 => Pw(18)( 91*8-1 downto  90*8), w92 => Pw(18)( 92*8-1 downto  91*8), w93 => Pw(18)( 93*8-1 downto  92*8), w94 => Pw(18)( 94*8-1 downto  93*8), w95 => Pw(18)( 95*8-1 downto  94*8), w96 => Pw(18)( 96*8-1 downto  95*8), 
w97 => Pw(18)( 97*8-1 downto  96*8), w98 => Pw(18)( 98*8-1 downto  97*8), w99 => Pw(18)( 99*8-1 downto  98*8), w100=> Pw(18)(100*8-1 downto  99*8), w101=> Pw(18)(101*8-1 downto 100*8), w102=> Pw(18)(102*8-1 downto 101*8), w103=> Pw(18)(103*8-1 downto 102*8), w104=> Pw(18)(104*8-1 downto 103*8), 
w105=> Pw(18)(105*8-1 downto 104*8), w106=> Pw(18)(106*8-1 downto 105*8), w107=> Pw(18)(107*8-1 downto 106*8), w108=> Pw(18)(108*8-1 downto 107*8), w109=> Pw(18)(109*8-1 downto 108*8), w110=> Pw(18)(110*8-1 downto 109*8), w111=> Pw(18)(111*8-1 downto 110*8), w112=> Pw(18)(112*8-1 downto 111*8), 
w113=> Pw(18)(113*8-1 downto 112*8), w114=> Pw(18)(114*8-1 downto 113*8), w115=> Pw(18)(115*8-1 downto 114*8), w116=> Pw(18)(116*8-1 downto 115*8), w117=> Pw(18)(117*8-1 downto 116*8), w118=> Pw(18)(118*8-1 downto 117*8), w119=> Pw(18)(119*8-1 downto 118*8), w120=> Pw(18)(120*8-1 downto 119*8), 
w121=> Pw(18)(121*8-1 downto 120*8), w122=> Pw(18)(122*8-1 downto 121*8), w123=> Pw(18)(123*8-1 downto 122*8), w124=> Pw(18)(124*8-1 downto 123*8), w125=> Pw(18)(125*8-1 downto 124*8), w126=> Pw(18)(126*8-1 downto 125*8), w127=> Pw(18)(127*8-1 downto 126*8), w128=> Pw(18)(128*8-1 downto 127*8), 

           d_out   => pca_d18_out   ,
           en_out  => open  ,
           sof_out => open );

  
  PCA128_19_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(19)(     7 downto    0), w02 => Pw(19)( 2*8-1 downto    8), w03 => Pw(19)( 3*8-1 downto  2*8), w04 => Pw(19)( 4*8-1 downto  3*8), w05 => Pw(19)( 5*8-1 downto  4*8), w06 => Pw(19)( 6*8-1 downto  5*8), w07 => Pw(19)( 7*8-1 downto  6*8), w08 => Pw(19)( 8*8-1 downto  7*8),  
w09 => Pw(19)( 9*8-1 downto  8*8), w10 => Pw(19)(10*8-1 downto  9*8), w11 => Pw(19)(11*8-1 downto 10*8), w12 => Pw(19)(12*8-1 downto 11*8), w13 => Pw(19)(13*8-1 downto 12*8), w14 => Pw(19)(14*8-1 downto 13*8), w15 => Pw(19)(15*8-1 downto 14*8), w16 => Pw(19)(16*8-1 downto 15*8),  
w17 => Pw(19)(17*8-1 downto 16*8), w18 => Pw(19)(18*8-1 downto 17*8), w19 => Pw(19)(19*8-1 downto 18*8), w20 => Pw(19)(20*8-1 downto 19*8), w21 => Pw(19)(21*8-1 downto 20*8), w22 => Pw(19)(22*8-1 downto 21*8), w23 => Pw(19)(23*8-1 downto 22*8), w24 => Pw(19)(24*8-1 downto 23*8),  
w25 => Pw(19)(25*8-1 downto 24*8), w26 => Pw(19)(26*8-1 downto 25*8), w27 => Pw(19)(27*8-1 downto 26*8), w28 => Pw(19)(28*8-1 downto 27*8), w29 => Pw(19)(29*8-1 downto 28*8), w30 => Pw(19)(30*8-1 downto 29*8), w31 => Pw(19)(31*8-1 downto 30*8), w32 => Pw(19)(32*8-1 downto 31*8),  
w33 => Pw(19)(33*8-1 downto 32*8), w34 => Pw(19)(34*8-1 downto 33*8), w35 => Pw(19)(35*8-1 downto 34*8), w36 => Pw(19)(36*8-1 downto 35*8), w37 => Pw(19)(37*8-1 downto 36*8), w38 => Pw(19)(38*8-1 downto 37*8), w39 => Pw(19)(39*8-1 downto 38*8), w40 => Pw(19)(40*8-1 downto 39*8),  
w41 => Pw(19)(41*8-1 downto 40*8), w42 => Pw(19)(42*8-1 downto 41*8), w43 => Pw(19)(43*8-1 downto 42*8), w44 => Pw(19)(44*8-1 downto 43*8), w45 => Pw(19)(45*8-1 downto 44*8), w46 => Pw(19)(46*8-1 downto 45*8), w47 => Pw(19)(47*8-1 downto 46*8), w48 => Pw(19)(48*8-1 downto 47*8),  
w49 => Pw(19)(49*8-1 downto 48*8), w50 => Pw(19)(50*8-1 downto 49*8), w51 => Pw(19)(51*8-1 downto 50*8), w52 => Pw(19)(52*8-1 downto 51*8), w53 => Pw(19)(53*8-1 downto 52*8), w54 => Pw(19)(54*8-1 downto 53*8), w55 => Pw(19)(55*8-1 downto 54*8), w56 => Pw(19)(56*8-1 downto 55*8),  
w57 => Pw(19)(57*8-1 downto 56*8), w58 => Pw(19)(58*8-1 downto 57*8), w59 => Pw(19)(59*8-1 downto 58*8), w60 => Pw(19)(60*8-1 downto 59*8), w61 => Pw(19)(61*8-1 downto 60*8), w62 => Pw(19)(62*8-1 downto 61*8), w63 => Pw(19)(63*8-1 downto 62*8), w64 => Pw(19)(64*8-1 downto 63*8), 
w65 => Pw(19)( 65*8-1 downto  64*8), w66 => Pw(19)( 66*8-1 downto  65*8), w67 => Pw(19)( 67*8-1 downto  66*8), w68 => Pw(19)( 68*8-1 downto  67*8), w69 => Pw(19)( 69*8-1 downto  68*8), w70 => Pw(19)( 70*8-1 downto  69*8), w71 => Pw(19)( 71*8-1 downto  70*8), w72 => Pw(19)( 72*8-1 downto  71*8), 
w73 => Pw(19)( 73*8-1 downto  72*8), w74 => Pw(19)( 74*8-1 downto  73*8), w75 => Pw(19)( 75*8-1 downto  74*8), w76 => Pw(19)( 76*8-1 downto  75*8), w77 => Pw(19)( 77*8-1 downto  76*8), w78 => Pw(19)( 78*8-1 downto  77*8), w79 => Pw(19)( 79*8-1 downto  78*8), w80 => Pw(19)( 80*8-1 downto  79*8), 
w81 => Pw(19)( 81*8-1 downto  80*8), w82 => Pw(19)( 82*8-1 downto  81*8), w83 => Pw(19)( 83*8-1 downto  82*8), w84 => Pw(19)( 84*8-1 downto  83*8), w85 => Pw(19)( 85*8-1 downto  84*8), w86 => Pw(19)( 86*8-1 downto  85*8), w87 => Pw(19)( 87*8-1 downto  86*8), w88 => Pw(19)( 88*8-1 downto  87*8), 
w89 => Pw(19)( 89*8-1 downto  88*8), w90 => Pw(19)( 90*8-1 downto  89*8), w91 => Pw(19)( 91*8-1 downto  90*8), w92 => Pw(19)( 92*8-1 downto  91*8), w93 => Pw(19)( 93*8-1 downto  92*8), w94 => Pw(19)( 94*8-1 downto  93*8), w95 => Pw(19)( 95*8-1 downto  94*8), w96 => Pw(19)( 96*8-1 downto  95*8), 
w97 => Pw(19)( 97*8-1 downto  96*8), w98 => Pw(19)( 98*8-1 downto  97*8), w99 => Pw(19)( 99*8-1 downto  98*8), w100=> Pw(19)(100*8-1 downto  99*8), w101=> Pw(19)(101*8-1 downto 100*8), w102=> Pw(19)(102*8-1 downto 101*8), w103=> Pw(19)(103*8-1 downto 102*8), w104=> Pw(19)(104*8-1 downto 103*8), 
w105=> Pw(19)(105*8-1 downto 104*8), w106=> Pw(19)(106*8-1 downto 105*8), w107=> Pw(19)(107*8-1 downto 106*8), w108=> Pw(19)(108*8-1 downto 107*8), w109=> Pw(19)(109*8-1 downto 108*8), w110=> Pw(19)(110*8-1 downto 109*8), w111=> Pw(19)(111*8-1 downto 110*8), w112=> Pw(19)(112*8-1 downto 111*8), 
w113=> Pw(19)(113*8-1 downto 112*8), w114=> Pw(19)(114*8-1 downto 113*8), w115=> Pw(19)(115*8-1 downto 114*8), w116=> Pw(19)(116*8-1 downto 115*8), w117=> Pw(19)(117*8-1 downto 116*8), w118=> Pw(19)(118*8-1 downto 117*8), w119=> Pw(19)(119*8-1 downto 118*8), w120=> Pw(19)(120*8-1 downto 119*8), 
w121=> Pw(19)(121*8-1 downto 120*8), w122=> Pw(19)(122*8-1 downto 121*8), w123=> Pw(19)(123*8-1 downto 122*8), w124=> Pw(19)(124*8-1 downto 123*8), w125=> Pw(19)(125*8-1 downto 124*8), w126=> Pw(19)(126*8-1 downto 125*8), w127=> Pw(19)(127*8-1 downto 126*8), w128=> Pw(19)(128*8-1 downto 127*8), 

           d_out   => pca_d19_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_20_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(20)(     7 downto    0), w02 => Pw(20)( 2*8-1 downto    8), w03 => Pw(20)( 3*8-1 downto  2*8), w04 => Pw(20)( 4*8-1 downto  3*8), w05 => Pw(20)( 5*8-1 downto  4*8), w06 => Pw(20)( 6*8-1 downto  5*8), w07 => Pw(20)( 7*8-1 downto  6*8), w08 => Pw(20)( 8*8-1 downto  7*8),  
w09 => Pw(20)( 9*8-1 downto  8*8), w10 => Pw(20)(10*8-1 downto  9*8), w11 => Pw(20)(11*8-1 downto 10*8), w12 => Pw(20)(12*8-1 downto 11*8), w13 => Pw(20)(13*8-1 downto 12*8), w14 => Pw(20)(14*8-1 downto 13*8), w15 => Pw(20)(15*8-1 downto 14*8), w16 => Pw(20)(16*8-1 downto 15*8),  
w17 => Pw(20)(17*8-1 downto 16*8), w18 => Pw(20)(18*8-1 downto 17*8), w19 => Pw(20)(19*8-1 downto 18*8), w20 => Pw(20)(20*8-1 downto 19*8), w21 => Pw(20)(21*8-1 downto 20*8), w22 => Pw(20)(22*8-1 downto 21*8), w23 => Pw(20)(23*8-1 downto 22*8), w24 => Pw(20)(24*8-1 downto 23*8),  
w25 => Pw(20)(25*8-1 downto 24*8), w26 => Pw(20)(26*8-1 downto 25*8), w27 => Pw(20)(27*8-1 downto 26*8), w28 => Pw(20)(28*8-1 downto 27*8), w29 => Pw(20)(29*8-1 downto 28*8), w30 => Pw(20)(30*8-1 downto 29*8), w31 => Pw(20)(31*8-1 downto 30*8), w32 => Pw(20)(32*8-1 downto 31*8),  
w33 => Pw(20)(33*8-1 downto 32*8), w34 => Pw(20)(34*8-1 downto 33*8), w35 => Pw(20)(35*8-1 downto 34*8), w36 => Pw(20)(36*8-1 downto 35*8), w37 => Pw(20)(37*8-1 downto 36*8), w38 => Pw(20)(38*8-1 downto 37*8), w39 => Pw(20)(39*8-1 downto 38*8), w40 => Pw(20)(40*8-1 downto 39*8),  
w41 => Pw(20)(41*8-1 downto 40*8), w42 => Pw(20)(42*8-1 downto 41*8), w43 => Pw(20)(43*8-1 downto 42*8), w44 => Pw(20)(44*8-1 downto 43*8), w45 => Pw(20)(45*8-1 downto 44*8), w46 => Pw(20)(46*8-1 downto 45*8), w47 => Pw(20)(47*8-1 downto 46*8), w48 => Pw(20)(48*8-1 downto 47*8),  
w49 => Pw(20)(49*8-1 downto 48*8), w50 => Pw(20)(50*8-1 downto 49*8), w51 => Pw(20)(51*8-1 downto 50*8), w52 => Pw(20)(52*8-1 downto 51*8), w53 => Pw(20)(53*8-1 downto 52*8), w54 => Pw(20)(54*8-1 downto 53*8), w55 => Pw(20)(55*8-1 downto 54*8), w56 => Pw(20)(56*8-1 downto 55*8),  
w57 => Pw(20)(57*8-1 downto 56*8), w58 => Pw(20)(58*8-1 downto 57*8), w59 => Pw(20)(59*8-1 downto 58*8), w60 => Pw(20)(60*8-1 downto 59*8), w61 => Pw(20)(61*8-1 downto 60*8), w62 => Pw(20)(62*8-1 downto 61*8), w63 => Pw(20)(63*8-1 downto 62*8), w64 => Pw(20)(64*8-1 downto 63*8), 
w65 => Pw(20)( 65*8-1 downto  64*8), w66 => Pw(20)( 66*8-1 downto  65*8), w67 => Pw(20)( 67*8-1 downto  66*8), w68 => Pw(20)( 68*8-1 downto  67*8), w69 => Pw(20)( 69*8-1 downto  68*8), w70 => Pw(20)( 70*8-1 downto  69*8), w71 => Pw(20)( 71*8-1 downto  70*8), w72 => Pw(20)( 72*8-1 downto  71*8), 
w73 => Pw(20)( 73*8-1 downto  72*8), w74 => Pw(20)( 74*8-1 downto  73*8), w75 => Pw(20)( 75*8-1 downto  74*8), w76 => Pw(20)( 76*8-1 downto  75*8), w77 => Pw(20)( 77*8-1 downto  76*8), w78 => Pw(20)( 78*8-1 downto  77*8), w79 => Pw(20)( 79*8-1 downto  78*8), w80 => Pw(20)( 80*8-1 downto  79*8), 
w81 => Pw(20)( 81*8-1 downto  80*8), w82 => Pw(20)( 82*8-1 downto  81*8), w83 => Pw(20)( 83*8-1 downto  82*8), w84 => Pw(20)( 84*8-1 downto  83*8), w85 => Pw(20)( 85*8-1 downto  84*8), w86 => Pw(20)( 86*8-1 downto  85*8), w87 => Pw(20)( 87*8-1 downto  86*8), w88 => Pw(20)( 88*8-1 downto  87*8), 
w89 => Pw(20)( 89*8-1 downto  88*8), w90 => Pw(20)( 90*8-1 downto  89*8), w91 => Pw(20)( 91*8-1 downto  90*8), w92 => Pw(20)( 92*8-1 downto  91*8), w93 => Pw(20)( 93*8-1 downto  92*8), w94 => Pw(20)( 94*8-1 downto  93*8), w95 => Pw(20)( 95*8-1 downto  94*8), w96 => Pw(20)( 96*8-1 downto  95*8), 
w97 => Pw(20)( 97*8-1 downto  96*8), w98 => Pw(20)( 98*8-1 downto  97*8), w99 => Pw(20)( 99*8-1 downto  98*8), w100=> Pw(20)(100*8-1 downto  99*8), w101=> Pw(20)(101*8-1 downto 100*8), w102=> Pw(20)(102*8-1 downto 101*8), w103=> Pw(20)(103*8-1 downto 102*8), w104=> Pw(20)(104*8-1 downto 103*8), 
w105=> Pw(20)(105*8-1 downto 104*8), w106=> Pw(20)(106*8-1 downto 105*8), w107=> Pw(20)(107*8-1 downto 106*8), w108=> Pw(20)(108*8-1 downto 107*8), w109=> Pw(20)(109*8-1 downto 108*8), w110=> Pw(20)(110*8-1 downto 109*8), w111=> Pw(20)(111*8-1 downto 110*8), w112=> Pw(20)(112*8-1 downto 111*8), 
w113=> Pw(20)(113*8-1 downto 112*8), w114=> Pw(20)(114*8-1 downto 113*8), w115=> Pw(20)(115*8-1 downto 114*8), w116=> Pw(20)(116*8-1 downto 115*8), w117=> Pw(20)(117*8-1 downto 116*8), w118=> Pw(20)(118*8-1 downto 117*8), w119=> Pw(20)(119*8-1 downto 118*8), w120=> Pw(20)(120*8-1 downto 119*8), 
w121=> Pw(20)(121*8-1 downto 120*8), w122=> Pw(20)(122*8-1 downto 121*8), w123=> Pw(20)(123*8-1 downto 122*8), w124=> Pw(20)(124*8-1 downto 123*8), w125=> Pw(20)(125*8-1 downto 124*8), w126=> Pw(20)(126*8-1 downto 125*8), w127=> Pw(20)(127*8-1 downto 126*8), w128=> Pw(20)(128*8-1 downto 127*8), 

           d_out   => pca_d20_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_21_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(21)(     7 downto    0), w02 => Pw(21)( 2*8-1 downto    8), w03 => Pw(21)( 3*8-1 downto  2*8), w04 => Pw(21)( 4*8-1 downto  3*8), w05 => Pw(21)( 5*8-1 downto  4*8), w06 => Pw(21)( 6*8-1 downto  5*8), w07 => Pw(21)( 7*8-1 downto  6*8), w08 => Pw(21)( 8*8-1 downto  7*8),  
w09 => Pw(21)( 9*8-1 downto  8*8), w10 => Pw(21)(10*8-1 downto  9*8), w11 => Pw(21)(11*8-1 downto 10*8), w12 => Pw(21)(12*8-1 downto 11*8), w13 => Pw(21)(13*8-1 downto 12*8), w14 => Pw(21)(14*8-1 downto 13*8), w15 => Pw(21)(15*8-1 downto 14*8), w16 => Pw(21)(16*8-1 downto 15*8),  
w17 => Pw(21)(17*8-1 downto 16*8), w18 => Pw(21)(18*8-1 downto 17*8), w19 => Pw(21)(19*8-1 downto 18*8), w20 => Pw(21)(20*8-1 downto 19*8), w21 => Pw(21)(21*8-1 downto 20*8), w22 => Pw(21)(22*8-1 downto 21*8), w23 => Pw(21)(23*8-1 downto 22*8), w24 => Pw(21)(24*8-1 downto 23*8),  
w25 => Pw(21)(25*8-1 downto 24*8), w26 => Pw(21)(26*8-1 downto 25*8), w27 => Pw(21)(27*8-1 downto 26*8), w28 => Pw(21)(28*8-1 downto 27*8), w29 => Pw(21)(29*8-1 downto 28*8), w30 => Pw(21)(30*8-1 downto 29*8), w31 => Pw(21)(31*8-1 downto 30*8), w32 => Pw(21)(32*8-1 downto 31*8),  
w33 => Pw(21)(33*8-1 downto 32*8), w34 => Pw(21)(34*8-1 downto 33*8), w35 => Pw(21)(35*8-1 downto 34*8), w36 => Pw(21)(36*8-1 downto 35*8), w37 => Pw(21)(37*8-1 downto 36*8), w38 => Pw(21)(38*8-1 downto 37*8), w39 => Pw(21)(39*8-1 downto 38*8), w40 => Pw(21)(40*8-1 downto 39*8),  
w41 => Pw(21)(41*8-1 downto 40*8), w42 => Pw(21)(42*8-1 downto 41*8), w43 => Pw(21)(43*8-1 downto 42*8), w44 => Pw(21)(44*8-1 downto 43*8), w45 => Pw(21)(45*8-1 downto 44*8), w46 => Pw(21)(46*8-1 downto 45*8), w47 => Pw(21)(47*8-1 downto 46*8), w48 => Pw(21)(48*8-1 downto 47*8),  
w49 => Pw(21)(49*8-1 downto 48*8), w50 => Pw(21)(50*8-1 downto 49*8), w51 => Pw(21)(51*8-1 downto 50*8), w52 => Pw(21)(52*8-1 downto 51*8), w53 => Pw(21)(53*8-1 downto 52*8), w54 => Pw(21)(54*8-1 downto 53*8), w55 => Pw(21)(55*8-1 downto 54*8), w56 => Pw(21)(56*8-1 downto 55*8),  
w57 => Pw(21)(57*8-1 downto 56*8), w58 => Pw(21)(58*8-1 downto 57*8), w59 => Pw(21)(59*8-1 downto 58*8), w60 => Pw(21)(60*8-1 downto 59*8), w61 => Pw(21)(61*8-1 downto 60*8), w62 => Pw(21)(62*8-1 downto 61*8), w63 => Pw(21)(63*8-1 downto 62*8), w64 => Pw(21)(64*8-1 downto 63*8), 
w65 => Pw(21)( 65*8-1 downto  64*8), w66 => Pw(21)( 66*8-1 downto  65*8), w67 => Pw(21)( 67*8-1 downto  66*8), w68 => Pw(21)( 68*8-1 downto  67*8), w69 => Pw(21)( 69*8-1 downto  68*8), w70 => Pw(21)( 70*8-1 downto  69*8), w71 => Pw(21)( 71*8-1 downto  70*8), w72 => Pw(21)( 72*8-1 downto  71*8), 
w73 => Pw(21)( 73*8-1 downto  72*8), w74 => Pw(21)( 74*8-1 downto  73*8), w75 => Pw(21)( 75*8-1 downto  74*8), w76 => Pw(21)( 76*8-1 downto  75*8), w77 => Pw(21)( 77*8-1 downto  76*8), w78 => Pw(21)( 78*8-1 downto  77*8), w79 => Pw(21)( 79*8-1 downto  78*8), w80 => Pw(21)( 80*8-1 downto  79*8), 
w81 => Pw(21)( 81*8-1 downto  80*8), w82 => Pw(21)( 82*8-1 downto  81*8), w83 => Pw(21)( 83*8-1 downto  82*8), w84 => Pw(21)( 84*8-1 downto  83*8), w85 => Pw(21)( 85*8-1 downto  84*8), w86 => Pw(21)( 86*8-1 downto  85*8), w87 => Pw(21)( 87*8-1 downto  86*8), w88 => Pw(21)( 88*8-1 downto  87*8), 
w89 => Pw(21)( 89*8-1 downto  88*8), w90 => Pw(21)( 90*8-1 downto  89*8), w91 => Pw(21)( 91*8-1 downto  90*8), w92 => Pw(21)( 92*8-1 downto  91*8), w93 => Pw(21)( 93*8-1 downto  92*8), w94 => Pw(21)( 94*8-1 downto  93*8), w95 => Pw(21)( 95*8-1 downto  94*8), w96 => Pw(21)( 96*8-1 downto  95*8), 
w97 => Pw(21)( 97*8-1 downto  96*8), w98 => Pw(21)( 98*8-1 downto  97*8), w99 => Pw(21)( 99*8-1 downto  98*8), w100=> Pw(21)(100*8-1 downto  99*8), w101=> Pw(21)(101*8-1 downto 100*8), w102=> Pw(21)(102*8-1 downto 101*8), w103=> Pw(21)(103*8-1 downto 102*8), w104=> Pw(21)(104*8-1 downto 103*8), 
w105=> Pw(21)(105*8-1 downto 104*8), w106=> Pw(21)(106*8-1 downto 105*8), w107=> Pw(21)(107*8-1 downto 106*8), w108=> Pw(21)(108*8-1 downto 107*8), w109=> Pw(21)(109*8-1 downto 108*8), w110=> Pw(21)(110*8-1 downto 109*8), w111=> Pw(21)(111*8-1 downto 110*8), w112=> Pw(21)(112*8-1 downto 111*8), 
w113=> Pw(21)(113*8-1 downto 112*8), w114=> Pw(21)(114*8-1 downto 113*8), w115=> Pw(21)(115*8-1 downto 114*8), w116=> Pw(21)(116*8-1 downto 115*8), w117=> Pw(21)(117*8-1 downto 116*8), w118=> Pw(21)(118*8-1 downto 117*8), w119=> Pw(21)(119*8-1 downto 118*8), w120=> Pw(21)(120*8-1 downto 119*8), 
w121=> Pw(21)(121*8-1 downto 120*8), w122=> Pw(21)(122*8-1 downto 121*8), w123=> Pw(21)(123*8-1 downto 122*8), w124=> Pw(21)(124*8-1 downto 123*8), w125=> Pw(21)(125*8-1 downto 124*8), w126=> Pw(21)(126*8-1 downto 125*8), w127=> Pw(21)(127*8-1 downto 126*8), w128=> Pw(21)(128*8-1 downto 127*8), 

           d_out   => pca_d21_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_22_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(22)(     7 downto    0), w02 => Pw(22)( 2*8-1 downto    8), w03 => Pw(22)( 3*8-1 downto  2*8), w04 => Pw(22)( 4*8-1 downto  3*8), w05 => Pw(22)( 5*8-1 downto  4*8), w06 => Pw(22)( 6*8-1 downto  5*8), w07 => Pw(22)( 7*8-1 downto  6*8), w08 => Pw(22)( 8*8-1 downto  7*8),  
w09 => Pw(22)( 9*8-1 downto  8*8), w10 => Pw(22)(10*8-1 downto  9*8), w11 => Pw(22)(11*8-1 downto 10*8), w12 => Pw(22)(12*8-1 downto 11*8), w13 => Pw(22)(13*8-1 downto 12*8), w14 => Pw(22)(14*8-1 downto 13*8), w15 => Pw(22)(15*8-1 downto 14*8), w16 => Pw(22)(16*8-1 downto 15*8),  
w17 => Pw(22)(17*8-1 downto 16*8), w18 => Pw(22)(18*8-1 downto 17*8), w19 => Pw(22)(19*8-1 downto 18*8), w20 => Pw(22)(20*8-1 downto 19*8), w21 => Pw(22)(21*8-1 downto 20*8), w22 => Pw(22)(22*8-1 downto 21*8), w23 => Pw(22)(23*8-1 downto 22*8), w24 => Pw(22)(24*8-1 downto 23*8),  
w25 => Pw(22)(25*8-1 downto 24*8), w26 => Pw(22)(26*8-1 downto 25*8), w27 => Pw(22)(27*8-1 downto 26*8), w28 => Pw(22)(28*8-1 downto 27*8), w29 => Pw(22)(29*8-1 downto 28*8), w30 => Pw(22)(30*8-1 downto 29*8), w31 => Pw(22)(31*8-1 downto 30*8), w32 => Pw(22)(32*8-1 downto 31*8),  
w33 => Pw(22)(33*8-1 downto 32*8), w34 => Pw(22)(34*8-1 downto 33*8), w35 => Pw(22)(35*8-1 downto 34*8), w36 => Pw(22)(36*8-1 downto 35*8), w37 => Pw(22)(37*8-1 downto 36*8), w38 => Pw(22)(38*8-1 downto 37*8), w39 => Pw(22)(39*8-1 downto 38*8), w40 => Pw(22)(40*8-1 downto 39*8),  
w41 => Pw(22)(41*8-1 downto 40*8), w42 => Pw(22)(42*8-1 downto 41*8), w43 => Pw(22)(43*8-1 downto 42*8), w44 => Pw(22)(44*8-1 downto 43*8), w45 => Pw(22)(45*8-1 downto 44*8), w46 => Pw(22)(46*8-1 downto 45*8), w47 => Pw(22)(47*8-1 downto 46*8), w48 => Pw(22)(48*8-1 downto 47*8),  
w49 => Pw(22)(49*8-1 downto 48*8), w50 => Pw(22)(50*8-1 downto 49*8), w51 => Pw(22)(51*8-1 downto 50*8), w52 => Pw(22)(52*8-1 downto 51*8), w53 => Pw(22)(53*8-1 downto 52*8), w54 => Pw(22)(54*8-1 downto 53*8), w55 => Pw(22)(55*8-1 downto 54*8), w56 => Pw(22)(56*8-1 downto 55*8),  
w57 => Pw(22)(57*8-1 downto 56*8), w58 => Pw(22)(58*8-1 downto 57*8), w59 => Pw(22)(59*8-1 downto 58*8), w60 => Pw(22)(60*8-1 downto 59*8), w61 => Pw(22)(61*8-1 downto 60*8), w62 => Pw(22)(62*8-1 downto 61*8), w63 => Pw(22)(63*8-1 downto 62*8), w64 => Pw(22)(64*8-1 downto 63*8), 
w65 => Pw(22)( 65*8-1 downto  64*8), w66 => Pw(22)( 66*8-1 downto  65*8), w67 => Pw(22)( 67*8-1 downto  66*8), w68 => Pw(22)( 68*8-1 downto  67*8), w69 => Pw(22)( 69*8-1 downto  68*8), w70 => Pw(22)( 70*8-1 downto  69*8), w71 => Pw(22)( 71*8-1 downto  70*8), w72 => Pw(22)( 72*8-1 downto  71*8), 
w73 => Pw(22)( 73*8-1 downto  72*8), w74 => Pw(22)( 74*8-1 downto  73*8), w75 => Pw(22)( 75*8-1 downto  74*8), w76 => Pw(22)( 76*8-1 downto  75*8), w77 => Pw(22)( 77*8-1 downto  76*8), w78 => Pw(22)( 78*8-1 downto  77*8), w79 => Pw(22)( 79*8-1 downto  78*8), w80 => Pw(22)( 80*8-1 downto  79*8), 
w81 => Pw(22)( 81*8-1 downto  80*8), w82 => Pw(22)( 82*8-1 downto  81*8), w83 => Pw(22)( 83*8-1 downto  82*8), w84 => Pw(22)( 84*8-1 downto  83*8), w85 => Pw(22)( 85*8-1 downto  84*8), w86 => Pw(22)( 86*8-1 downto  85*8), w87 => Pw(22)( 87*8-1 downto  86*8), w88 => Pw(22)( 88*8-1 downto  87*8), 
w89 => Pw(22)( 89*8-1 downto  88*8), w90 => Pw(22)( 90*8-1 downto  89*8), w91 => Pw(22)( 91*8-1 downto  90*8), w92 => Pw(22)( 92*8-1 downto  91*8), w93 => Pw(22)( 93*8-1 downto  92*8), w94 => Pw(22)( 94*8-1 downto  93*8), w95 => Pw(22)( 95*8-1 downto  94*8), w96 => Pw(22)( 96*8-1 downto  95*8), 
w97 => Pw(22)( 97*8-1 downto  96*8), w98 => Pw(22)( 98*8-1 downto  97*8), w99 => Pw(22)( 99*8-1 downto  98*8), w100=> Pw(22)(100*8-1 downto  99*8), w101=> Pw(22)(101*8-1 downto 100*8), w102=> Pw(22)(102*8-1 downto 101*8), w103=> Pw(22)(103*8-1 downto 102*8), w104=> Pw(22)(104*8-1 downto 103*8), 
w105=> Pw(22)(105*8-1 downto 104*8), w106=> Pw(22)(106*8-1 downto 105*8), w107=> Pw(22)(107*8-1 downto 106*8), w108=> Pw(22)(108*8-1 downto 107*8), w109=> Pw(22)(109*8-1 downto 108*8), w110=> Pw(22)(110*8-1 downto 109*8), w111=> Pw(22)(111*8-1 downto 110*8), w112=> Pw(22)(112*8-1 downto 111*8), 
w113=> Pw(22)(113*8-1 downto 112*8), w114=> Pw(22)(114*8-1 downto 113*8), w115=> Pw(22)(115*8-1 downto 114*8), w116=> Pw(22)(116*8-1 downto 115*8), w117=> Pw(22)(117*8-1 downto 116*8), w118=> Pw(22)(118*8-1 downto 117*8), w119=> Pw(22)(119*8-1 downto 118*8), w120=> Pw(22)(120*8-1 downto 119*8), 
w121=> Pw(22)(121*8-1 downto 120*8), w122=> Pw(22)(122*8-1 downto 121*8), w123=> Pw(22)(123*8-1 downto 122*8), w124=> Pw(22)(124*8-1 downto 123*8), w125=> Pw(22)(125*8-1 downto 124*8), w126=> Pw(22)(126*8-1 downto 125*8), w127=> Pw(22)(127*8-1 downto 126*8), w128=> Pw(22)(128*8-1 downto 127*8), 

           d_out   => pca_d22_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_23_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(23)(     7 downto    0), w02 => Pw(23)( 2*8-1 downto    8), w03 => Pw(23)( 3*8-1 downto  2*8), w04 => Pw(23)( 4*8-1 downto  3*8), w05 => Pw(23)( 5*8-1 downto  4*8), w06 => Pw(23)( 6*8-1 downto  5*8), w07 => Pw(23)( 7*8-1 downto  6*8), w08 => Pw(23)( 8*8-1 downto  7*8),  
w09 => Pw(23)( 9*8-1 downto  8*8), w10 => Pw(23)(10*8-1 downto  9*8), w11 => Pw(23)(11*8-1 downto 10*8), w12 => Pw(23)(12*8-1 downto 11*8), w13 => Pw(23)(13*8-1 downto 12*8), w14 => Pw(23)(14*8-1 downto 13*8), w15 => Pw(23)(15*8-1 downto 14*8), w16 => Pw(23)(16*8-1 downto 15*8),  
w17 => Pw(23)(17*8-1 downto 16*8), w18 => Pw(23)(18*8-1 downto 17*8), w19 => Pw(23)(19*8-1 downto 18*8), w20 => Pw(23)(20*8-1 downto 19*8), w21 => Pw(23)(21*8-1 downto 20*8), w22 => Pw(23)(22*8-1 downto 21*8), w23 => Pw(23)(23*8-1 downto 22*8), w24 => Pw(23)(24*8-1 downto 23*8),  
w25 => Pw(23)(25*8-1 downto 24*8), w26 => Pw(23)(26*8-1 downto 25*8), w27 => Pw(23)(27*8-1 downto 26*8), w28 => Pw(23)(28*8-1 downto 27*8), w29 => Pw(23)(29*8-1 downto 28*8), w30 => Pw(23)(30*8-1 downto 29*8), w31 => Pw(23)(31*8-1 downto 30*8), w32 => Pw(23)(32*8-1 downto 31*8),  
w33 => Pw(23)(33*8-1 downto 32*8), w34 => Pw(23)(34*8-1 downto 33*8), w35 => Pw(23)(35*8-1 downto 34*8), w36 => Pw(23)(36*8-1 downto 35*8), w37 => Pw(23)(37*8-1 downto 36*8), w38 => Pw(23)(38*8-1 downto 37*8), w39 => Pw(23)(39*8-1 downto 38*8), w40 => Pw(23)(40*8-1 downto 39*8),  
w41 => Pw(23)(41*8-1 downto 40*8), w42 => Pw(23)(42*8-1 downto 41*8), w43 => Pw(23)(43*8-1 downto 42*8), w44 => Pw(23)(44*8-1 downto 43*8), w45 => Pw(23)(45*8-1 downto 44*8), w46 => Pw(23)(46*8-1 downto 45*8), w47 => Pw(23)(47*8-1 downto 46*8), w48 => Pw(23)(48*8-1 downto 47*8),  
w49 => Pw(23)(49*8-1 downto 48*8), w50 => Pw(23)(50*8-1 downto 49*8), w51 => Pw(23)(51*8-1 downto 50*8), w52 => Pw(23)(52*8-1 downto 51*8), w53 => Pw(23)(53*8-1 downto 52*8), w54 => Pw(23)(54*8-1 downto 53*8), w55 => Pw(23)(55*8-1 downto 54*8), w56 => Pw(23)(56*8-1 downto 55*8),  
w57 => Pw(23)(57*8-1 downto 56*8), w58 => Pw(23)(58*8-1 downto 57*8), w59 => Pw(23)(59*8-1 downto 58*8), w60 => Pw(23)(60*8-1 downto 59*8), w61 => Pw(23)(61*8-1 downto 60*8), w62 => Pw(23)(62*8-1 downto 61*8), w63 => Pw(23)(63*8-1 downto 62*8), w64 => Pw(23)(64*8-1 downto 63*8), 
w65 => Pw(23)( 65*8-1 downto  64*8), w66 => Pw(23)( 66*8-1 downto  65*8), w67 => Pw(23)( 67*8-1 downto  66*8), w68 => Pw(23)( 68*8-1 downto  67*8), w69 => Pw(23)( 69*8-1 downto  68*8), w70 => Pw(23)( 70*8-1 downto  69*8), w71 => Pw(23)( 71*8-1 downto  70*8), w72 => Pw(23)( 72*8-1 downto  71*8), 
w73 => Pw(23)( 73*8-1 downto  72*8), w74 => Pw(23)( 74*8-1 downto  73*8), w75 => Pw(23)( 75*8-1 downto  74*8), w76 => Pw(23)( 76*8-1 downto  75*8), w77 => Pw(23)( 77*8-1 downto  76*8), w78 => Pw(23)( 78*8-1 downto  77*8), w79 => Pw(23)( 79*8-1 downto  78*8), w80 => Pw(23)( 80*8-1 downto  79*8), 
w81 => Pw(23)( 81*8-1 downto  80*8), w82 => Pw(23)( 82*8-1 downto  81*8), w83 => Pw(23)( 83*8-1 downto  82*8), w84 => Pw(23)( 84*8-1 downto  83*8), w85 => Pw(23)( 85*8-1 downto  84*8), w86 => Pw(23)( 86*8-1 downto  85*8), w87 => Pw(23)( 87*8-1 downto  86*8), w88 => Pw(23)( 88*8-1 downto  87*8), 
w89 => Pw(23)( 89*8-1 downto  88*8), w90 => Pw(23)( 90*8-1 downto  89*8), w91 => Pw(23)( 91*8-1 downto  90*8), w92 => Pw(23)( 92*8-1 downto  91*8), w93 => Pw(23)( 93*8-1 downto  92*8), w94 => Pw(23)( 94*8-1 downto  93*8), w95 => Pw(23)( 95*8-1 downto  94*8), w96 => Pw(23)( 96*8-1 downto  95*8), 
w97 => Pw(23)( 97*8-1 downto  96*8), w98 => Pw(23)( 98*8-1 downto  97*8), w99 => Pw(23)( 99*8-1 downto  98*8), w100=> Pw(23)(100*8-1 downto  99*8), w101=> Pw(23)(101*8-1 downto 100*8), w102=> Pw(23)(102*8-1 downto 101*8), w103=> Pw(23)(103*8-1 downto 102*8), w104=> Pw(23)(104*8-1 downto 103*8), 
w105=> Pw(23)(105*8-1 downto 104*8), w106=> Pw(23)(106*8-1 downto 105*8), w107=> Pw(23)(107*8-1 downto 106*8), w108=> Pw(23)(108*8-1 downto 107*8), w109=> Pw(23)(109*8-1 downto 108*8), w110=> Pw(23)(110*8-1 downto 109*8), w111=> Pw(23)(111*8-1 downto 110*8), w112=> Pw(23)(112*8-1 downto 111*8), 
w113=> Pw(23)(113*8-1 downto 112*8), w114=> Pw(23)(114*8-1 downto 113*8), w115=> Pw(23)(115*8-1 downto 114*8), w116=> Pw(23)(116*8-1 downto 115*8), w117=> Pw(23)(117*8-1 downto 116*8), w118=> Pw(23)(118*8-1 downto 117*8), w119=> Pw(23)(119*8-1 downto 118*8), w120=> Pw(23)(120*8-1 downto 119*8), 
w121=> Pw(23)(121*8-1 downto 120*8), w122=> Pw(23)(122*8-1 downto 121*8), w123=> Pw(23)(123*8-1 downto 122*8), w124=> Pw(23)(124*8-1 downto 123*8), w125=> Pw(23)(125*8-1 downto 124*8), w126=> Pw(23)(126*8-1 downto 125*8), w127=> Pw(23)(127*8-1 downto 126*8), w128=> Pw(23)(128*8-1 downto 127*8), 

           d_out   => pca_d23_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_24_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(24)(     7 downto    0), w02 => Pw(24)( 2*8-1 downto    8), w03 => Pw(24)( 3*8-1 downto  2*8), w04 => Pw(24)( 4*8-1 downto  3*8), w05 => Pw(24)( 5*8-1 downto  4*8), w06 => Pw(24)( 6*8-1 downto  5*8), w07 => Pw(24)( 7*8-1 downto  6*8), w08 => Pw(24)( 8*8-1 downto  7*8),  
w09 => Pw(24)( 9*8-1 downto  8*8), w10 => Pw(24)(10*8-1 downto  9*8), w11 => Pw(24)(11*8-1 downto 10*8), w12 => Pw(24)(12*8-1 downto 11*8), w13 => Pw(24)(13*8-1 downto 12*8), w14 => Pw(24)(14*8-1 downto 13*8), w15 => Pw(24)(15*8-1 downto 14*8), w16 => Pw(24)(16*8-1 downto 15*8),  
w17 => Pw(24)(17*8-1 downto 16*8), w18 => Pw(24)(18*8-1 downto 17*8), w19 => Pw(24)(19*8-1 downto 18*8), w20 => Pw(24)(20*8-1 downto 19*8), w21 => Pw(24)(21*8-1 downto 20*8), w22 => Pw(24)(22*8-1 downto 21*8), w23 => Pw(24)(23*8-1 downto 22*8), w24 => Pw(24)(24*8-1 downto 23*8),  
w25 => Pw(24)(25*8-1 downto 24*8), w26 => Pw(24)(26*8-1 downto 25*8), w27 => Pw(24)(27*8-1 downto 26*8), w28 => Pw(24)(28*8-1 downto 27*8), w29 => Pw(24)(29*8-1 downto 28*8), w30 => Pw(24)(30*8-1 downto 29*8), w31 => Pw(24)(31*8-1 downto 30*8), w32 => Pw(24)(32*8-1 downto 31*8),  
w33 => Pw(24)(33*8-1 downto 32*8), w34 => Pw(24)(34*8-1 downto 33*8), w35 => Pw(24)(35*8-1 downto 34*8), w36 => Pw(24)(36*8-1 downto 35*8), w37 => Pw(24)(37*8-1 downto 36*8), w38 => Pw(24)(38*8-1 downto 37*8), w39 => Pw(24)(39*8-1 downto 38*8), w40 => Pw(24)(40*8-1 downto 39*8),  
w41 => Pw(24)(41*8-1 downto 40*8), w42 => Pw(24)(42*8-1 downto 41*8), w43 => Pw(24)(43*8-1 downto 42*8), w44 => Pw(24)(44*8-1 downto 43*8), w45 => Pw(24)(45*8-1 downto 44*8), w46 => Pw(24)(46*8-1 downto 45*8), w47 => Pw(24)(47*8-1 downto 46*8), w48 => Pw(24)(48*8-1 downto 47*8),  
w49 => Pw(24)(49*8-1 downto 48*8), w50 => Pw(24)(50*8-1 downto 49*8), w51 => Pw(24)(51*8-1 downto 50*8), w52 => Pw(24)(52*8-1 downto 51*8), w53 => Pw(24)(53*8-1 downto 52*8), w54 => Pw(24)(54*8-1 downto 53*8), w55 => Pw(24)(55*8-1 downto 54*8), w56 => Pw(24)(56*8-1 downto 55*8),  
w57 => Pw(24)(57*8-1 downto 56*8), w58 => Pw(24)(58*8-1 downto 57*8), w59 => Pw(24)(59*8-1 downto 58*8), w60 => Pw(24)(60*8-1 downto 59*8), w61 => Pw(24)(61*8-1 downto 60*8), w62 => Pw(24)(62*8-1 downto 61*8), w63 => Pw(24)(63*8-1 downto 62*8), w64 => Pw(24)(64*8-1 downto 63*8), 
w65 => Pw(24)( 65*8-1 downto  64*8), w66 => Pw(24)( 66*8-1 downto  65*8), w67 => Pw(24)( 67*8-1 downto  66*8), w68 => Pw(24)( 68*8-1 downto  67*8), w69 => Pw(24)( 69*8-1 downto  68*8), w70 => Pw(24)( 70*8-1 downto  69*8), w71 => Pw(24)( 71*8-1 downto  70*8), w72 => Pw(24)( 72*8-1 downto  71*8), 
w73 => Pw(24)( 73*8-1 downto  72*8), w74 => Pw(24)( 74*8-1 downto  73*8), w75 => Pw(24)( 75*8-1 downto  74*8), w76 => Pw(24)( 76*8-1 downto  75*8), w77 => Pw(24)( 77*8-1 downto  76*8), w78 => Pw(24)( 78*8-1 downto  77*8), w79 => Pw(24)( 79*8-1 downto  78*8), w80 => Pw(24)( 80*8-1 downto  79*8), 
w81 => Pw(24)( 81*8-1 downto  80*8), w82 => Pw(24)( 82*8-1 downto  81*8), w83 => Pw(24)( 83*8-1 downto  82*8), w84 => Pw(24)( 84*8-1 downto  83*8), w85 => Pw(24)( 85*8-1 downto  84*8), w86 => Pw(24)( 86*8-1 downto  85*8), w87 => Pw(24)( 87*8-1 downto  86*8), w88 => Pw(24)( 88*8-1 downto  87*8), 
w89 => Pw(24)( 89*8-1 downto  88*8), w90 => Pw(24)( 90*8-1 downto  89*8), w91 => Pw(24)( 91*8-1 downto  90*8), w92 => Pw(24)( 92*8-1 downto  91*8), w93 => Pw(24)( 93*8-1 downto  92*8), w94 => Pw(24)( 94*8-1 downto  93*8), w95 => Pw(24)( 95*8-1 downto  94*8), w96 => Pw(24)( 96*8-1 downto  95*8), 
w97 => Pw(24)( 97*8-1 downto  96*8), w98 => Pw(24)( 98*8-1 downto  97*8), w99 => Pw(24)( 99*8-1 downto  98*8), w100=> Pw(24)(100*8-1 downto  99*8), w101=> Pw(24)(101*8-1 downto 100*8), w102=> Pw(24)(102*8-1 downto 101*8), w103=> Pw(24)(103*8-1 downto 102*8), w104=> Pw(24)(104*8-1 downto 103*8), 
w105=> Pw(24)(105*8-1 downto 104*8), w106=> Pw(24)(106*8-1 downto 105*8), w107=> Pw(24)(107*8-1 downto 106*8), w108=> Pw(24)(108*8-1 downto 107*8), w109=> Pw(24)(109*8-1 downto 108*8), w110=> Pw(24)(110*8-1 downto 109*8), w111=> Pw(24)(111*8-1 downto 110*8), w112=> Pw(24)(112*8-1 downto 111*8), 
w113=> Pw(24)(113*8-1 downto 112*8), w114=> Pw(24)(114*8-1 downto 113*8), w115=> Pw(24)(115*8-1 downto 114*8), w116=> Pw(24)(116*8-1 downto 115*8), w117=> Pw(24)(117*8-1 downto 116*8), w118=> Pw(24)(118*8-1 downto 117*8), w119=> Pw(24)(119*8-1 downto 118*8), w120=> Pw(24)(120*8-1 downto 119*8), 
w121=> Pw(24)(121*8-1 downto 120*8), w122=> Pw(24)(122*8-1 downto 121*8), w123=> Pw(24)(123*8-1 downto 122*8), w124=> Pw(24)(124*8-1 downto 123*8), w125=> Pw(24)(125*8-1 downto 124*8), w126=> Pw(24)(126*8-1 downto 125*8), w127=> Pw(24)(127*8-1 downto 126*8), w128=> Pw(24)(128*8-1 downto 127*8), 

           d_out   => pca_d24_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_25_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(25)(     7 downto    0), w02 => Pw(25)( 2*8-1 downto    8), w03 => Pw(25)( 3*8-1 downto  2*8), w04 => Pw(25)( 4*8-1 downto  3*8), w05 => Pw(25)( 5*8-1 downto  4*8), w06 => Pw(25)( 6*8-1 downto  5*8), w07 => Pw(25)( 7*8-1 downto  6*8), w08 => Pw(25)( 8*8-1 downto  7*8),  
w09 => Pw(25)( 9*8-1 downto  8*8), w10 => Pw(25)(10*8-1 downto  9*8), w11 => Pw(25)(11*8-1 downto 10*8), w12 => Pw(25)(12*8-1 downto 11*8), w13 => Pw(25)(13*8-1 downto 12*8), w14 => Pw(25)(14*8-1 downto 13*8), w15 => Pw(25)(15*8-1 downto 14*8), w16 => Pw(25)(16*8-1 downto 15*8),  
w17 => Pw(25)(17*8-1 downto 16*8), w18 => Pw(25)(18*8-1 downto 17*8), w19 => Pw(25)(19*8-1 downto 18*8), w20 => Pw(25)(20*8-1 downto 19*8), w21 => Pw(25)(21*8-1 downto 20*8), w22 => Pw(25)(22*8-1 downto 21*8), w23 => Pw(25)(23*8-1 downto 22*8), w24 => Pw(25)(24*8-1 downto 23*8),  
w25 => Pw(25)(25*8-1 downto 24*8), w26 => Pw(25)(26*8-1 downto 25*8), w27 => Pw(25)(27*8-1 downto 26*8), w28 => Pw(25)(28*8-1 downto 27*8), w29 => Pw(25)(29*8-1 downto 28*8), w30 => Pw(25)(30*8-1 downto 29*8), w31 => Pw(25)(31*8-1 downto 30*8), w32 => Pw(25)(32*8-1 downto 31*8),  
w33 => Pw(25)(33*8-1 downto 32*8), w34 => Pw(25)(34*8-1 downto 33*8), w35 => Pw(25)(35*8-1 downto 34*8), w36 => Pw(25)(36*8-1 downto 35*8), w37 => Pw(25)(37*8-1 downto 36*8), w38 => Pw(25)(38*8-1 downto 37*8), w39 => Pw(25)(39*8-1 downto 38*8), w40 => Pw(25)(40*8-1 downto 39*8),  
w41 => Pw(25)(41*8-1 downto 40*8), w42 => Pw(25)(42*8-1 downto 41*8), w43 => Pw(25)(43*8-1 downto 42*8), w44 => Pw(25)(44*8-1 downto 43*8), w45 => Pw(25)(45*8-1 downto 44*8), w46 => Pw(25)(46*8-1 downto 45*8), w47 => Pw(25)(47*8-1 downto 46*8), w48 => Pw(25)(48*8-1 downto 47*8),  
w49 => Pw(25)(49*8-1 downto 48*8), w50 => Pw(25)(50*8-1 downto 49*8), w51 => Pw(25)(51*8-1 downto 50*8), w52 => Pw(25)(52*8-1 downto 51*8), w53 => Pw(25)(53*8-1 downto 52*8), w54 => Pw(25)(54*8-1 downto 53*8), w55 => Pw(25)(55*8-1 downto 54*8), w56 => Pw(25)(56*8-1 downto 55*8),  
w57 => Pw(25)(57*8-1 downto 56*8), w58 => Pw(25)(58*8-1 downto 57*8), w59 => Pw(25)(59*8-1 downto 58*8), w60 => Pw(25)(60*8-1 downto 59*8), w61 => Pw(25)(61*8-1 downto 60*8), w62 => Pw(25)(62*8-1 downto 61*8), w63 => Pw(25)(63*8-1 downto 62*8), w64 => Pw(25)(64*8-1 downto 63*8), 
w65 => Pw(25)( 65*8-1 downto  64*8), w66 => Pw(25)( 66*8-1 downto  65*8), w67 => Pw(25)( 67*8-1 downto  66*8), w68 => Pw(25)( 68*8-1 downto  67*8), w69 => Pw(25)( 69*8-1 downto  68*8), w70 => Pw(25)( 70*8-1 downto  69*8), w71 => Pw(25)( 71*8-1 downto  70*8), w72 => Pw(25)( 72*8-1 downto  71*8), 
w73 => Pw(25)( 73*8-1 downto  72*8), w74 => Pw(25)( 74*8-1 downto  73*8), w75 => Pw(25)( 75*8-1 downto  74*8), w76 => Pw(25)( 76*8-1 downto  75*8), w77 => Pw(25)( 77*8-1 downto  76*8), w78 => Pw(25)( 78*8-1 downto  77*8), w79 => Pw(25)( 79*8-1 downto  78*8), w80 => Pw(25)( 80*8-1 downto  79*8), 
w81 => Pw(25)( 81*8-1 downto  80*8), w82 => Pw(25)( 82*8-1 downto  81*8), w83 => Pw(25)( 83*8-1 downto  82*8), w84 => Pw(25)( 84*8-1 downto  83*8), w85 => Pw(25)( 85*8-1 downto  84*8), w86 => Pw(25)( 86*8-1 downto  85*8), w87 => Pw(25)( 87*8-1 downto  86*8), w88 => Pw(25)( 88*8-1 downto  87*8), 
w89 => Pw(25)( 89*8-1 downto  88*8), w90 => Pw(25)( 90*8-1 downto  89*8), w91 => Pw(25)( 91*8-1 downto  90*8), w92 => Pw(25)( 92*8-1 downto  91*8), w93 => Pw(25)( 93*8-1 downto  92*8), w94 => Pw(25)( 94*8-1 downto  93*8), w95 => Pw(25)( 95*8-1 downto  94*8), w96 => Pw(25)( 96*8-1 downto  95*8), 
w97 => Pw(25)( 97*8-1 downto  96*8), w98 => Pw(25)( 98*8-1 downto  97*8), w99 => Pw(25)( 99*8-1 downto  98*8), w100=> Pw(25)(100*8-1 downto  99*8), w101=> Pw(25)(101*8-1 downto 100*8), w102=> Pw(25)(102*8-1 downto 101*8), w103=> Pw(25)(103*8-1 downto 102*8), w104=> Pw(25)(104*8-1 downto 103*8), 
w105=> Pw(25)(105*8-1 downto 104*8), w106=> Pw(25)(106*8-1 downto 105*8), w107=> Pw(25)(107*8-1 downto 106*8), w108=> Pw(25)(108*8-1 downto 107*8), w109=> Pw(25)(109*8-1 downto 108*8), w110=> Pw(25)(110*8-1 downto 109*8), w111=> Pw(25)(111*8-1 downto 110*8), w112=> Pw(25)(112*8-1 downto 111*8), 
w113=> Pw(25)(113*8-1 downto 112*8), w114=> Pw(25)(114*8-1 downto 113*8), w115=> Pw(25)(115*8-1 downto 114*8), w116=> Pw(25)(116*8-1 downto 115*8), w117=> Pw(25)(117*8-1 downto 116*8), w118=> Pw(25)(118*8-1 downto 117*8), w119=> Pw(25)(119*8-1 downto 118*8), w120=> Pw(25)(120*8-1 downto 119*8), 
w121=> Pw(25)(121*8-1 downto 120*8), w122=> Pw(25)(122*8-1 downto 121*8), w123=> Pw(25)(123*8-1 downto 122*8), w124=> Pw(25)(124*8-1 downto 123*8), w125=> Pw(25)(125*8-1 downto 124*8), w126=> Pw(25)(126*8-1 downto 125*8), w127=> Pw(25)(127*8-1 downto 126*8), w128=> Pw(25)(128*8-1 downto 127*8), 

           d_out   => pca_d25_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_26_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 

d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(26)(     7 downto    0), w02 => Pw(26)( 2*8-1 downto    8), w03 => Pw(26)( 3*8-1 downto  2*8), w04 => Pw(26)( 4*8-1 downto  3*8), w05 => Pw(26)( 5*8-1 downto  4*8), w06 => Pw(26)( 6*8-1 downto  5*8), w07 => Pw(26)( 7*8-1 downto  6*8), w08 => Pw(26)( 8*8-1 downto  7*8),  
w09 => Pw(26)( 9*8-1 downto  8*8), w10 => Pw(26)(10*8-1 downto  9*8), w11 => Pw(26)(11*8-1 downto 10*8), w12 => Pw(26)(12*8-1 downto 11*8), w13 => Pw(26)(13*8-1 downto 12*8), w14 => Pw(26)(14*8-1 downto 13*8), w15 => Pw(26)(15*8-1 downto 14*8), w16 => Pw(26)(16*8-1 downto 15*8),  
w17 => Pw(26)(17*8-1 downto 16*8), w18 => Pw(26)(18*8-1 downto 17*8), w19 => Pw(26)(19*8-1 downto 18*8), w20 => Pw(26)(20*8-1 downto 19*8), w21 => Pw(26)(21*8-1 downto 20*8), w22 => Pw(26)(22*8-1 downto 21*8), w23 => Pw(26)(23*8-1 downto 22*8), w24 => Pw(26)(24*8-1 downto 23*8),  
w25 => Pw(26)(25*8-1 downto 24*8), w26 => Pw(26)(26*8-1 downto 25*8), w27 => Pw(26)(27*8-1 downto 26*8), w28 => Pw(26)(28*8-1 downto 27*8), w29 => Pw(26)(29*8-1 downto 28*8), w30 => Pw(26)(30*8-1 downto 29*8), w31 => Pw(26)(31*8-1 downto 30*8), w32 => Pw(26)(32*8-1 downto 31*8),  
w33 => Pw(26)(33*8-1 downto 32*8), w34 => Pw(26)(34*8-1 downto 33*8), w35 => Pw(26)(35*8-1 downto 34*8), w36 => Pw(26)(36*8-1 downto 35*8), w37 => Pw(26)(37*8-1 downto 36*8), w38 => Pw(26)(38*8-1 downto 37*8), w39 => Pw(26)(39*8-1 downto 38*8), w40 => Pw(26)(40*8-1 downto 39*8),  
w41 => Pw(26)(41*8-1 downto 40*8), w42 => Pw(26)(42*8-1 downto 41*8), w43 => Pw(26)(43*8-1 downto 42*8), w44 => Pw(26)(44*8-1 downto 43*8), w45 => Pw(26)(45*8-1 downto 44*8), w46 => Pw(26)(46*8-1 downto 45*8), w47 => Pw(26)(47*8-1 downto 46*8), w48 => Pw(26)(48*8-1 downto 47*8),  
w49 => Pw(26)(49*8-1 downto 48*8), w50 => Pw(26)(50*8-1 downto 49*8), w51 => Pw(26)(51*8-1 downto 50*8), w52 => Pw(26)(52*8-1 downto 51*8), w53 => Pw(26)(53*8-1 downto 52*8), w54 => Pw(26)(54*8-1 downto 53*8), w55 => Pw(26)(55*8-1 downto 54*8), w56 => Pw(26)(56*8-1 downto 55*8),  
w57 => Pw(26)(57*8-1 downto 56*8), w58 => Pw(26)(58*8-1 downto 57*8), w59 => Pw(26)(59*8-1 downto 58*8), w60 => Pw(26)(60*8-1 downto 59*8), w61 => Pw(26)(61*8-1 downto 60*8), w62 => Pw(26)(62*8-1 downto 61*8), w63 => Pw(26)(63*8-1 downto 62*8), w64 => Pw(26)(64*8-1 downto 63*8), 
w65 => Pw(26)( 65*8-1 downto  64*8), w66 => Pw(26)( 66*8-1 downto  65*8), w67 => Pw(26)( 67*8-1 downto  66*8), w68 => Pw(26)( 68*8-1 downto  67*8), w69 => Pw(26)( 69*8-1 downto  68*8), w70 => Pw(26)( 70*8-1 downto  69*8), w71 => Pw(26)( 71*8-1 downto  70*8), w72 => Pw(26)( 72*8-1 downto  71*8), 
w73 => Pw(26)( 73*8-1 downto  72*8), w74 => Pw(26)( 74*8-1 downto  73*8), w75 => Pw(26)( 75*8-1 downto  74*8), w76 => Pw(26)( 76*8-1 downto  75*8), w77 => Pw(26)( 77*8-1 downto  76*8), w78 => Pw(26)( 78*8-1 downto  77*8), w79 => Pw(26)( 79*8-1 downto  78*8), w80 => Pw(26)( 80*8-1 downto  79*8), 
w81 => Pw(26)( 81*8-1 downto  80*8), w82 => Pw(26)( 82*8-1 downto  81*8), w83 => Pw(26)( 83*8-1 downto  82*8), w84 => Pw(26)( 84*8-1 downto  83*8), w85 => Pw(26)( 85*8-1 downto  84*8), w86 => Pw(26)( 86*8-1 downto  85*8), w87 => Pw(26)( 87*8-1 downto  86*8), w88 => Pw(26)( 88*8-1 downto  87*8), 
w89 => Pw(26)( 89*8-1 downto  88*8), w90 => Pw(26)( 90*8-1 downto  89*8), w91 => Pw(26)( 91*8-1 downto  90*8), w92 => Pw(26)( 92*8-1 downto  91*8), w93 => Pw(26)( 93*8-1 downto  92*8), w94 => Pw(26)( 94*8-1 downto  93*8), w95 => Pw(26)( 95*8-1 downto  94*8), w96 => Pw(26)( 96*8-1 downto  95*8), 
w97 => Pw(26)( 97*8-1 downto  96*8), w98 => Pw(26)( 98*8-1 downto  97*8), w99 => Pw(26)( 99*8-1 downto  98*8), w100=> Pw(26)(100*8-1 downto  99*8), w101=> Pw(26)(101*8-1 downto 100*8), w102=> Pw(26)(102*8-1 downto 101*8), w103=> Pw(26)(103*8-1 downto 102*8), w104=> Pw(26)(104*8-1 downto 103*8), 
w105=> Pw(26)(105*8-1 downto 104*8), w106=> Pw(26)(106*8-1 downto 105*8), w107=> Pw(26)(107*8-1 downto 106*8), w108=> Pw(26)(108*8-1 downto 107*8), w109=> Pw(26)(109*8-1 downto 108*8), w110=> Pw(26)(110*8-1 downto 109*8), w111=> Pw(26)(111*8-1 downto 110*8), w112=> Pw(26)(112*8-1 downto 111*8), 
w113=> Pw(26)(113*8-1 downto 112*8), w114=> Pw(26)(114*8-1 downto 113*8), w115=> Pw(26)(115*8-1 downto 114*8), w116=> Pw(26)(116*8-1 downto 115*8), w117=> Pw(26)(117*8-1 downto 116*8), w118=> Pw(26)(118*8-1 downto 117*8), w119=> Pw(26)(119*8-1 downto 118*8), w120=> Pw(26)(120*8-1 downto 119*8), 
w121=> Pw(26)(121*8-1 downto 120*8), w122=> Pw(26)(122*8-1 downto 121*8), w123=> Pw(26)(123*8-1 downto 122*8), w124=> Pw(26)(124*8-1 downto 123*8), w125=> Pw(26)(125*8-1 downto 124*8), w126=> Pw(26)(126*8-1 downto 125*8), w127=> Pw(26)(127*8-1 downto 126*8), w128=> Pw(26)(128*8-1 downto 127*8), 

           d_out   => pca_d26_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_27_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 

d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(27)(     7 downto    0), w02 => Pw(27)( 2*8-1 downto    8), w03 => Pw(27)( 3*8-1 downto  2*8), w04 => Pw(27)( 4*8-1 downto  3*8), w05 => Pw(27)( 5*8-1 downto  4*8), w06 => Pw(27)( 6*8-1 downto  5*8), w07 => Pw(27)( 7*8-1 downto  6*8), w08 => Pw(27)( 8*8-1 downto  7*8),  
w09 => Pw(27)( 9*8-1 downto  8*8), w10 => Pw(27)(10*8-1 downto  9*8), w11 => Pw(27)(11*8-1 downto 10*8), w12 => Pw(27)(12*8-1 downto 11*8), w13 => Pw(27)(13*8-1 downto 12*8), w14 => Pw(27)(14*8-1 downto 13*8), w15 => Pw(27)(15*8-1 downto 14*8), w16 => Pw(27)(16*8-1 downto 15*8),  
w17 => Pw(27)(17*8-1 downto 16*8), w18 => Pw(27)(18*8-1 downto 17*8), w19 => Pw(27)(19*8-1 downto 18*8), w20 => Pw(27)(20*8-1 downto 19*8), w21 => Pw(27)(21*8-1 downto 20*8), w22 => Pw(27)(22*8-1 downto 21*8), w23 => Pw(27)(23*8-1 downto 22*8), w24 => Pw(27)(24*8-1 downto 23*8),  
w25 => Pw(27)(25*8-1 downto 24*8), w26 => Pw(27)(26*8-1 downto 25*8), w27 => Pw(27)(27*8-1 downto 26*8), w28 => Pw(27)(28*8-1 downto 27*8), w29 => Pw(27)(29*8-1 downto 28*8), w30 => Pw(27)(30*8-1 downto 29*8), w31 => Pw(27)(31*8-1 downto 30*8), w32 => Pw(27)(32*8-1 downto 31*8),  
w33 => Pw(27)(33*8-1 downto 32*8), w34 => Pw(27)(34*8-1 downto 33*8), w35 => Pw(27)(35*8-1 downto 34*8), w36 => Pw(27)(36*8-1 downto 35*8), w37 => Pw(27)(37*8-1 downto 36*8), w38 => Pw(27)(38*8-1 downto 37*8), w39 => Pw(27)(39*8-1 downto 38*8), w40 => Pw(27)(40*8-1 downto 39*8),  
w41 => Pw(27)(41*8-1 downto 40*8), w42 => Pw(27)(42*8-1 downto 41*8), w43 => Pw(27)(43*8-1 downto 42*8), w44 => Pw(27)(44*8-1 downto 43*8), w45 => Pw(27)(45*8-1 downto 44*8), w46 => Pw(27)(46*8-1 downto 45*8), w47 => Pw(27)(47*8-1 downto 46*8), w48 => Pw(27)(48*8-1 downto 47*8),  
w49 => Pw(27)(49*8-1 downto 48*8), w50 => Pw(27)(50*8-1 downto 49*8), w51 => Pw(27)(51*8-1 downto 50*8), w52 => Pw(27)(52*8-1 downto 51*8), w53 => Pw(27)(53*8-1 downto 52*8), w54 => Pw(27)(54*8-1 downto 53*8), w55 => Pw(27)(55*8-1 downto 54*8), w56 => Pw(27)(56*8-1 downto 55*8),  
w57 => Pw(27)(57*8-1 downto 56*8), w58 => Pw(27)(58*8-1 downto 57*8), w59 => Pw(27)(59*8-1 downto 58*8), w60 => Pw(27)(60*8-1 downto 59*8), w61 => Pw(27)(61*8-1 downto 60*8), w62 => Pw(27)(62*8-1 downto 61*8), w63 => Pw(27)(63*8-1 downto 62*8), w64 => Pw(27)(64*8-1 downto 63*8), 
w65 => Pw(27)( 65*8-1 downto  64*8), w66 => Pw(27)( 66*8-1 downto  65*8), w67 => Pw(27)( 67*8-1 downto  66*8), w68 => Pw(27)( 68*8-1 downto  67*8), w69 => Pw(27)( 69*8-1 downto  68*8), w70 => Pw(27)( 70*8-1 downto  69*8), w71 => Pw(27)( 71*8-1 downto  70*8), w72 => Pw(27)( 72*8-1 downto  71*8), 
w73 => Pw(27)( 73*8-1 downto  72*8), w74 => Pw(27)( 74*8-1 downto  73*8), w75 => Pw(27)( 75*8-1 downto  74*8), w76 => Pw(27)( 76*8-1 downto  75*8), w77 => Pw(27)( 77*8-1 downto  76*8), w78 => Pw(27)( 78*8-1 downto  77*8), w79 => Pw(27)( 79*8-1 downto  78*8), w80 => Pw(27)( 80*8-1 downto  79*8), 
w81 => Pw(27)( 81*8-1 downto  80*8), w82 => Pw(27)( 82*8-1 downto  81*8), w83 => Pw(27)( 83*8-1 downto  82*8), w84 => Pw(27)( 84*8-1 downto  83*8), w85 => Pw(27)( 85*8-1 downto  84*8), w86 => Pw(27)( 86*8-1 downto  85*8), w87 => Pw(27)( 87*8-1 downto  86*8), w88 => Pw(27)( 88*8-1 downto  87*8), 
w89 => Pw(27)( 89*8-1 downto  88*8), w90 => Pw(27)( 90*8-1 downto  89*8), w91 => Pw(27)( 91*8-1 downto  90*8), w92 => Pw(27)( 92*8-1 downto  91*8), w93 => Pw(27)( 93*8-1 downto  92*8), w94 => Pw(27)( 94*8-1 downto  93*8), w95 => Pw(27)( 95*8-1 downto  94*8), w96 => Pw(27)( 96*8-1 downto  95*8), 
w97 => Pw(27)( 97*8-1 downto  96*8), w98 => Pw(27)( 98*8-1 downto  97*8), w99 => Pw(27)( 99*8-1 downto  98*8), w100=> Pw(27)(100*8-1 downto  99*8), w101=> Pw(27)(101*8-1 downto 100*8), w102=> Pw(27)(102*8-1 downto 101*8), w103=> Pw(27)(103*8-1 downto 102*8), w104=> Pw(27)(104*8-1 downto 103*8), 
w105=> Pw(27)(105*8-1 downto 104*8), w106=> Pw(27)(106*8-1 downto 105*8), w107=> Pw(27)(107*8-1 downto 106*8), w108=> Pw(27)(108*8-1 downto 107*8), w109=> Pw(27)(109*8-1 downto 108*8), w110=> Pw(27)(110*8-1 downto 109*8), w111=> Pw(27)(111*8-1 downto 110*8), w112=> Pw(27)(112*8-1 downto 111*8), 
w113=> Pw(27)(113*8-1 downto 112*8), w114=> Pw(27)(114*8-1 downto 113*8), w115=> Pw(27)(115*8-1 downto 114*8), w116=> Pw(27)(116*8-1 downto 115*8), w117=> Pw(27)(117*8-1 downto 116*8), w118=> Pw(27)(118*8-1 downto 117*8), w119=> Pw(27)(119*8-1 downto 118*8), w120=> Pw(27)(120*8-1 downto 119*8), 
w121=> Pw(27)(121*8-1 downto 120*8), w122=> Pw(27)(122*8-1 downto 121*8), w123=> Pw(27)(123*8-1 downto 122*8), w124=> Pw(27)(124*8-1 downto 123*8), w125=> Pw(27)(125*8-1 downto 124*8), w126=> Pw(27)(126*8-1 downto 125*8), w127=> Pw(27)(127*8-1 downto 126*8), w128=> Pw(27)(128*8-1 downto 127*8), 

           d_out   => pca_d27_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_28_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(28)(     7 downto    0), w02 => Pw(28)( 2*8-1 downto    8), w03 => Pw(28)( 3*8-1 downto  2*8), w04 => Pw(28)( 4*8-1 downto  3*8), w05 => Pw(28)( 5*8-1 downto  4*8), w06 => Pw(28)( 6*8-1 downto  5*8), w07 => Pw(28)( 7*8-1 downto  6*8), w08 => Pw(28)( 8*8-1 downto  7*8),  
w09 => Pw(28)( 9*8-1 downto  8*8), w10 => Pw(28)(10*8-1 downto  9*8), w11 => Pw(28)(11*8-1 downto 10*8), w12 => Pw(28)(12*8-1 downto 11*8), w13 => Pw(28)(13*8-1 downto 12*8), w14 => Pw(28)(14*8-1 downto 13*8), w15 => Pw(28)(15*8-1 downto 14*8), w16 => Pw(28)(16*8-1 downto 15*8),  
w17 => Pw(28)(17*8-1 downto 16*8), w18 => Pw(28)(18*8-1 downto 17*8), w19 => Pw(28)(19*8-1 downto 18*8), w20 => Pw(28)(20*8-1 downto 19*8), w21 => Pw(28)(21*8-1 downto 20*8), w22 => Pw(28)(22*8-1 downto 21*8), w23 => Pw(28)(23*8-1 downto 22*8), w24 => Pw(28)(24*8-1 downto 23*8),  
w25 => Pw(28)(25*8-1 downto 24*8), w26 => Pw(28)(26*8-1 downto 25*8), w27 => Pw(28)(27*8-1 downto 26*8), w28 => Pw(28)(28*8-1 downto 27*8), w29 => Pw(28)(29*8-1 downto 28*8), w30 => Pw(28)(30*8-1 downto 29*8), w31 => Pw(28)(31*8-1 downto 30*8), w32 => Pw(28)(32*8-1 downto 31*8),  
w33 => Pw(28)(33*8-1 downto 32*8), w34 => Pw(28)(34*8-1 downto 33*8), w35 => Pw(28)(35*8-1 downto 34*8), w36 => Pw(28)(36*8-1 downto 35*8), w37 => Pw(28)(37*8-1 downto 36*8), w38 => Pw(28)(38*8-1 downto 37*8), w39 => Pw(28)(39*8-1 downto 38*8), w40 => Pw(28)(40*8-1 downto 39*8),  
w41 => Pw(28)(41*8-1 downto 40*8), w42 => Pw(28)(42*8-1 downto 41*8), w43 => Pw(28)(43*8-1 downto 42*8), w44 => Pw(28)(44*8-1 downto 43*8), w45 => Pw(28)(45*8-1 downto 44*8), w46 => Pw(28)(46*8-1 downto 45*8), w47 => Pw(28)(47*8-1 downto 46*8), w48 => Pw(28)(48*8-1 downto 47*8),  
w49 => Pw(28)(49*8-1 downto 48*8), w50 => Pw(28)(50*8-1 downto 49*8), w51 => Pw(28)(51*8-1 downto 50*8), w52 => Pw(28)(52*8-1 downto 51*8), w53 => Pw(28)(53*8-1 downto 52*8), w54 => Pw(28)(54*8-1 downto 53*8), w55 => Pw(28)(55*8-1 downto 54*8), w56 => Pw(28)(56*8-1 downto 55*8),  
w57 => Pw(28)(57*8-1 downto 56*8), w58 => Pw(28)(58*8-1 downto 57*8), w59 => Pw(28)(59*8-1 downto 58*8), w60 => Pw(28)(60*8-1 downto 59*8), w61 => Pw(28)(61*8-1 downto 60*8), w62 => Pw(28)(62*8-1 downto 61*8), w63 => Pw(28)(63*8-1 downto 62*8), w64 => Pw(28)(64*8-1 downto 63*8), 
w65 => Pw(28)( 65*8-1 downto  64*8), w66 => Pw(28)( 66*8-1 downto  65*8), w67 => Pw(28)( 67*8-1 downto  66*8), w68 => Pw(28)( 68*8-1 downto  67*8), w69 => Pw(28)( 69*8-1 downto  68*8), w70 => Pw(28)( 70*8-1 downto  69*8), w71 => Pw(28)( 71*8-1 downto  70*8), w72 => Pw(28)( 72*8-1 downto  71*8), 
w73 => Pw(28)( 73*8-1 downto  72*8), w74 => Pw(28)( 74*8-1 downto  73*8), w75 => Pw(28)( 75*8-1 downto  74*8), w76 => Pw(28)( 76*8-1 downto  75*8), w77 => Pw(28)( 77*8-1 downto  76*8), w78 => Pw(28)( 78*8-1 downto  77*8), w79 => Pw(28)( 79*8-1 downto  78*8), w80 => Pw(28)( 80*8-1 downto  79*8), 
w81 => Pw(28)( 81*8-1 downto  80*8), w82 => Pw(28)( 82*8-1 downto  81*8), w83 => Pw(28)( 83*8-1 downto  82*8), w84 => Pw(28)( 84*8-1 downto  83*8), w85 => Pw(28)( 85*8-1 downto  84*8), w86 => Pw(28)( 86*8-1 downto  85*8), w87 => Pw(28)( 87*8-1 downto  86*8), w88 => Pw(28)( 88*8-1 downto  87*8), 
w89 => Pw(28)( 89*8-1 downto  88*8), w90 => Pw(28)( 90*8-1 downto  89*8), w91 => Pw(28)( 91*8-1 downto  90*8), w92 => Pw(28)( 92*8-1 downto  91*8), w93 => Pw(28)( 93*8-1 downto  92*8), w94 => Pw(28)( 94*8-1 downto  93*8), w95 => Pw(28)( 95*8-1 downto  94*8), w96 => Pw(28)( 96*8-1 downto  95*8), 
w97 => Pw(28)( 97*8-1 downto  96*8), w98 => Pw(28)( 98*8-1 downto  97*8), w99 => Pw(28)( 99*8-1 downto  98*8), w100=> Pw(28)(100*8-1 downto  99*8), w101=> Pw(28)(101*8-1 downto 100*8), w102=> Pw(28)(102*8-1 downto 101*8), w103=> Pw(28)(103*8-1 downto 102*8), w104=> Pw(28)(104*8-1 downto 103*8), 
w105=> Pw(28)(105*8-1 downto 104*8), w106=> Pw(28)(106*8-1 downto 105*8), w107=> Pw(28)(107*8-1 downto 106*8), w108=> Pw(28)(108*8-1 downto 107*8), w109=> Pw(28)(109*8-1 downto 108*8), w110=> Pw(28)(110*8-1 downto 109*8), w111=> Pw(28)(111*8-1 downto 110*8), w112=> Pw(28)(112*8-1 downto 111*8), 
w113=> Pw(28)(113*8-1 downto 112*8), w114=> Pw(28)(114*8-1 downto 113*8), w115=> Pw(28)(115*8-1 downto 114*8), w116=> Pw(28)(116*8-1 downto 115*8), w117=> Pw(28)(117*8-1 downto 116*8), w118=> Pw(28)(118*8-1 downto 117*8), w119=> Pw(28)(119*8-1 downto 118*8), w120=> Pw(28)(120*8-1 downto 119*8), 
w121=> Pw(28)(121*8-1 downto 120*8), w122=> Pw(28)(122*8-1 downto 121*8), w123=> Pw(28)(123*8-1 downto 122*8), w124=> Pw(28)(124*8-1 downto 123*8), w125=> Pw(28)(125*8-1 downto 124*8), w126=> Pw(28)(126*8-1 downto 125*8), w127=> Pw(28)(127*8-1 downto 126*8), w128=> Pw(28)(128*8-1 downto 127*8), 

           d_out   => pca_d28_out   ,
           en_out  => open  ,
           sof_out => open );

  
  PCA128_29_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(29)(     7 downto    0), w02 => Pw(29)( 2*8-1 downto    8), w03 => Pw(29)( 3*8-1 downto  2*8), w04 => Pw(29)( 4*8-1 downto  3*8), w05 => Pw(29)( 5*8-1 downto  4*8), w06 => Pw(29)( 6*8-1 downto  5*8), w07 => Pw(29)( 7*8-1 downto  6*8), w08 => Pw(29)( 8*8-1 downto  7*8),  
w09 => Pw(29)( 9*8-1 downto  8*8), w10 => Pw(29)(10*8-1 downto  9*8), w11 => Pw(29)(11*8-1 downto 10*8), w12 => Pw(29)(12*8-1 downto 11*8), w13 => Pw(29)(13*8-1 downto 12*8), w14 => Pw(29)(14*8-1 downto 13*8), w15 => Pw(29)(15*8-1 downto 14*8), w16 => Pw(29)(16*8-1 downto 15*8),  
w17 => Pw(29)(17*8-1 downto 16*8), w18 => Pw(29)(18*8-1 downto 17*8), w19 => Pw(29)(19*8-1 downto 18*8), w20 => Pw(29)(20*8-1 downto 19*8), w21 => Pw(29)(21*8-1 downto 20*8), w22 => Pw(29)(22*8-1 downto 21*8), w23 => Pw(29)(23*8-1 downto 22*8), w24 => Pw(29)(24*8-1 downto 23*8),  
w25 => Pw(29)(25*8-1 downto 24*8), w26 => Pw(29)(26*8-1 downto 25*8), w27 => Pw(29)(27*8-1 downto 26*8), w28 => Pw(29)(28*8-1 downto 27*8), w29 => Pw(29)(29*8-1 downto 28*8), w30 => Pw(29)(30*8-1 downto 29*8), w31 => Pw(29)(31*8-1 downto 30*8), w32 => Pw(29)(32*8-1 downto 31*8),  
w33 => Pw(29)(33*8-1 downto 32*8), w34 => Pw(29)(34*8-1 downto 33*8), w35 => Pw(29)(35*8-1 downto 34*8), w36 => Pw(29)(36*8-1 downto 35*8), w37 => Pw(29)(37*8-1 downto 36*8), w38 => Pw(29)(38*8-1 downto 37*8), w39 => Pw(29)(39*8-1 downto 38*8), w40 => Pw(29)(40*8-1 downto 39*8),  
w41 => Pw(29)(41*8-1 downto 40*8), w42 => Pw(29)(42*8-1 downto 41*8), w43 => Pw(29)(43*8-1 downto 42*8), w44 => Pw(29)(44*8-1 downto 43*8), w45 => Pw(29)(45*8-1 downto 44*8), w46 => Pw(29)(46*8-1 downto 45*8), w47 => Pw(29)(47*8-1 downto 46*8), w48 => Pw(29)(48*8-1 downto 47*8),  
w49 => Pw(29)(49*8-1 downto 48*8), w50 => Pw(29)(50*8-1 downto 49*8), w51 => Pw(29)(51*8-1 downto 50*8), w52 => Pw(29)(52*8-1 downto 51*8), w53 => Pw(29)(53*8-1 downto 52*8), w54 => Pw(29)(54*8-1 downto 53*8), w55 => Pw(29)(55*8-1 downto 54*8), w56 => Pw(29)(56*8-1 downto 55*8),  
w57 => Pw(29)(57*8-1 downto 56*8), w58 => Pw(29)(58*8-1 downto 57*8), w59 => Pw(29)(59*8-1 downto 58*8), w60 => Pw(29)(60*8-1 downto 59*8), w61 => Pw(29)(61*8-1 downto 60*8), w62 => Pw(29)(62*8-1 downto 61*8), w63 => Pw(29)(63*8-1 downto 62*8), w64 => Pw(29)(64*8-1 downto 63*8), 
w65 => Pw(29)( 65*8-1 downto  64*8), w66 => Pw(29)( 66*8-1 downto  65*8), w67 => Pw(29)( 67*8-1 downto  66*8), w68 => Pw(29)( 68*8-1 downto  67*8), w69 => Pw(29)( 69*8-1 downto  68*8), w70 => Pw(29)( 70*8-1 downto  69*8), w71 => Pw(29)( 71*8-1 downto  70*8), w72 => Pw(29)( 72*8-1 downto  71*8), 
w73 => Pw(29)( 73*8-1 downto  72*8), w74 => Pw(29)( 74*8-1 downto  73*8), w75 => Pw(29)( 75*8-1 downto  74*8), w76 => Pw(29)( 76*8-1 downto  75*8), w77 => Pw(29)( 77*8-1 downto  76*8), w78 => Pw(29)( 78*8-1 downto  77*8), w79 => Pw(29)( 79*8-1 downto  78*8), w80 => Pw(29)( 80*8-1 downto  79*8), 
w81 => Pw(29)( 81*8-1 downto  80*8), w82 => Pw(29)( 82*8-1 downto  81*8), w83 => Pw(29)( 83*8-1 downto  82*8), w84 => Pw(29)( 84*8-1 downto  83*8), w85 => Pw(29)( 85*8-1 downto  84*8), w86 => Pw(29)( 86*8-1 downto  85*8), w87 => Pw(29)( 87*8-1 downto  86*8), w88 => Pw(29)( 88*8-1 downto  87*8), 
w89 => Pw(29)( 89*8-1 downto  88*8), w90 => Pw(29)( 90*8-1 downto  89*8), w91 => Pw(29)( 91*8-1 downto  90*8), w92 => Pw(29)( 92*8-1 downto  91*8), w93 => Pw(29)( 93*8-1 downto  92*8), w94 => Pw(29)( 94*8-1 downto  93*8), w95 => Pw(29)( 95*8-1 downto  94*8), w96 => Pw(29)( 96*8-1 downto  95*8), 
w97 => Pw(29)( 97*8-1 downto  96*8), w98 => Pw(29)( 98*8-1 downto  97*8), w99 => Pw(29)( 99*8-1 downto  98*8), w100=> Pw(29)(100*8-1 downto  99*8), w101=> Pw(29)(101*8-1 downto 100*8), w102=> Pw(29)(102*8-1 downto 101*8), w103=> Pw(29)(103*8-1 downto 102*8), w104=> Pw(29)(104*8-1 downto 103*8), 
w105=> Pw(29)(105*8-1 downto 104*8), w106=> Pw(29)(106*8-1 downto 105*8), w107=> Pw(29)(107*8-1 downto 106*8), w108=> Pw(29)(108*8-1 downto 107*8), w109=> Pw(29)(109*8-1 downto 108*8), w110=> Pw(29)(110*8-1 downto 109*8), w111=> Pw(29)(111*8-1 downto 110*8), w112=> Pw(29)(112*8-1 downto 111*8), 
w113=> Pw(29)(113*8-1 downto 112*8), w114=> Pw(29)(114*8-1 downto 113*8), w115=> Pw(29)(115*8-1 downto 114*8), w116=> Pw(29)(116*8-1 downto 115*8), w117=> Pw(29)(117*8-1 downto 116*8), w118=> Pw(29)(118*8-1 downto 117*8), w119=> Pw(29)(119*8-1 downto 118*8), w120=> Pw(29)(120*8-1 downto 119*8), 
w121=> Pw(29)(121*8-1 downto 120*8), w122=> Pw(29)(122*8-1 downto 121*8), w123=> Pw(29)(123*8-1 downto 122*8), w124=> Pw(29)(124*8-1 downto 123*8), w125=> Pw(29)(125*8-1 downto 124*8), w126=> Pw(29)(126*8-1 downto 125*8), w127=> Pw(29)(127*8-1 downto 126*8), w128=> Pw(29)(128*8-1 downto 127*8), 

           d_out   => pca_d29_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_30_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(30)(     7 downto    0), w02 => Pw(30)( 2*8-1 downto    8), w03 => Pw(30)( 3*8-1 downto  2*8), w04 => Pw(30)( 4*8-1 downto  3*8), w05 => Pw(30)( 5*8-1 downto  4*8), w06 => Pw(30)( 6*8-1 downto  5*8), w07 => Pw(30)( 7*8-1 downto  6*8), w08 => Pw(30)( 8*8-1 downto  7*8),  
w09 => Pw(30)( 9*8-1 downto  8*8), w10 => Pw(30)(10*8-1 downto  9*8), w11 => Pw(30)(11*8-1 downto 10*8), w12 => Pw(30)(12*8-1 downto 11*8), w13 => Pw(30)(13*8-1 downto 12*8), w14 => Pw(30)(14*8-1 downto 13*8), w15 => Pw(30)(15*8-1 downto 14*8), w16 => Pw(30)(16*8-1 downto 15*8),  
w17 => Pw(30)(17*8-1 downto 16*8), w18 => Pw(30)(18*8-1 downto 17*8), w19 => Pw(30)(19*8-1 downto 18*8), w20 => Pw(30)(20*8-1 downto 19*8), w21 => Pw(30)(21*8-1 downto 20*8), w22 => Pw(30)(22*8-1 downto 21*8), w23 => Pw(30)(23*8-1 downto 22*8), w24 => Pw(30)(24*8-1 downto 23*8),  
w25 => Pw(30)(25*8-1 downto 24*8), w26 => Pw(30)(26*8-1 downto 25*8), w27 => Pw(30)(27*8-1 downto 26*8), w28 => Pw(30)(28*8-1 downto 27*8), w29 => Pw(30)(29*8-1 downto 28*8), w30 => Pw(30)(30*8-1 downto 29*8), w31 => Pw(30)(31*8-1 downto 30*8), w32 => Pw(30)(32*8-1 downto 31*8),  
w33 => Pw(30)(33*8-1 downto 32*8), w34 => Pw(30)(34*8-1 downto 33*8), w35 => Pw(30)(35*8-1 downto 34*8), w36 => Pw(30)(36*8-1 downto 35*8), w37 => Pw(30)(37*8-1 downto 36*8), w38 => Pw(30)(38*8-1 downto 37*8), w39 => Pw(30)(39*8-1 downto 38*8), w40 => Pw(30)(40*8-1 downto 39*8),  
w41 => Pw(30)(41*8-1 downto 40*8), w42 => Pw(30)(42*8-1 downto 41*8), w43 => Pw(30)(43*8-1 downto 42*8), w44 => Pw(30)(44*8-1 downto 43*8), w45 => Pw(30)(45*8-1 downto 44*8), w46 => Pw(30)(46*8-1 downto 45*8), w47 => Pw(30)(47*8-1 downto 46*8), w48 => Pw(30)(48*8-1 downto 47*8),  
w49 => Pw(30)(49*8-1 downto 48*8), w50 => Pw(30)(50*8-1 downto 49*8), w51 => Pw(30)(51*8-1 downto 50*8), w52 => Pw(30)(52*8-1 downto 51*8), w53 => Pw(30)(53*8-1 downto 52*8), w54 => Pw(30)(54*8-1 downto 53*8), w55 => Pw(30)(55*8-1 downto 54*8), w56 => Pw(30)(56*8-1 downto 55*8),  
w57 => Pw(30)(57*8-1 downto 56*8), w58 => Pw(30)(58*8-1 downto 57*8), w59 => Pw(30)(59*8-1 downto 58*8), w60 => Pw(30)(60*8-1 downto 59*8), w61 => Pw(30)(61*8-1 downto 60*8), w62 => Pw(30)(62*8-1 downto 61*8), w63 => Pw(30)(63*8-1 downto 62*8), w64 => Pw(30)(64*8-1 downto 63*8), 
w65 => Pw(30)( 65*8-1 downto  64*8), w66 => Pw(30)( 66*8-1 downto  65*8), w67 => Pw(30)( 67*8-1 downto  66*8), w68 => Pw(30)( 68*8-1 downto  67*8), w69 => Pw(30)( 69*8-1 downto  68*8), w70 => Pw(30)( 70*8-1 downto  69*8), w71 => Pw(30)( 71*8-1 downto  70*8), w72 => Pw(30)( 72*8-1 downto  71*8), 
w73 => Pw(30)( 73*8-1 downto  72*8), w74 => Pw(30)( 74*8-1 downto  73*8), w75 => Pw(30)( 75*8-1 downto  74*8), w76 => Pw(30)( 76*8-1 downto  75*8), w77 => Pw(30)( 77*8-1 downto  76*8), w78 => Pw(30)( 78*8-1 downto  77*8), w79 => Pw(30)( 79*8-1 downto  78*8), w80 => Pw(30)( 80*8-1 downto  79*8), 
w81 => Pw(30)( 81*8-1 downto  80*8), w82 => Pw(30)( 82*8-1 downto  81*8), w83 => Pw(30)( 83*8-1 downto  82*8), w84 => Pw(30)( 84*8-1 downto  83*8), w85 => Pw(30)( 85*8-1 downto  84*8), w86 => Pw(30)( 86*8-1 downto  85*8), w87 => Pw(30)( 87*8-1 downto  86*8), w88 => Pw(30)( 88*8-1 downto  87*8), 
w89 => Pw(30)( 89*8-1 downto  88*8), w90 => Pw(30)( 90*8-1 downto  89*8), w91 => Pw(30)( 91*8-1 downto  90*8), w92 => Pw(30)( 92*8-1 downto  91*8), w93 => Pw(30)( 93*8-1 downto  92*8), w94 => Pw(30)( 94*8-1 downto  93*8), w95 => Pw(30)( 95*8-1 downto  94*8), w96 => Pw(30)( 96*8-1 downto  95*8), 
w97 => Pw(30)( 97*8-1 downto  96*8), w98 => Pw(30)( 98*8-1 downto  97*8), w99 => Pw(30)( 99*8-1 downto  98*8), w100=> Pw(30)(100*8-1 downto  99*8), w101=> Pw(30)(101*8-1 downto 100*8), w102=> Pw(30)(102*8-1 downto 101*8), w103=> Pw(30)(103*8-1 downto 102*8), w104=> Pw(30)(104*8-1 downto 103*8), 
w105=> Pw(30)(105*8-1 downto 104*8), w106=> Pw(30)(106*8-1 downto 105*8), w107=> Pw(30)(107*8-1 downto 106*8), w108=> Pw(30)(108*8-1 downto 107*8), w109=> Pw(30)(109*8-1 downto 108*8), w110=> Pw(30)(110*8-1 downto 109*8), w111=> Pw(30)(111*8-1 downto 110*8), w112=> Pw(30)(112*8-1 downto 111*8), 
w113=> Pw(30)(113*8-1 downto 112*8), w114=> Pw(30)(114*8-1 downto 113*8), w115=> Pw(30)(115*8-1 downto 114*8), w116=> Pw(30)(116*8-1 downto 115*8), w117=> Pw(30)(117*8-1 downto 116*8), w118=> Pw(30)(118*8-1 downto 117*8), w119=> Pw(30)(119*8-1 downto 118*8), w120=> Pw(30)(120*8-1 downto 119*8), 
w121=> Pw(30)(121*8-1 downto 120*8), w122=> Pw(30)(122*8-1 downto 121*8), w123=> Pw(30)(123*8-1 downto 122*8), w124=> Pw(30)(124*8-1 downto 123*8), w125=> Pw(30)(125*8-1 downto 124*8), w126=> Pw(30)(126*8-1 downto 125*8), w127=> Pw(30)(127*8-1 downto 126*8), w128=> Pw(30)(128*8-1 downto 127*8), 

           d_out   => pca_d30_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_31_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(31)(     7 downto    0), w02 => Pw(31)( 2*8-1 downto    8), w03 => Pw(31)( 3*8-1 downto  2*8), w04 => Pw(31)( 4*8-1 downto  3*8), w05 => Pw(31)( 5*8-1 downto  4*8), w06 => Pw(31)( 6*8-1 downto  5*8), w07 => Pw(31)( 7*8-1 downto  6*8), w08 => Pw(31)( 8*8-1 downto  7*8),  
w09 => Pw(31)( 9*8-1 downto  8*8), w10 => Pw(31)(10*8-1 downto  9*8), w11 => Pw(31)(11*8-1 downto 10*8), w12 => Pw(31)(12*8-1 downto 11*8), w13 => Pw(31)(13*8-1 downto 12*8), w14 => Pw(31)(14*8-1 downto 13*8), w15 => Pw(31)(15*8-1 downto 14*8), w16 => Pw(31)(16*8-1 downto 15*8),  
w17 => Pw(31)(17*8-1 downto 16*8), w18 => Pw(31)(18*8-1 downto 17*8), w19 => Pw(31)(19*8-1 downto 18*8), w20 => Pw(31)(20*8-1 downto 19*8), w21 => Pw(31)(21*8-1 downto 20*8), w22 => Pw(31)(22*8-1 downto 21*8), w23 => Pw(31)(23*8-1 downto 22*8), w24 => Pw(31)(24*8-1 downto 23*8),  
w25 => Pw(31)(25*8-1 downto 24*8), w26 => Pw(31)(26*8-1 downto 25*8), w27 => Pw(31)(27*8-1 downto 26*8), w28 => Pw(31)(28*8-1 downto 27*8), w29 => Pw(31)(29*8-1 downto 28*8), w30 => Pw(31)(30*8-1 downto 29*8), w31 => Pw(31)(31*8-1 downto 30*8), w32 => Pw(31)(32*8-1 downto 31*8),  
w33 => Pw(31)(33*8-1 downto 32*8), w34 => Pw(31)(34*8-1 downto 33*8), w35 => Pw(31)(35*8-1 downto 34*8), w36 => Pw(31)(36*8-1 downto 35*8), w37 => Pw(31)(37*8-1 downto 36*8), w38 => Pw(31)(38*8-1 downto 37*8), w39 => Pw(31)(39*8-1 downto 38*8), w40 => Pw(31)(40*8-1 downto 39*8),  
w41 => Pw(31)(41*8-1 downto 40*8), w42 => Pw(31)(42*8-1 downto 41*8), w43 => Pw(31)(43*8-1 downto 42*8), w44 => Pw(31)(44*8-1 downto 43*8), w45 => Pw(31)(45*8-1 downto 44*8), w46 => Pw(31)(46*8-1 downto 45*8), w47 => Pw(31)(47*8-1 downto 46*8), w48 => Pw(31)(48*8-1 downto 47*8),  
w49 => Pw(31)(49*8-1 downto 48*8), w50 => Pw(31)(50*8-1 downto 49*8), w51 => Pw(31)(51*8-1 downto 50*8), w52 => Pw(31)(52*8-1 downto 51*8), w53 => Pw(31)(53*8-1 downto 52*8), w54 => Pw(31)(54*8-1 downto 53*8), w55 => Pw(31)(55*8-1 downto 54*8), w56 => Pw(31)(56*8-1 downto 55*8),  
w57 => Pw(31)(57*8-1 downto 56*8), w58 => Pw(31)(58*8-1 downto 57*8), w59 => Pw(31)(59*8-1 downto 58*8), w60 => Pw(31)(60*8-1 downto 59*8), w61 => Pw(31)(61*8-1 downto 60*8), w62 => Pw(31)(62*8-1 downto 61*8), w63 => Pw(31)(63*8-1 downto 62*8), w64 => Pw(31)(64*8-1 downto 63*8), 
w65 => Pw(31)( 65*8-1 downto  64*8), w66 => Pw(31)( 66*8-1 downto  65*8), w67 => Pw(31)( 67*8-1 downto  66*8), w68 => Pw(31)( 68*8-1 downto  67*8), w69 => Pw(31)( 69*8-1 downto  68*8), w70 => Pw(31)( 70*8-1 downto  69*8), w71 => Pw(31)( 71*8-1 downto  70*8), w72 => Pw(31)( 72*8-1 downto  71*8), 
w73 => Pw(31)( 73*8-1 downto  72*8), w74 => Pw(31)( 74*8-1 downto  73*8), w75 => Pw(31)( 75*8-1 downto  74*8), w76 => Pw(31)( 76*8-1 downto  75*8), w77 => Pw(31)( 77*8-1 downto  76*8), w78 => Pw(31)( 78*8-1 downto  77*8), w79 => Pw(31)( 79*8-1 downto  78*8), w80 => Pw(31)( 80*8-1 downto  79*8), 
w81 => Pw(31)( 81*8-1 downto  80*8), w82 => Pw(31)( 82*8-1 downto  81*8), w83 => Pw(31)( 83*8-1 downto  82*8), w84 => Pw(31)( 84*8-1 downto  83*8), w85 => Pw(31)( 85*8-1 downto  84*8), w86 => Pw(31)( 86*8-1 downto  85*8), w87 => Pw(31)( 87*8-1 downto  86*8), w88 => Pw(31)( 88*8-1 downto  87*8), 
w89 => Pw(31)( 89*8-1 downto  88*8), w90 => Pw(31)( 90*8-1 downto  89*8), w91 => Pw(31)( 91*8-1 downto  90*8), w92 => Pw(31)( 92*8-1 downto  91*8), w93 => Pw(31)( 93*8-1 downto  92*8), w94 => Pw(31)( 94*8-1 downto  93*8), w95 => Pw(31)( 95*8-1 downto  94*8), w96 => Pw(31)( 96*8-1 downto  95*8), 
w97 => Pw(31)( 97*8-1 downto  96*8), w98 => Pw(31)( 98*8-1 downto  97*8), w99 => Pw(31)( 99*8-1 downto  98*8), w100=> Pw(31)(100*8-1 downto  99*8), w101=> Pw(31)(101*8-1 downto 100*8), w102=> Pw(31)(102*8-1 downto 101*8), w103=> Pw(31)(103*8-1 downto 102*8), w104=> Pw(31)(104*8-1 downto 103*8), 
w105=> Pw(31)(105*8-1 downto 104*8), w106=> Pw(31)(106*8-1 downto 105*8), w107=> Pw(31)(107*8-1 downto 106*8), w108=> Pw(31)(108*8-1 downto 107*8), w109=> Pw(31)(109*8-1 downto 108*8), w110=> Pw(31)(110*8-1 downto 109*8), w111=> Pw(31)(111*8-1 downto 110*8), w112=> Pw(31)(112*8-1 downto 111*8), 
w113=> Pw(31)(113*8-1 downto 112*8), w114=> Pw(31)(114*8-1 downto 113*8), w115=> Pw(31)(115*8-1 downto 114*8), w116=> Pw(31)(116*8-1 downto 115*8), w117=> Pw(31)(117*8-1 downto 116*8), w118=> Pw(31)(118*8-1 downto 117*8), w119=> Pw(31)(119*8-1 downto 118*8), w120=> Pw(31)(120*8-1 downto 119*8), 
w121=> Pw(31)(121*8-1 downto 120*8), w122=> Pw(31)(122*8-1 downto 121*8), w123=> Pw(31)(123*8-1 downto 122*8), w124=> Pw(31)(124*8-1 downto 123*8), w125=> Pw(31)(125*8-1 downto 124*8), w126=> Pw(31)(126*8-1 downto 125*8), w127=> Pw(31)(127*8-1 downto 126*8), w128=> Pw(31)(128*8-1 downto 127*8), 

           d_out   => pca_d31_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_32_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(32)(     7 downto    0), w02 => Pw(32)( 2*8-1 downto    8), w03 => Pw(32)( 3*8-1 downto  2*8), w04 => Pw(32)( 4*8-1 downto  3*8), w05 => Pw(32)( 5*8-1 downto  4*8), w06 => Pw(32)( 6*8-1 downto  5*8), w07 => Pw(32)( 7*8-1 downto  6*8), w08 => Pw(32)( 8*8-1 downto  7*8),  
w09 => Pw(32)( 9*8-1 downto  8*8), w10 => Pw(32)(10*8-1 downto  9*8), w11 => Pw(32)(11*8-1 downto 10*8), w12 => Pw(32)(12*8-1 downto 11*8), w13 => Pw(32)(13*8-1 downto 12*8), w14 => Pw(32)(14*8-1 downto 13*8), w15 => Pw(32)(15*8-1 downto 14*8), w16 => Pw(32)(16*8-1 downto 15*8),  
w17 => Pw(32)(17*8-1 downto 16*8), w18 => Pw(32)(18*8-1 downto 17*8), w19 => Pw(32)(19*8-1 downto 18*8), w20 => Pw(32)(20*8-1 downto 19*8), w21 => Pw(32)(21*8-1 downto 20*8), w22 => Pw(32)(22*8-1 downto 21*8), w23 => Pw(32)(23*8-1 downto 22*8), w24 => Pw(32)(24*8-1 downto 23*8),  
w25 => Pw(32)(25*8-1 downto 24*8), w26 => Pw(32)(26*8-1 downto 25*8), w27 => Pw(32)(27*8-1 downto 26*8), w28 => Pw(32)(28*8-1 downto 27*8), w29 => Pw(32)(29*8-1 downto 28*8), w30 => Pw(32)(30*8-1 downto 29*8), w31 => Pw(32)(31*8-1 downto 30*8), w32 => Pw(32)(32*8-1 downto 31*8),  
w33 => Pw(32)(33*8-1 downto 32*8), w34 => Pw(32)(34*8-1 downto 33*8), w35 => Pw(32)(35*8-1 downto 34*8), w36 => Pw(32)(36*8-1 downto 35*8), w37 => Pw(32)(37*8-1 downto 36*8), w38 => Pw(32)(38*8-1 downto 37*8), w39 => Pw(32)(39*8-1 downto 38*8), w40 => Pw(32)(40*8-1 downto 39*8),  
w41 => Pw(32)(41*8-1 downto 40*8), w42 => Pw(32)(42*8-1 downto 41*8), w43 => Pw(32)(43*8-1 downto 42*8), w44 => Pw(32)(44*8-1 downto 43*8), w45 => Pw(32)(45*8-1 downto 44*8), w46 => Pw(32)(46*8-1 downto 45*8), w47 => Pw(32)(47*8-1 downto 46*8), w48 => Pw(32)(48*8-1 downto 47*8),  
w49 => Pw(32)(49*8-1 downto 48*8), w50 => Pw(32)(50*8-1 downto 49*8), w51 => Pw(32)(51*8-1 downto 50*8), w52 => Pw(32)(52*8-1 downto 51*8), w53 => Pw(32)(53*8-1 downto 52*8), w54 => Pw(32)(54*8-1 downto 53*8), w55 => Pw(32)(55*8-1 downto 54*8), w56 => Pw(32)(56*8-1 downto 55*8),  
w57 => Pw(32)(57*8-1 downto 56*8), w58 => Pw(32)(58*8-1 downto 57*8), w59 => Pw(32)(59*8-1 downto 58*8), w60 => Pw(32)(60*8-1 downto 59*8), w61 => Pw(32)(61*8-1 downto 60*8), w62 => Pw(32)(62*8-1 downto 61*8), w63 => Pw(32)(63*8-1 downto 62*8), w64 => Pw(32)(64*8-1 downto 63*8), 
w65 => Pw(32)( 65*8-1 downto  64*8), w66 => Pw(32)( 66*8-1 downto  65*8), w67 => Pw(32)( 67*8-1 downto  66*8), w68 => Pw(32)( 68*8-1 downto  67*8), w69 => Pw(32)( 69*8-1 downto  68*8), w70 => Pw(32)( 70*8-1 downto  69*8), w71 => Pw(32)( 71*8-1 downto  70*8), w72 => Pw(32)( 72*8-1 downto  71*8), 
w73 => Pw(32)( 73*8-1 downto  72*8), w74 => Pw(32)( 74*8-1 downto  73*8), w75 => Pw(32)( 75*8-1 downto  74*8), w76 => Pw(32)( 76*8-1 downto  75*8), w77 => Pw(32)( 77*8-1 downto  76*8), w78 => Pw(32)( 78*8-1 downto  77*8), w79 => Pw(32)( 79*8-1 downto  78*8), w80 => Pw(32)( 80*8-1 downto  79*8), 
w81 => Pw(32)( 81*8-1 downto  80*8), w82 => Pw(32)( 82*8-1 downto  81*8), w83 => Pw(32)( 83*8-1 downto  82*8), w84 => Pw(32)( 84*8-1 downto  83*8), w85 => Pw(32)( 85*8-1 downto  84*8), w86 => Pw(32)( 86*8-1 downto  85*8), w87 => Pw(32)( 87*8-1 downto  86*8), w88 => Pw(32)( 88*8-1 downto  87*8), 
w89 => Pw(32)( 89*8-1 downto  88*8), w90 => Pw(32)( 90*8-1 downto  89*8), w91 => Pw(32)( 91*8-1 downto  90*8), w92 => Pw(32)( 92*8-1 downto  91*8), w93 => Pw(32)( 93*8-1 downto  92*8), w94 => Pw(32)( 94*8-1 downto  93*8), w95 => Pw(32)( 95*8-1 downto  94*8), w96 => Pw(32)( 96*8-1 downto  95*8), 
w97 => Pw(32)( 97*8-1 downto  96*8), w98 => Pw(32)( 98*8-1 downto  97*8), w99 => Pw(32)( 99*8-1 downto  98*8), w100=> Pw(32)(100*8-1 downto  99*8), w101=> Pw(32)(101*8-1 downto 100*8), w102=> Pw(32)(102*8-1 downto 101*8), w103=> Pw(32)(103*8-1 downto 102*8), w104=> Pw(32)(104*8-1 downto 103*8), 
w105=> Pw(32)(105*8-1 downto 104*8), w106=> Pw(32)(106*8-1 downto 105*8), w107=> Pw(32)(107*8-1 downto 106*8), w108=> Pw(32)(108*8-1 downto 107*8), w109=> Pw(32)(109*8-1 downto 108*8), w110=> Pw(32)(110*8-1 downto 109*8), w111=> Pw(32)(111*8-1 downto 110*8), w112=> Pw(32)(112*8-1 downto 111*8), 
w113=> Pw(32)(113*8-1 downto 112*8), w114=> Pw(32)(114*8-1 downto 113*8), w115=> Pw(32)(115*8-1 downto 114*8), w116=> Pw(32)(116*8-1 downto 115*8), w117=> Pw(32)(117*8-1 downto 116*8), w118=> Pw(32)(118*8-1 downto 117*8), w119=> Pw(32)(119*8-1 downto 118*8), w120=> Pw(32)(120*8-1 downto 119*8), 
w121=> Pw(32)(121*8-1 downto 120*8), w122=> Pw(32)(122*8-1 downto 121*8), w123=> Pw(32)(123*8-1 downto 122*8), w124=> Pw(32)(124*8-1 downto 123*8), w125=> Pw(32)(125*8-1 downto 124*8), w126=> Pw(32)(126*8-1 downto 125*8), w127=> Pw(32)(127*8-1 downto 126*8), w128=> Pw(32)(128*8-1 downto 127*8), 

           d_out   => pca_d32_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_33_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(33)(     7 downto    0), w02 => Pw(33)( 2*8-1 downto    8), w03 => Pw(33)( 3*8-1 downto  2*8), w04 => Pw(33)( 4*8-1 downto  3*8), w05 => Pw(33)( 5*8-1 downto  4*8), w06 => Pw(33)( 6*8-1 downto  5*8), w07 => Pw(33)( 7*8-1 downto  6*8), w08 => Pw(33)( 8*8-1 downto  7*8),  
w09 => Pw(33)( 9*8-1 downto  8*8), w10 => Pw(33)(10*8-1 downto  9*8), w11 => Pw(33)(11*8-1 downto 10*8), w12 => Pw(33)(12*8-1 downto 11*8), w13 => Pw(33)(13*8-1 downto 12*8), w14 => Pw(33)(14*8-1 downto 13*8), w15 => Pw(33)(15*8-1 downto 14*8), w16 => Pw(33)(16*8-1 downto 15*8),  
w17 => Pw(33)(17*8-1 downto 16*8), w18 => Pw(33)(18*8-1 downto 17*8), w19 => Pw(33)(19*8-1 downto 18*8), w20 => Pw(33)(20*8-1 downto 19*8), w21 => Pw(33)(21*8-1 downto 20*8), w22 => Pw(33)(22*8-1 downto 21*8), w23 => Pw(33)(23*8-1 downto 22*8), w24 => Pw(33)(24*8-1 downto 23*8),  
w25 => Pw(33)(25*8-1 downto 24*8), w26 => Pw(33)(26*8-1 downto 25*8), w27 => Pw(33)(27*8-1 downto 26*8), w28 => Pw(33)(28*8-1 downto 27*8), w29 => Pw(33)(29*8-1 downto 28*8), w30 => Pw(33)(30*8-1 downto 29*8), w31 => Pw(33)(31*8-1 downto 30*8), w32 => Pw(33)(32*8-1 downto 31*8),  
w33 => Pw(33)(33*8-1 downto 32*8), w34 => Pw(33)(34*8-1 downto 33*8), w35 => Pw(33)(35*8-1 downto 34*8), w36 => Pw(33)(36*8-1 downto 35*8), w37 => Pw(33)(37*8-1 downto 36*8), w38 => Pw(33)(38*8-1 downto 37*8), w39 => Pw(33)(39*8-1 downto 38*8), w40 => Pw(33)(40*8-1 downto 39*8),  
w41 => Pw(33)(41*8-1 downto 40*8), w42 => Pw(33)(42*8-1 downto 41*8), w43 => Pw(33)(43*8-1 downto 42*8), w44 => Pw(33)(44*8-1 downto 43*8), w45 => Pw(33)(45*8-1 downto 44*8), w46 => Pw(33)(46*8-1 downto 45*8), w47 => Pw(33)(47*8-1 downto 46*8), w48 => Pw(33)(48*8-1 downto 47*8),  
w49 => Pw(33)(49*8-1 downto 48*8), w50 => Pw(33)(50*8-1 downto 49*8), w51 => Pw(33)(51*8-1 downto 50*8), w52 => Pw(33)(52*8-1 downto 51*8), w53 => Pw(33)(53*8-1 downto 52*8), w54 => Pw(33)(54*8-1 downto 53*8), w55 => Pw(33)(55*8-1 downto 54*8), w56 => Pw(33)(56*8-1 downto 55*8),  
w57 => Pw(33)(57*8-1 downto 56*8), w58 => Pw(33)(58*8-1 downto 57*8), w59 => Pw(33)(59*8-1 downto 58*8), w60 => Pw(33)(60*8-1 downto 59*8), w61 => Pw(33)(61*8-1 downto 60*8), w62 => Pw(33)(62*8-1 downto 61*8), w63 => Pw(33)(63*8-1 downto 62*8), w64 => Pw(33)(64*8-1 downto 63*8), 
w65 => Pw(33)( 65*8-1 downto  64*8), w66 => Pw(33)( 66*8-1 downto  65*8), w67 => Pw(33)( 67*8-1 downto  66*8), w68 => Pw(33)( 68*8-1 downto  67*8), w69 => Pw(33)( 69*8-1 downto  68*8), w70 => Pw(33)( 70*8-1 downto  69*8), w71 => Pw(33)( 71*8-1 downto  70*8), w72 => Pw(33)( 72*8-1 downto  71*8), 
w73 => Pw(33)( 73*8-1 downto  72*8), w74 => Pw(33)( 74*8-1 downto  73*8), w75 => Pw(33)( 75*8-1 downto  74*8), w76 => Pw(33)( 76*8-1 downto  75*8), w77 => Pw(33)( 77*8-1 downto  76*8), w78 => Pw(33)( 78*8-1 downto  77*8), w79 => Pw(33)( 79*8-1 downto  78*8), w80 => Pw(33)( 80*8-1 downto  79*8), 
w81 => Pw(33)( 81*8-1 downto  80*8), w82 => Pw(33)( 82*8-1 downto  81*8), w83 => Pw(33)( 83*8-1 downto  82*8), w84 => Pw(33)( 84*8-1 downto  83*8), w85 => Pw(33)( 85*8-1 downto  84*8), w86 => Pw(33)( 86*8-1 downto  85*8), w87 => Pw(33)( 87*8-1 downto  86*8), w88 => Pw(33)( 88*8-1 downto  87*8), 
w89 => Pw(33)( 89*8-1 downto  88*8), w90 => Pw(33)( 90*8-1 downto  89*8), w91 => Pw(33)( 91*8-1 downto  90*8), w92 => Pw(33)( 92*8-1 downto  91*8), w93 => Pw(33)( 93*8-1 downto  92*8), w94 => Pw(33)( 94*8-1 downto  93*8), w95 => Pw(33)( 95*8-1 downto  94*8), w96 => Pw(33)( 96*8-1 downto  95*8), 
w97 => Pw(33)( 97*8-1 downto  96*8), w98 => Pw(33)( 98*8-1 downto  97*8), w99 => Pw(33)( 99*8-1 downto  98*8), w100=> Pw(33)(100*8-1 downto  99*8), w101=> Pw(33)(101*8-1 downto 100*8), w102=> Pw(33)(102*8-1 downto 101*8), w103=> Pw(33)(103*8-1 downto 102*8), w104=> Pw(33)(104*8-1 downto 103*8), 
w105=> Pw(33)(105*8-1 downto 104*8), w106=> Pw(33)(106*8-1 downto 105*8), w107=> Pw(33)(107*8-1 downto 106*8), w108=> Pw(33)(108*8-1 downto 107*8), w109=> Pw(33)(109*8-1 downto 108*8), w110=> Pw(33)(110*8-1 downto 109*8), w111=> Pw(33)(111*8-1 downto 110*8), w112=> Pw(33)(112*8-1 downto 111*8), 
w113=> Pw(33)(113*8-1 downto 112*8), w114=> Pw(33)(114*8-1 downto 113*8), w115=> Pw(33)(115*8-1 downto 114*8), w116=> Pw(33)(116*8-1 downto 115*8), w117=> Pw(33)(117*8-1 downto 116*8), w118=> Pw(33)(118*8-1 downto 117*8), w119=> Pw(33)(119*8-1 downto 118*8), w120=> Pw(33)(120*8-1 downto 119*8), 
w121=> Pw(33)(121*8-1 downto 120*8), w122=> Pw(33)(122*8-1 downto 121*8), w123=> Pw(33)(123*8-1 downto 122*8), w124=> Pw(33)(124*8-1 downto 123*8), w125=> Pw(33)(125*8-1 downto 124*8), w126=> Pw(33)(126*8-1 downto 125*8), w127=> Pw(33)(127*8-1 downto 126*8), w128=> Pw(33)(128*8-1 downto 127*8), 

           d_out   => pca_d33_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_34_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(34)(     7 downto    0), w02 => Pw(34)( 2*8-1 downto    8), w03 => Pw(34)( 3*8-1 downto  2*8), w04 => Pw(34)( 4*8-1 downto  3*8), w05 => Pw(34)( 5*8-1 downto  4*8), w06 => Pw(34)( 6*8-1 downto  5*8), w07 => Pw(34)( 7*8-1 downto  6*8), w08 => Pw(34)( 8*8-1 downto  7*8),  
w09 => Pw(34)( 9*8-1 downto  8*8), w10 => Pw(34)(10*8-1 downto  9*8), w11 => Pw(34)(11*8-1 downto 10*8), w12 => Pw(34)(12*8-1 downto 11*8), w13 => Pw(34)(13*8-1 downto 12*8), w14 => Pw(34)(14*8-1 downto 13*8), w15 => Pw(34)(15*8-1 downto 14*8), w16 => Pw(34)(16*8-1 downto 15*8),  
w17 => Pw(34)(17*8-1 downto 16*8), w18 => Pw(34)(18*8-1 downto 17*8), w19 => Pw(34)(19*8-1 downto 18*8), w20 => Pw(34)(20*8-1 downto 19*8), w21 => Pw(34)(21*8-1 downto 20*8), w22 => Pw(34)(22*8-1 downto 21*8), w23 => Pw(34)(23*8-1 downto 22*8), w24 => Pw(34)(24*8-1 downto 23*8),  
w25 => Pw(34)(25*8-1 downto 24*8), w26 => Pw(34)(26*8-1 downto 25*8), w27 => Pw(34)(27*8-1 downto 26*8), w28 => Pw(34)(28*8-1 downto 27*8), w29 => Pw(34)(29*8-1 downto 28*8), w30 => Pw(34)(30*8-1 downto 29*8), w31 => Pw(34)(31*8-1 downto 30*8), w32 => Pw(34)(32*8-1 downto 31*8),  
w33 => Pw(34)(33*8-1 downto 32*8), w34 => Pw(34)(34*8-1 downto 33*8), w35 => Pw(34)(35*8-1 downto 34*8), w36 => Pw(34)(36*8-1 downto 35*8), w37 => Pw(34)(37*8-1 downto 36*8), w38 => Pw(34)(38*8-1 downto 37*8), w39 => Pw(34)(39*8-1 downto 38*8), w40 => Pw(34)(40*8-1 downto 39*8),  
w41 => Pw(34)(41*8-1 downto 40*8), w42 => Pw(34)(42*8-1 downto 41*8), w43 => Pw(34)(43*8-1 downto 42*8), w44 => Pw(34)(44*8-1 downto 43*8), w45 => Pw(34)(45*8-1 downto 44*8), w46 => Pw(34)(46*8-1 downto 45*8), w47 => Pw(34)(47*8-1 downto 46*8), w48 => Pw(34)(48*8-1 downto 47*8),  
w49 => Pw(34)(49*8-1 downto 48*8), w50 => Pw(34)(50*8-1 downto 49*8), w51 => Pw(34)(51*8-1 downto 50*8), w52 => Pw(34)(52*8-1 downto 51*8), w53 => Pw(34)(53*8-1 downto 52*8), w54 => Pw(34)(54*8-1 downto 53*8), w55 => Pw(34)(55*8-1 downto 54*8), w56 => Pw(34)(56*8-1 downto 55*8),  
w57 => Pw(34)(57*8-1 downto 56*8), w58 => Pw(34)(58*8-1 downto 57*8), w59 => Pw(34)(59*8-1 downto 58*8), w60 => Pw(34)(60*8-1 downto 59*8), w61 => Pw(34)(61*8-1 downto 60*8), w62 => Pw(34)(62*8-1 downto 61*8), w63 => Pw(34)(63*8-1 downto 62*8), w64 => Pw(34)(64*8-1 downto 63*8), 
w65 => Pw(34)( 65*8-1 downto  64*8), w66 => Pw(34)( 66*8-1 downto  65*8), w67 => Pw(34)( 67*8-1 downto  66*8), w68 => Pw(34)( 68*8-1 downto  67*8), w69 => Pw(34)( 69*8-1 downto  68*8), w70 => Pw(34)( 70*8-1 downto  69*8), w71 => Pw(34)( 71*8-1 downto  70*8), w72 => Pw(34)( 72*8-1 downto  71*8), 
w73 => Pw(34)( 73*8-1 downto  72*8), w74 => Pw(34)( 74*8-1 downto  73*8), w75 => Pw(34)( 75*8-1 downto  74*8), w76 => Pw(34)( 76*8-1 downto  75*8), w77 => Pw(34)( 77*8-1 downto  76*8), w78 => Pw(34)( 78*8-1 downto  77*8), w79 => Pw(34)( 79*8-1 downto  78*8), w80 => Pw(34)( 80*8-1 downto  79*8), 
w81 => Pw(34)( 81*8-1 downto  80*8), w82 => Pw(34)( 82*8-1 downto  81*8), w83 => Pw(34)( 83*8-1 downto  82*8), w84 => Pw(34)( 84*8-1 downto  83*8), w85 => Pw(34)( 85*8-1 downto  84*8), w86 => Pw(34)( 86*8-1 downto  85*8), w87 => Pw(34)( 87*8-1 downto  86*8), w88 => Pw(34)( 88*8-1 downto  87*8), 
w89 => Pw(34)( 89*8-1 downto  88*8), w90 => Pw(34)( 90*8-1 downto  89*8), w91 => Pw(34)( 91*8-1 downto  90*8), w92 => Pw(34)( 92*8-1 downto  91*8), w93 => Pw(34)( 93*8-1 downto  92*8), w94 => Pw(34)( 94*8-1 downto  93*8), w95 => Pw(34)( 95*8-1 downto  94*8), w96 => Pw(34)( 96*8-1 downto  95*8), 
w97 => Pw(34)( 97*8-1 downto  96*8), w98 => Pw(34)( 98*8-1 downto  97*8), w99 => Pw(34)( 99*8-1 downto  98*8), w100=> Pw(34)(100*8-1 downto  99*8), w101=> Pw(34)(101*8-1 downto 100*8), w102=> Pw(34)(102*8-1 downto 101*8), w103=> Pw(34)(103*8-1 downto 102*8), w104=> Pw(34)(104*8-1 downto 103*8), 
w105=> Pw(34)(105*8-1 downto 104*8), w106=> Pw(34)(106*8-1 downto 105*8), w107=> Pw(34)(107*8-1 downto 106*8), w108=> Pw(34)(108*8-1 downto 107*8), w109=> Pw(34)(109*8-1 downto 108*8), w110=> Pw(34)(110*8-1 downto 109*8), w111=> Pw(34)(111*8-1 downto 110*8), w112=> Pw(34)(112*8-1 downto 111*8), 
w113=> Pw(34)(113*8-1 downto 112*8), w114=> Pw(34)(114*8-1 downto 113*8), w115=> Pw(34)(115*8-1 downto 114*8), w116=> Pw(34)(116*8-1 downto 115*8), w117=> Pw(34)(117*8-1 downto 116*8), w118=> Pw(34)(118*8-1 downto 117*8), w119=> Pw(34)(119*8-1 downto 118*8), w120=> Pw(34)(120*8-1 downto 119*8), 
w121=> Pw(34)(121*8-1 downto 120*8), w122=> Pw(34)(122*8-1 downto 121*8), w123=> Pw(34)(123*8-1 downto 122*8), w124=> Pw(34)(124*8-1 downto 123*8), w125=> Pw(34)(125*8-1 downto 124*8), w126=> Pw(34)(126*8-1 downto 125*8), w127=> Pw(34)(127*8-1 downto 126*8), w128=> Pw(34)(128*8-1 downto 127*8), 

           d_out   => pca_d34_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_35_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(35)(     7 downto    0), w02 => Pw(35)( 2*8-1 downto    8), w03 => Pw(35)( 3*8-1 downto  2*8), w04 => Pw(35)( 4*8-1 downto  3*8), w05 => Pw(35)( 5*8-1 downto  4*8), w06 => Pw(35)( 6*8-1 downto  5*8), w07 => Pw(35)( 7*8-1 downto  6*8), w08 => Pw(35)( 8*8-1 downto  7*8),  
w09 => Pw(35)( 9*8-1 downto  8*8), w10 => Pw(35)(10*8-1 downto  9*8), w11 => Pw(35)(11*8-1 downto 10*8), w12 => Pw(35)(12*8-1 downto 11*8), w13 => Pw(35)(13*8-1 downto 12*8), w14 => Pw(35)(14*8-1 downto 13*8), w15 => Pw(35)(15*8-1 downto 14*8), w16 => Pw(35)(16*8-1 downto 15*8),  
w17 => Pw(35)(17*8-1 downto 16*8), w18 => Pw(35)(18*8-1 downto 17*8), w19 => Pw(35)(19*8-1 downto 18*8), w20 => Pw(35)(20*8-1 downto 19*8), w21 => Pw(35)(21*8-1 downto 20*8), w22 => Pw(35)(22*8-1 downto 21*8), w23 => Pw(35)(23*8-1 downto 22*8), w24 => Pw(35)(24*8-1 downto 23*8),  
w25 => Pw(35)(25*8-1 downto 24*8), w26 => Pw(35)(26*8-1 downto 25*8), w27 => Pw(35)(27*8-1 downto 26*8), w28 => Pw(35)(28*8-1 downto 27*8), w29 => Pw(35)(29*8-1 downto 28*8), w30 => Pw(35)(30*8-1 downto 29*8), w31 => Pw(35)(31*8-1 downto 30*8), w32 => Pw(35)(32*8-1 downto 31*8),  
w33 => Pw(35)(33*8-1 downto 32*8), w34 => Pw(35)(34*8-1 downto 33*8), w35 => Pw(35)(35*8-1 downto 34*8), w36 => Pw(35)(36*8-1 downto 35*8), w37 => Pw(35)(37*8-1 downto 36*8), w38 => Pw(35)(38*8-1 downto 37*8), w39 => Pw(35)(39*8-1 downto 38*8), w40 => Pw(35)(40*8-1 downto 39*8),  
w41 => Pw(35)(41*8-1 downto 40*8), w42 => Pw(35)(42*8-1 downto 41*8), w43 => Pw(35)(43*8-1 downto 42*8), w44 => Pw(35)(44*8-1 downto 43*8), w45 => Pw(35)(45*8-1 downto 44*8), w46 => Pw(35)(46*8-1 downto 45*8), w47 => Pw(35)(47*8-1 downto 46*8), w48 => Pw(35)(48*8-1 downto 47*8),  
w49 => Pw(35)(49*8-1 downto 48*8), w50 => Pw(35)(50*8-1 downto 49*8), w51 => Pw(35)(51*8-1 downto 50*8), w52 => Pw(35)(52*8-1 downto 51*8), w53 => Pw(35)(53*8-1 downto 52*8), w54 => Pw(35)(54*8-1 downto 53*8), w55 => Pw(35)(55*8-1 downto 54*8), w56 => Pw(35)(56*8-1 downto 55*8),  
w57 => Pw(35)(57*8-1 downto 56*8), w58 => Pw(35)(58*8-1 downto 57*8), w59 => Pw(35)(59*8-1 downto 58*8), w60 => Pw(35)(60*8-1 downto 59*8), w61 => Pw(35)(61*8-1 downto 60*8), w62 => Pw(35)(62*8-1 downto 61*8), w63 => Pw(35)(63*8-1 downto 62*8), w64 => Pw(35)(64*8-1 downto 63*8), 
w65 => Pw(35)( 65*8-1 downto  64*8), w66 => Pw(35)( 66*8-1 downto  65*8), w67 => Pw(35)( 67*8-1 downto  66*8), w68 => Pw(35)( 68*8-1 downto  67*8), w69 => Pw(35)( 69*8-1 downto  68*8), w70 => Pw(35)( 70*8-1 downto  69*8), w71 => Pw(35)( 71*8-1 downto  70*8), w72 => Pw(35)( 72*8-1 downto  71*8), 
w73 => Pw(35)( 73*8-1 downto  72*8), w74 => Pw(35)( 74*8-1 downto  73*8), w75 => Pw(35)( 75*8-1 downto  74*8), w76 => Pw(35)( 76*8-1 downto  75*8), w77 => Pw(35)( 77*8-1 downto  76*8), w78 => Pw(35)( 78*8-1 downto  77*8), w79 => Pw(35)( 79*8-1 downto  78*8), w80 => Pw(35)( 80*8-1 downto  79*8), 
w81 => Pw(35)( 81*8-1 downto  80*8), w82 => Pw(35)( 82*8-1 downto  81*8), w83 => Pw(35)( 83*8-1 downto  82*8), w84 => Pw(35)( 84*8-1 downto  83*8), w85 => Pw(35)( 85*8-1 downto  84*8), w86 => Pw(35)( 86*8-1 downto  85*8), w87 => Pw(35)( 87*8-1 downto  86*8), w88 => Pw(35)( 88*8-1 downto  87*8), 
w89 => Pw(35)( 89*8-1 downto  88*8), w90 => Pw(35)( 90*8-1 downto  89*8), w91 => Pw(35)( 91*8-1 downto  90*8), w92 => Pw(35)( 92*8-1 downto  91*8), w93 => Pw(35)( 93*8-1 downto  92*8), w94 => Pw(35)( 94*8-1 downto  93*8), w95 => Pw(35)( 95*8-1 downto  94*8), w96 => Pw(35)( 96*8-1 downto  95*8), 
w97 => Pw(35)( 97*8-1 downto  96*8), w98 => Pw(35)( 98*8-1 downto  97*8), w99 => Pw(35)( 99*8-1 downto  98*8), w100=> Pw(35)(100*8-1 downto  99*8), w101=> Pw(35)(101*8-1 downto 100*8), w102=> Pw(35)(102*8-1 downto 101*8), w103=> Pw(35)(103*8-1 downto 102*8), w104=> Pw(35)(104*8-1 downto 103*8), 
w105=> Pw(35)(105*8-1 downto 104*8), w106=> Pw(35)(106*8-1 downto 105*8), w107=> Pw(35)(107*8-1 downto 106*8), w108=> Pw(35)(108*8-1 downto 107*8), w109=> Pw(35)(109*8-1 downto 108*8), w110=> Pw(35)(110*8-1 downto 109*8), w111=> Pw(35)(111*8-1 downto 110*8), w112=> Pw(35)(112*8-1 downto 111*8), 
w113=> Pw(35)(113*8-1 downto 112*8), w114=> Pw(35)(114*8-1 downto 113*8), w115=> Pw(35)(115*8-1 downto 114*8), w116=> Pw(35)(116*8-1 downto 115*8), w117=> Pw(35)(117*8-1 downto 116*8), w118=> Pw(35)(118*8-1 downto 117*8), w119=> Pw(35)(119*8-1 downto 118*8), w120=> Pw(35)(120*8-1 downto 119*8), 
w121=> Pw(35)(121*8-1 downto 120*8), w122=> Pw(35)(122*8-1 downto 121*8), w123=> Pw(35)(123*8-1 downto 122*8), w124=> Pw(35)(124*8-1 downto 123*8), w125=> Pw(35)(125*8-1 downto 124*8), w126=> Pw(35)(126*8-1 downto 125*8), w127=> Pw(35)(127*8-1 downto 126*8), w128=> Pw(35)(128*8-1 downto 127*8), 

           d_out   => pca_d35_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_36_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(36)(     7 downto    0), w02 => Pw(36)( 2*8-1 downto    8), w03 => Pw(36)( 3*8-1 downto  2*8), w04 => Pw(36)( 4*8-1 downto  3*8), w05 => Pw(36)( 5*8-1 downto  4*8), w06 => Pw(36)( 6*8-1 downto  5*8), w07 => Pw(36)( 7*8-1 downto  6*8), w08 => Pw(36)( 8*8-1 downto  7*8),  
w09 => Pw(36)( 9*8-1 downto  8*8), w10 => Pw(36)(10*8-1 downto  9*8), w11 => Pw(36)(11*8-1 downto 10*8), w12 => Pw(36)(12*8-1 downto 11*8), w13 => Pw(36)(13*8-1 downto 12*8), w14 => Pw(36)(14*8-1 downto 13*8), w15 => Pw(36)(15*8-1 downto 14*8), w16 => Pw(36)(16*8-1 downto 15*8),  
w17 => Pw(36)(17*8-1 downto 16*8), w18 => Pw(36)(18*8-1 downto 17*8), w19 => Pw(36)(19*8-1 downto 18*8), w20 => Pw(36)(20*8-1 downto 19*8), w21 => Pw(36)(21*8-1 downto 20*8), w22 => Pw(36)(22*8-1 downto 21*8), w23 => Pw(36)(23*8-1 downto 22*8), w24 => Pw(36)(24*8-1 downto 23*8),  
w25 => Pw(36)(25*8-1 downto 24*8), w26 => Pw(36)(26*8-1 downto 25*8), w27 => Pw(36)(27*8-1 downto 26*8), w28 => Pw(36)(28*8-1 downto 27*8), w29 => Pw(36)(29*8-1 downto 28*8), w30 => Pw(36)(30*8-1 downto 29*8), w31 => Pw(36)(31*8-1 downto 30*8), w32 => Pw(36)(32*8-1 downto 31*8),  
w33 => Pw(36)(33*8-1 downto 32*8), w34 => Pw(36)(34*8-1 downto 33*8), w35 => Pw(36)(35*8-1 downto 34*8), w36 => Pw(36)(36*8-1 downto 35*8), w37 => Pw(36)(37*8-1 downto 36*8), w38 => Pw(36)(38*8-1 downto 37*8), w39 => Pw(36)(39*8-1 downto 38*8), w40 => Pw(36)(40*8-1 downto 39*8),  
w41 => Pw(36)(41*8-1 downto 40*8), w42 => Pw(36)(42*8-1 downto 41*8), w43 => Pw(36)(43*8-1 downto 42*8), w44 => Pw(36)(44*8-1 downto 43*8), w45 => Pw(36)(45*8-1 downto 44*8), w46 => Pw(36)(46*8-1 downto 45*8), w47 => Pw(36)(47*8-1 downto 46*8), w48 => Pw(36)(48*8-1 downto 47*8),  
w49 => Pw(36)(49*8-1 downto 48*8), w50 => Pw(36)(50*8-1 downto 49*8), w51 => Pw(36)(51*8-1 downto 50*8), w52 => Pw(36)(52*8-1 downto 51*8), w53 => Pw(36)(53*8-1 downto 52*8), w54 => Pw(36)(54*8-1 downto 53*8), w55 => Pw(36)(55*8-1 downto 54*8), w56 => Pw(36)(56*8-1 downto 55*8),  
w57 => Pw(36)(57*8-1 downto 56*8), w58 => Pw(36)(58*8-1 downto 57*8), w59 => Pw(36)(59*8-1 downto 58*8), w60 => Pw(36)(60*8-1 downto 59*8), w61 => Pw(36)(61*8-1 downto 60*8), w62 => Pw(36)(62*8-1 downto 61*8), w63 => Pw(36)(63*8-1 downto 62*8), w64 => Pw(36)(64*8-1 downto 63*8), 
w65 => Pw(36)( 65*8-1 downto  64*8), w66 => Pw(36)( 66*8-1 downto  65*8), w67 => Pw(36)( 67*8-1 downto  66*8), w68 => Pw(36)( 68*8-1 downto  67*8), w69 => Pw(36)( 69*8-1 downto  68*8), w70 => Pw(36)( 70*8-1 downto  69*8), w71 => Pw(36)( 71*8-1 downto  70*8), w72 => Pw(36)( 72*8-1 downto  71*8), 
w73 => Pw(36)( 73*8-1 downto  72*8), w74 => Pw(36)( 74*8-1 downto  73*8), w75 => Pw(36)( 75*8-1 downto  74*8), w76 => Pw(36)( 76*8-1 downto  75*8), w77 => Pw(36)( 77*8-1 downto  76*8), w78 => Pw(36)( 78*8-1 downto  77*8), w79 => Pw(36)( 79*8-1 downto  78*8), w80 => Pw(36)( 80*8-1 downto  79*8), 
w81 => Pw(36)( 81*8-1 downto  80*8), w82 => Pw(36)( 82*8-1 downto  81*8), w83 => Pw(36)( 83*8-1 downto  82*8), w84 => Pw(36)( 84*8-1 downto  83*8), w85 => Pw(36)( 85*8-1 downto  84*8), w86 => Pw(36)( 86*8-1 downto  85*8), w87 => Pw(36)( 87*8-1 downto  86*8), w88 => Pw(36)( 88*8-1 downto  87*8), 
w89 => Pw(36)( 89*8-1 downto  88*8), w90 => Pw(36)( 90*8-1 downto  89*8), w91 => Pw(36)( 91*8-1 downto  90*8), w92 => Pw(36)( 92*8-1 downto  91*8), w93 => Pw(36)( 93*8-1 downto  92*8), w94 => Pw(36)( 94*8-1 downto  93*8), w95 => Pw(36)( 95*8-1 downto  94*8), w96 => Pw(36)( 96*8-1 downto  95*8), 
w97 => Pw(36)( 97*8-1 downto  96*8), w98 => Pw(36)( 98*8-1 downto  97*8), w99 => Pw(36)( 99*8-1 downto  98*8), w100=> Pw(36)(100*8-1 downto  99*8), w101=> Pw(36)(101*8-1 downto 100*8), w102=> Pw(36)(102*8-1 downto 101*8), w103=> Pw(36)(103*8-1 downto 102*8), w104=> Pw(36)(104*8-1 downto 103*8), 
w105=> Pw(36)(105*8-1 downto 104*8), w106=> Pw(36)(106*8-1 downto 105*8), w107=> Pw(36)(107*8-1 downto 106*8), w108=> Pw(36)(108*8-1 downto 107*8), w109=> Pw(36)(109*8-1 downto 108*8), w110=> Pw(36)(110*8-1 downto 109*8), w111=> Pw(36)(111*8-1 downto 110*8), w112=> Pw(36)(112*8-1 downto 111*8), 
w113=> Pw(36)(113*8-1 downto 112*8), w114=> Pw(36)(114*8-1 downto 113*8), w115=> Pw(36)(115*8-1 downto 114*8), w116=> Pw(36)(116*8-1 downto 115*8), w117=> Pw(36)(117*8-1 downto 116*8), w118=> Pw(36)(118*8-1 downto 117*8), w119=> Pw(36)(119*8-1 downto 118*8), w120=> Pw(36)(120*8-1 downto 119*8), 
w121=> Pw(36)(121*8-1 downto 120*8), w122=> Pw(36)(122*8-1 downto 121*8), w123=> Pw(36)(123*8-1 downto 122*8), w124=> Pw(36)(124*8-1 downto 123*8), w125=> Pw(36)(125*8-1 downto 124*8), w126=> Pw(36)(126*8-1 downto 125*8), w127=> Pw(36)(127*8-1 downto 126*8), w128=> Pw(36)(128*8-1 downto 127*8), 

           d_out   => pca_d36_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_37_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(37)(     7 downto    0), w02 => Pw(37)( 2*8-1 downto    8), w03 => Pw(37)( 3*8-1 downto  2*8), w04 => Pw(37)( 4*8-1 downto  3*8), w05 => Pw(37)( 5*8-1 downto  4*8), w06 => Pw(37)( 6*8-1 downto  5*8), w07 => Pw(37)( 7*8-1 downto  6*8), w08 => Pw(37)( 8*8-1 downto  7*8),  
w09 => Pw(37)( 9*8-1 downto  8*8), w10 => Pw(37)(10*8-1 downto  9*8), w11 => Pw(37)(11*8-1 downto 10*8), w12 => Pw(37)(12*8-1 downto 11*8), w13 => Pw(37)(13*8-1 downto 12*8), w14 => Pw(37)(14*8-1 downto 13*8), w15 => Pw(37)(15*8-1 downto 14*8), w16 => Pw(37)(16*8-1 downto 15*8),  
w17 => Pw(37)(17*8-1 downto 16*8), w18 => Pw(37)(18*8-1 downto 17*8), w19 => Pw(37)(19*8-1 downto 18*8), w20 => Pw(37)(20*8-1 downto 19*8), w21 => Pw(37)(21*8-1 downto 20*8), w22 => Pw(37)(22*8-1 downto 21*8), w23 => Pw(37)(23*8-1 downto 22*8), w24 => Pw(37)(24*8-1 downto 23*8),  
w25 => Pw(37)(25*8-1 downto 24*8), w26 => Pw(37)(26*8-1 downto 25*8), w27 => Pw(37)(27*8-1 downto 26*8), w28 => Pw(37)(28*8-1 downto 27*8), w29 => Pw(37)(29*8-1 downto 28*8), w30 => Pw(37)(30*8-1 downto 29*8), w31 => Pw(37)(31*8-1 downto 30*8), w32 => Pw(37)(32*8-1 downto 31*8),  
w33 => Pw(37)(33*8-1 downto 32*8), w34 => Pw(37)(34*8-1 downto 33*8), w35 => Pw(37)(35*8-1 downto 34*8), w36 => Pw(37)(36*8-1 downto 35*8), w37 => Pw(37)(37*8-1 downto 36*8), w38 => Pw(37)(38*8-1 downto 37*8), w39 => Pw(37)(39*8-1 downto 38*8), w40 => Pw(37)(40*8-1 downto 39*8),  
w41 => Pw(37)(41*8-1 downto 40*8), w42 => Pw(37)(42*8-1 downto 41*8), w43 => Pw(37)(43*8-1 downto 42*8), w44 => Pw(37)(44*8-1 downto 43*8), w45 => Pw(37)(45*8-1 downto 44*8), w46 => Pw(37)(46*8-1 downto 45*8), w47 => Pw(37)(47*8-1 downto 46*8), w48 => Pw(37)(48*8-1 downto 47*8),  
w49 => Pw(37)(49*8-1 downto 48*8), w50 => Pw(37)(50*8-1 downto 49*8), w51 => Pw(37)(51*8-1 downto 50*8), w52 => Pw(37)(52*8-1 downto 51*8), w53 => Pw(37)(53*8-1 downto 52*8), w54 => Pw(37)(54*8-1 downto 53*8), w55 => Pw(37)(55*8-1 downto 54*8), w56 => Pw(37)(56*8-1 downto 55*8),  
w57 => Pw(37)(57*8-1 downto 56*8), w58 => Pw(37)(58*8-1 downto 57*8), w59 => Pw(37)(59*8-1 downto 58*8), w60 => Pw(37)(60*8-1 downto 59*8), w61 => Pw(37)(61*8-1 downto 60*8), w62 => Pw(37)(62*8-1 downto 61*8), w63 => Pw(37)(63*8-1 downto 62*8), w64 => Pw(37)(64*8-1 downto 63*8), 
w65 => Pw(37)( 65*8-1 downto  64*8), w66 => Pw(37)( 66*8-1 downto  65*8), w67 => Pw(37)( 67*8-1 downto  66*8), w68 => Pw(37)( 68*8-1 downto  67*8), w69 => Pw(37)( 69*8-1 downto  68*8), w70 => Pw(37)( 70*8-1 downto  69*8), w71 => Pw(37)( 71*8-1 downto  70*8), w72 => Pw(37)( 72*8-1 downto  71*8), 
w73 => Pw(37)( 73*8-1 downto  72*8), w74 => Pw(37)( 74*8-1 downto  73*8), w75 => Pw(37)( 75*8-1 downto  74*8), w76 => Pw(37)( 76*8-1 downto  75*8), w77 => Pw(37)( 77*8-1 downto  76*8), w78 => Pw(37)( 78*8-1 downto  77*8), w79 => Pw(37)( 79*8-1 downto  78*8), w80 => Pw(37)( 80*8-1 downto  79*8), 
w81 => Pw(37)( 81*8-1 downto  80*8), w82 => Pw(37)( 82*8-1 downto  81*8), w83 => Pw(37)( 83*8-1 downto  82*8), w84 => Pw(37)( 84*8-1 downto  83*8), w85 => Pw(37)( 85*8-1 downto  84*8), w86 => Pw(37)( 86*8-1 downto  85*8), w87 => Pw(37)( 87*8-1 downto  86*8), w88 => Pw(37)( 88*8-1 downto  87*8), 
w89 => Pw(37)( 89*8-1 downto  88*8), w90 => Pw(37)( 90*8-1 downto  89*8), w91 => Pw(37)( 91*8-1 downto  90*8), w92 => Pw(37)( 92*8-1 downto  91*8), w93 => Pw(37)( 93*8-1 downto  92*8), w94 => Pw(37)( 94*8-1 downto  93*8), w95 => Pw(37)( 95*8-1 downto  94*8), w96 => Pw(37)( 96*8-1 downto  95*8), 
w97 => Pw(37)( 97*8-1 downto  96*8), w98 => Pw(37)( 98*8-1 downto  97*8), w99 => Pw(37)( 99*8-1 downto  98*8), w100=> Pw(37)(100*8-1 downto  99*8), w101=> Pw(37)(101*8-1 downto 100*8), w102=> Pw(37)(102*8-1 downto 101*8), w103=> Pw(37)(103*8-1 downto 102*8), w104=> Pw(37)(104*8-1 downto 103*8), 
w105=> Pw(37)(105*8-1 downto 104*8), w106=> Pw(37)(106*8-1 downto 105*8), w107=> Pw(37)(107*8-1 downto 106*8), w108=> Pw(37)(108*8-1 downto 107*8), w109=> Pw(37)(109*8-1 downto 108*8), w110=> Pw(37)(110*8-1 downto 109*8), w111=> Pw(37)(111*8-1 downto 110*8), w112=> Pw(37)(112*8-1 downto 111*8), 
w113=> Pw(37)(113*8-1 downto 112*8), w114=> Pw(37)(114*8-1 downto 113*8), w115=> Pw(37)(115*8-1 downto 114*8), w116=> Pw(37)(116*8-1 downto 115*8), w117=> Pw(37)(117*8-1 downto 116*8), w118=> Pw(37)(118*8-1 downto 117*8), w119=> Pw(37)(119*8-1 downto 118*8), w120=> Pw(37)(120*8-1 downto 119*8), 
w121=> Pw(37)(121*8-1 downto 120*8), w122=> Pw(37)(122*8-1 downto 121*8), w123=> Pw(37)(123*8-1 downto 122*8), w124=> Pw(37)(124*8-1 downto 123*8), w125=> Pw(37)(125*8-1 downto 124*8), w126=> Pw(37)(126*8-1 downto 125*8), w127=> Pw(37)(127*8-1 downto 126*8), w128=> Pw(37)(128*8-1 downto 127*8), 

           d_out   => pca_d37_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_38_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(38)(     7 downto    0), w02 => Pw(38)( 2*8-1 downto    8), w03 => Pw(38)( 3*8-1 downto  2*8), w04 => Pw(38)( 4*8-1 downto  3*8), w05 => Pw(38)( 5*8-1 downto  4*8), w06 => Pw(38)( 6*8-1 downto  5*8), w07 => Pw(38)( 7*8-1 downto  6*8), w08 => Pw(38)( 8*8-1 downto  7*8),  
w09 => Pw(38)( 9*8-1 downto  8*8), w10 => Pw(38)(10*8-1 downto  9*8), w11 => Pw(38)(11*8-1 downto 10*8), w12 => Pw(38)(12*8-1 downto 11*8), w13 => Pw(38)(13*8-1 downto 12*8), w14 => Pw(38)(14*8-1 downto 13*8), w15 => Pw(38)(15*8-1 downto 14*8), w16 => Pw(38)(16*8-1 downto 15*8),  
w17 => Pw(38)(17*8-1 downto 16*8), w18 => Pw(38)(18*8-1 downto 17*8), w19 => Pw(38)(19*8-1 downto 18*8), w20 => Pw(38)(20*8-1 downto 19*8), w21 => Pw(38)(21*8-1 downto 20*8), w22 => Pw(38)(22*8-1 downto 21*8), w23 => Pw(38)(23*8-1 downto 22*8), w24 => Pw(38)(24*8-1 downto 23*8),  
w25 => Pw(38)(25*8-1 downto 24*8), w26 => Pw(38)(26*8-1 downto 25*8), w27 => Pw(38)(27*8-1 downto 26*8), w28 => Pw(38)(28*8-1 downto 27*8), w29 => Pw(38)(29*8-1 downto 28*8), w30 => Pw(38)(30*8-1 downto 29*8), w31 => Pw(38)(31*8-1 downto 30*8), w32 => Pw(38)(32*8-1 downto 31*8),  
w33 => Pw(38)(33*8-1 downto 32*8), w34 => Pw(38)(34*8-1 downto 33*8), w35 => Pw(38)(35*8-1 downto 34*8), w36 => Pw(38)(36*8-1 downto 35*8), w37 => Pw(38)(37*8-1 downto 36*8), w38 => Pw(38)(38*8-1 downto 37*8), w39 => Pw(38)(39*8-1 downto 38*8), w40 => Pw(38)(40*8-1 downto 39*8),  
w41 => Pw(38)(41*8-1 downto 40*8), w42 => Pw(38)(42*8-1 downto 41*8), w43 => Pw(38)(43*8-1 downto 42*8), w44 => Pw(38)(44*8-1 downto 43*8), w45 => Pw(38)(45*8-1 downto 44*8), w46 => Pw(38)(46*8-1 downto 45*8), w47 => Pw(38)(47*8-1 downto 46*8), w48 => Pw(38)(48*8-1 downto 47*8),  
w49 => Pw(38)(49*8-1 downto 48*8), w50 => Pw(38)(50*8-1 downto 49*8), w51 => Pw(38)(51*8-1 downto 50*8), w52 => Pw(38)(52*8-1 downto 51*8), w53 => Pw(38)(53*8-1 downto 52*8), w54 => Pw(38)(54*8-1 downto 53*8), w55 => Pw(38)(55*8-1 downto 54*8), w56 => Pw(38)(56*8-1 downto 55*8),  
w57 => Pw(38)(57*8-1 downto 56*8), w58 => Pw(38)(58*8-1 downto 57*8), w59 => Pw(38)(59*8-1 downto 58*8), w60 => Pw(38)(60*8-1 downto 59*8), w61 => Pw(38)(61*8-1 downto 60*8), w62 => Pw(38)(62*8-1 downto 61*8), w63 => Pw(38)(63*8-1 downto 62*8), w64 => Pw(38)(64*8-1 downto 63*8), 
w65 => Pw(38)( 65*8-1 downto  64*8), w66 => Pw(38)( 66*8-1 downto  65*8), w67 => Pw(38)( 67*8-1 downto  66*8), w68 => Pw(38)( 68*8-1 downto  67*8), w69 => Pw(38)( 69*8-1 downto  68*8), w70 => Pw(38)( 70*8-1 downto  69*8), w71 => Pw(38)( 71*8-1 downto  70*8), w72 => Pw(38)( 72*8-1 downto  71*8), 
w73 => Pw(38)( 73*8-1 downto  72*8), w74 => Pw(38)( 74*8-1 downto  73*8), w75 => Pw(38)( 75*8-1 downto  74*8), w76 => Pw(38)( 76*8-1 downto  75*8), w77 => Pw(38)( 77*8-1 downto  76*8), w78 => Pw(38)( 78*8-1 downto  77*8), w79 => Pw(38)( 79*8-1 downto  78*8), w80 => Pw(38)( 80*8-1 downto  79*8), 
w81 => Pw(38)( 81*8-1 downto  80*8), w82 => Pw(38)( 82*8-1 downto  81*8), w83 => Pw(38)( 83*8-1 downto  82*8), w84 => Pw(38)( 84*8-1 downto  83*8), w85 => Pw(38)( 85*8-1 downto  84*8), w86 => Pw(38)( 86*8-1 downto  85*8), w87 => Pw(38)( 87*8-1 downto  86*8), w88 => Pw(38)( 88*8-1 downto  87*8), 
w89 => Pw(38)( 89*8-1 downto  88*8), w90 => Pw(38)( 90*8-1 downto  89*8), w91 => Pw(38)( 91*8-1 downto  90*8), w92 => Pw(38)( 92*8-1 downto  91*8), w93 => Pw(38)( 93*8-1 downto  92*8), w94 => Pw(38)( 94*8-1 downto  93*8), w95 => Pw(38)( 95*8-1 downto  94*8), w96 => Pw(38)( 96*8-1 downto  95*8), 
w97 => Pw(38)( 97*8-1 downto  96*8), w98 => Pw(38)( 98*8-1 downto  97*8), w99 => Pw(38)( 99*8-1 downto  98*8), w100=> Pw(38)(100*8-1 downto  99*8), w101=> Pw(38)(101*8-1 downto 100*8), w102=> Pw(38)(102*8-1 downto 101*8), w103=> Pw(38)(103*8-1 downto 102*8), w104=> Pw(38)(104*8-1 downto 103*8), 
w105=> Pw(38)(105*8-1 downto 104*8), w106=> Pw(38)(106*8-1 downto 105*8), w107=> Pw(38)(107*8-1 downto 106*8), w108=> Pw(38)(108*8-1 downto 107*8), w109=> Pw(38)(109*8-1 downto 108*8), w110=> Pw(38)(110*8-1 downto 109*8), w111=> Pw(38)(111*8-1 downto 110*8), w112=> Pw(38)(112*8-1 downto 111*8), 
w113=> Pw(38)(113*8-1 downto 112*8), w114=> Pw(38)(114*8-1 downto 113*8), w115=> Pw(38)(115*8-1 downto 114*8), w116=> Pw(38)(116*8-1 downto 115*8), w117=> Pw(38)(117*8-1 downto 116*8), w118=> Pw(38)(118*8-1 downto 117*8), w119=> Pw(38)(119*8-1 downto 118*8), w120=> Pw(38)(120*8-1 downto 119*8), 
w121=> Pw(38)(121*8-1 downto 120*8), w122=> Pw(38)(122*8-1 downto 121*8), w123=> Pw(38)(123*8-1 downto 122*8), w124=> Pw(38)(124*8-1 downto 123*8), w125=> Pw(38)(125*8-1 downto 124*8), w126=> Pw(38)(126*8-1 downto 125*8), w127=> Pw(38)(127*8-1 downto 126*8), w128=> Pw(38)(128*8-1 downto 127*8), 

           d_out   => pca_d38_out   ,
           en_out  => open  ,
           sof_out => open );

  
  PCA128_39_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(39)(     7 downto    0), w02 => Pw(39)( 2*8-1 downto    8), w03 => Pw(39)( 3*8-1 downto  2*8), w04 => Pw(39)( 4*8-1 downto  3*8), w05 => Pw(39)( 5*8-1 downto  4*8), w06 => Pw(39)( 6*8-1 downto  5*8), w07 => Pw(39)( 7*8-1 downto  6*8), w08 => Pw(39)( 8*8-1 downto  7*8),  
w09 => Pw(39)( 9*8-1 downto  8*8), w10 => Pw(39)(10*8-1 downto  9*8), w11 => Pw(39)(11*8-1 downto 10*8), w12 => Pw(39)(12*8-1 downto 11*8), w13 => Pw(39)(13*8-1 downto 12*8), w14 => Pw(39)(14*8-1 downto 13*8), w15 => Pw(39)(15*8-1 downto 14*8), w16 => Pw(39)(16*8-1 downto 15*8),  
w17 => Pw(39)(17*8-1 downto 16*8), w18 => Pw(39)(18*8-1 downto 17*8), w19 => Pw(39)(19*8-1 downto 18*8), w20 => Pw(39)(20*8-1 downto 19*8), w21 => Pw(39)(21*8-1 downto 20*8), w22 => Pw(39)(22*8-1 downto 21*8), w23 => Pw(39)(23*8-1 downto 22*8), w24 => Pw(39)(24*8-1 downto 23*8),  
w25 => Pw(39)(25*8-1 downto 24*8), w26 => Pw(39)(26*8-1 downto 25*8), w27 => Pw(39)(27*8-1 downto 26*8), w28 => Pw(39)(28*8-1 downto 27*8), w29 => Pw(39)(29*8-1 downto 28*8), w30 => Pw(39)(30*8-1 downto 29*8), w31 => Pw(39)(31*8-1 downto 30*8), w32 => Pw(39)(32*8-1 downto 31*8),  
w33 => Pw(39)(33*8-1 downto 32*8), w34 => Pw(39)(34*8-1 downto 33*8), w35 => Pw(39)(35*8-1 downto 34*8), w36 => Pw(39)(36*8-1 downto 35*8), w37 => Pw(39)(37*8-1 downto 36*8), w38 => Pw(39)(38*8-1 downto 37*8), w39 => Pw(39)(39*8-1 downto 38*8), w40 => Pw(39)(40*8-1 downto 39*8),  
w41 => Pw(39)(41*8-1 downto 40*8), w42 => Pw(39)(42*8-1 downto 41*8), w43 => Pw(39)(43*8-1 downto 42*8), w44 => Pw(39)(44*8-1 downto 43*8), w45 => Pw(39)(45*8-1 downto 44*8), w46 => Pw(39)(46*8-1 downto 45*8), w47 => Pw(39)(47*8-1 downto 46*8), w48 => Pw(39)(48*8-1 downto 47*8),  
w49 => Pw(39)(49*8-1 downto 48*8), w50 => Pw(39)(50*8-1 downto 49*8), w51 => Pw(39)(51*8-1 downto 50*8), w52 => Pw(39)(52*8-1 downto 51*8), w53 => Pw(39)(53*8-1 downto 52*8), w54 => Pw(39)(54*8-1 downto 53*8), w55 => Pw(39)(55*8-1 downto 54*8), w56 => Pw(39)(56*8-1 downto 55*8),  
w57 => Pw(39)(57*8-1 downto 56*8), w58 => Pw(39)(58*8-1 downto 57*8), w59 => Pw(39)(59*8-1 downto 58*8), w60 => Pw(39)(60*8-1 downto 59*8), w61 => Pw(39)(61*8-1 downto 60*8), w62 => Pw(39)(62*8-1 downto 61*8), w63 => Pw(39)(63*8-1 downto 62*8), w64 => Pw(39)(64*8-1 downto 63*8), 
w65 => Pw(39)( 65*8-1 downto  64*8), w66 => Pw(39)( 66*8-1 downto  65*8), w67 => Pw(39)( 67*8-1 downto  66*8), w68 => Pw(39)( 68*8-1 downto  67*8), w69 => Pw(39)( 69*8-1 downto  68*8), w70 => Pw(39)( 70*8-1 downto  69*8), w71 => Pw(39)( 71*8-1 downto  70*8), w72 => Pw(39)( 72*8-1 downto  71*8), 
w73 => Pw(39)( 73*8-1 downto  72*8), w74 => Pw(39)( 74*8-1 downto  73*8), w75 => Pw(39)( 75*8-1 downto  74*8), w76 => Pw(39)( 76*8-1 downto  75*8), w77 => Pw(39)( 77*8-1 downto  76*8), w78 => Pw(39)( 78*8-1 downto  77*8), w79 => Pw(39)( 79*8-1 downto  78*8), w80 => Pw(39)( 80*8-1 downto  79*8), 
w81 => Pw(39)( 81*8-1 downto  80*8), w82 => Pw(39)( 82*8-1 downto  81*8), w83 => Pw(39)( 83*8-1 downto  82*8), w84 => Pw(39)( 84*8-1 downto  83*8), w85 => Pw(39)( 85*8-1 downto  84*8), w86 => Pw(39)( 86*8-1 downto  85*8), w87 => Pw(39)( 87*8-1 downto  86*8), w88 => Pw(39)( 88*8-1 downto  87*8), 
w89 => Pw(39)( 89*8-1 downto  88*8), w90 => Pw(39)( 90*8-1 downto  89*8), w91 => Pw(39)( 91*8-1 downto  90*8), w92 => Pw(39)( 92*8-1 downto  91*8), w93 => Pw(39)( 93*8-1 downto  92*8), w94 => Pw(39)( 94*8-1 downto  93*8), w95 => Pw(39)( 95*8-1 downto  94*8), w96 => Pw(39)( 96*8-1 downto  95*8), 
w97 => Pw(39)( 97*8-1 downto  96*8), w98 => Pw(39)( 98*8-1 downto  97*8), w99 => Pw(39)( 99*8-1 downto  98*8), w100=> Pw(39)(100*8-1 downto  99*8), w101=> Pw(39)(101*8-1 downto 100*8), w102=> Pw(39)(102*8-1 downto 101*8), w103=> Pw(39)(103*8-1 downto 102*8), w104=> Pw(39)(104*8-1 downto 103*8), 
w105=> Pw(39)(105*8-1 downto 104*8), w106=> Pw(39)(106*8-1 downto 105*8), w107=> Pw(39)(107*8-1 downto 106*8), w108=> Pw(39)(108*8-1 downto 107*8), w109=> Pw(39)(109*8-1 downto 108*8), w110=> Pw(39)(110*8-1 downto 109*8), w111=> Pw(39)(111*8-1 downto 110*8), w112=> Pw(39)(112*8-1 downto 111*8), 
w113=> Pw(39)(113*8-1 downto 112*8), w114=> Pw(39)(114*8-1 downto 113*8), w115=> Pw(39)(115*8-1 downto 114*8), w116=> Pw(39)(116*8-1 downto 115*8), w117=> Pw(39)(117*8-1 downto 116*8), w118=> Pw(39)(118*8-1 downto 117*8), w119=> Pw(39)(119*8-1 downto 118*8), w120=> Pw(39)(120*8-1 downto 119*8), 
w121=> Pw(39)(121*8-1 downto 120*8), w122=> Pw(39)(122*8-1 downto 121*8), w123=> Pw(39)(123*8-1 downto 122*8), w124=> Pw(39)(124*8-1 downto 123*8), w125=> Pw(39)(125*8-1 downto 124*8), w126=> Pw(39)(126*8-1 downto 125*8), w127=> Pw(39)(127*8-1 downto 126*8), w128=> Pw(39)(128*8-1 downto 127*8), 

           d_out   => pca_d39_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_40_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out, 

w01 => Pw(40)(     7 downto    0), w02 => Pw(40)( 2*8-1 downto    8), w03 => Pw(40)( 3*8-1 downto  2*8), w04 => Pw(40)( 4*8-1 downto  3*8), w05 => Pw(40)( 5*8-1 downto  4*8), w06 => Pw(40)( 6*8-1 downto  5*8), w07 => Pw(40)( 7*8-1 downto  6*8), w08 => Pw(40)( 8*8-1 downto  7*8),  
w09 => Pw(40)( 9*8-1 downto  8*8), w10 => Pw(40)(10*8-1 downto  9*8), w11 => Pw(40)(11*8-1 downto 10*8), w12 => Pw(40)(12*8-1 downto 11*8), w13 => Pw(40)(13*8-1 downto 12*8), w14 => Pw(40)(14*8-1 downto 13*8), w15 => Pw(40)(15*8-1 downto 14*8), w16 => Pw(40)(16*8-1 downto 15*8),  
w17 => Pw(40)(17*8-1 downto 16*8), w18 => Pw(40)(18*8-1 downto 17*8), w19 => Pw(40)(19*8-1 downto 18*8), w20 => Pw(40)(20*8-1 downto 19*8), w21 => Pw(40)(21*8-1 downto 20*8), w22 => Pw(40)(22*8-1 downto 21*8), w23 => Pw(40)(23*8-1 downto 22*8), w24 => Pw(40)(24*8-1 downto 23*8),  
w25 => Pw(40)(25*8-1 downto 24*8), w26 => Pw(40)(26*8-1 downto 25*8), w27 => Pw(40)(27*8-1 downto 26*8), w28 => Pw(40)(28*8-1 downto 27*8), w29 => Pw(40)(29*8-1 downto 28*8), w30 => Pw(40)(30*8-1 downto 29*8), w31 => Pw(40)(31*8-1 downto 30*8), w32 => Pw(40)(32*8-1 downto 31*8),  
w33 => Pw(40)(33*8-1 downto 32*8), w34 => Pw(40)(34*8-1 downto 33*8), w35 => Pw(40)(35*8-1 downto 34*8), w36 => Pw(40)(36*8-1 downto 35*8), w37 => Pw(40)(37*8-1 downto 36*8), w38 => Pw(40)(38*8-1 downto 37*8), w39 => Pw(40)(39*8-1 downto 38*8), w40 => Pw(40)(40*8-1 downto 39*8),  
w41 => Pw(40)(41*8-1 downto 40*8), w42 => Pw(40)(42*8-1 downto 41*8), w43 => Pw(40)(43*8-1 downto 42*8), w44 => Pw(40)(44*8-1 downto 43*8), w45 => Pw(40)(45*8-1 downto 44*8), w46 => Pw(40)(46*8-1 downto 45*8), w47 => Pw(40)(47*8-1 downto 46*8), w48 => Pw(40)(48*8-1 downto 47*8),  
w49 => Pw(40)(49*8-1 downto 48*8), w50 => Pw(40)(50*8-1 downto 49*8), w51 => Pw(40)(51*8-1 downto 50*8), w52 => Pw(40)(52*8-1 downto 51*8), w53 => Pw(40)(53*8-1 downto 52*8), w54 => Pw(40)(54*8-1 downto 53*8), w55 => Pw(40)(55*8-1 downto 54*8), w56 => Pw(40)(56*8-1 downto 55*8),  
w57 => Pw(40)(57*8-1 downto 56*8), w58 => Pw(40)(58*8-1 downto 57*8), w59 => Pw(40)(59*8-1 downto 58*8), w60 => Pw(40)(60*8-1 downto 59*8), w61 => Pw(40)(61*8-1 downto 60*8), w62 => Pw(40)(62*8-1 downto 61*8), w63 => Pw(40)(63*8-1 downto 62*8), w64 => Pw(40)(64*8-1 downto 63*8), 
w65 => Pw(40)( 65*8-1 downto  64*8), w66 => Pw(40)( 66*8-1 downto  65*8), w67 => Pw(40)( 67*8-1 downto  66*8), w68 => Pw(40)( 68*8-1 downto  67*8), w69 => Pw(40)( 69*8-1 downto  68*8), w70 => Pw(40)( 70*8-1 downto  69*8), w71 => Pw(40)( 71*8-1 downto  70*8), w72 => Pw(40)( 72*8-1 downto  71*8), 
w73 => Pw(40)( 73*8-1 downto  72*8), w74 => Pw(40)( 74*8-1 downto  73*8), w75 => Pw(40)( 75*8-1 downto  74*8), w76 => Pw(40)( 76*8-1 downto  75*8), w77 => Pw(40)( 77*8-1 downto  76*8), w78 => Pw(40)( 78*8-1 downto  77*8), w79 => Pw(40)( 79*8-1 downto  78*8), w80 => Pw(40)( 80*8-1 downto  79*8), 
w81 => Pw(40)( 81*8-1 downto  80*8), w82 => Pw(40)( 82*8-1 downto  81*8), w83 => Pw(40)( 83*8-1 downto  82*8), w84 => Pw(40)( 84*8-1 downto  83*8), w85 => Pw(40)( 85*8-1 downto  84*8), w86 => Pw(40)( 86*8-1 downto  85*8), w87 => Pw(40)( 87*8-1 downto  86*8), w88 => Pw(40)( 88*8-1 downto  87*8), 
w89 => Pw(40)( 89*8-1 downto  88*8), w90 => Pw(40)( 90*8-1 downto  89*8), w91 => Pw(40)( 91*8-1 downto  90*8), w92 => Pw(40)( 92*8-1 downto  91*8), w93 => Pw(40)( 93*8-1 downto  92*8), w94 => Pw(40)( 94*8-1 downto  93*8), w95 => Pw(40)( 95*8-1 downto  94*8), w96 => Pw(40)( 96*8-1 downto  95*8), 
w97 => Pw(40)( 97*8-1 downto  96*8), w98 => Pw(40)( 98*8-1 downto  97*8), w99 => Pw(40)( 99*8-1 downto  98*8), w100=> Pw(40)(100*8-1 downto  99*8), w101=> Pw(40)(101*8-1 downto 100*8), w102=> Pw(40)(102*8-1 downto 101*8), w103=> Pw(40)(103*8-1 downto 102*8), w104=> Pw(40)(104*8-1 downto 103*8), 
w105=> Pw(40)(105*8-1 downto 104*8), w106=> Pw(40)(106*8-1 downto 105*8), w107=> Pw(40)(107*8-1 downto 106*8), w108=> Pw(40)(108*8-1 downto 107*8), w109=> Pw(40)(109*8-1 downto 108*8), w110=> Pw(40)(110*8-1 downto 109*8), w111=> Pw(40)(111*8-1 downto 110*8), w112=> Pw(40)(112*8-1 downto 111*8), 
w113=> Pw(40)(113*8-1 downto 112*8), w114=> Pw(40)(114*8-1 downto 113*8), w115=> Pw(40)(115*8-1 downto 114*8), w116=> Pw(40)(116*8-1 downto 115*8), w117=> Pw(40)(117*8-1 downto 116*8), w118=> Pw(40)(118*8-1 downto 117*8), w119=> Pw(40)(119*8-1 downto 118*8), w120=> Pw(40)(120*8-1 downto 119*8), 
w121=> Pw(40)(121*8-1 downto 120*8), w122=> Pw(40)(122*8-1 downto 121*8), w123=> Pw(40)(123*8-1 downto 122*8), w124=> Pw(40)(124*8-1 downto 123*8), w125=> Pw(40)(125*8-1 downto 124*8), w126=> Pw(40)(126*8-1 downto 125*8), w127=> Pw(40)(127*8-1 downto 126*8), w128=> Pw(40)(128*8-1 downto 127*8), 

           d_out   => pca_d40_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_41_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(41)(     7 downto    0), w02 => Pw(41)( 2*8-1 downto    8), w03 => Pw(41)( 3*8-1 downto  2*8), w04 => Pw(41)( 4*8-1 downto  3*8), w05 => Pw(41)( 5*8-1 downto  4*8), w06 => Pw(41)( 6*8-1 downto  5*8), w07 => Pw(41)( 7*8-1 downto  6*8), w08 => Pw(41)( 8*8-1 downto  7*8),  
w09 => Pw(41)( 9*8-1 downto  8*8), w10 => Pw(41)(10*8-1 downto  9*8), w11 => Pw(41)(11*8-1 downto 10*8), w12 => Pw(41)(12*8-1 downto 11*8), w13 => Pw(41)(13*8-1 downto 12*8), w14 => Pw(41)(14*8-1 downto 13*8), w15 => Pw(41)(15*8-1 downto 14*8), w16 => Pw(41)(16*8-1 downto 15*8),  
w17 => Pw(41)(17*8-1 downto 16*8), w18 => Pw(41)(18*8-1 downto 17*8), w19 => Pw(41)(19*8-1 downto 18*8), w20 => Pw(41)(20*8-1 downto 19*8), w21 => Pw(41)(21*8-1 downto 20*8), w22 => Pw(41)(22*8-1 downto 21*8), w23 => Pw(41)(23*8-1 downto 22*8), w24 => Pw(41)(24*8-1 downto 23*8),  
w25 => Pw(41)(25*8-1 downto 24*8), w26 => Pw(41)(26*8-1 downto 25*8), w27 => Pw(41)(27*8-1 downto 26*8), w28 => Pw(41)(28*8-1 downto 27*8), w29 => Pw(41)(29*8-1 downto 28*8), w30 => Pw(41)(30*8-1 downto 29*8), w31 => Pw(41)(31*8-1 downto 30*8), w32 => Pw(41)(32*8-1 downto 31*8),  
w33 => Pw(41)(33*8-1 downto 32*8), w34 => Pw(41)(34*8-1 downto 33*8), w35 => Pw(41)(35*8-1 downto 34*8), w36 => Pw(41)(36*8-1 downto 35*8), w37 => Pw(41)(37*8-1 downto 36*8), w38 => Pw(41)(38*8-1 downto 37*8), w39 => Pw(41)(39*8-1 downto 38*8), w40 => Pw(41)(40*8-1 downto 39*8),  
w41 => Pw(41)(41*8-1 downto 40*8), w42 => Pw(41)(42*8-1 downto 41*8), w43 => Pw(41)(43*8-1 downto 42*8), w44 => Pw(41)(44*8-1 downto 43*8), w45 => Pw(41)(45*8-1 downto 44*8), w46 => Pw(41)(46*8-1 downto 45*8), w47 => Pw(41)(47*8-1 downto 46*8), w48 => Pw(41)(48*8-1 downto 47*8),  
w49 => Pw(41)(49*8-1 downto 48*8), w50 => Pw(41)(50*8-1 downto 49*8), w51 => Pw(41)(51*8-1 downto 50*8), w52 => Pw(41)(52*8-1 downto 51*8), w53 => Pw(41)(53*8-1 downto 52*8), w54 => Pw(41)(54*8-1 downto 53*8), w55 => Pw(41)(55*8-1 downto 54*8), w56 => Pw(41)(56*8-1 downto 55*8),  
w57 => Pw(41)(57*8-1 downto 56*8), w58 => Pw(41)(58*8-1 downto 57*8), w59 => Pw(41)(59*8-1 downto 58*8), w60 => Pw(41)(60*8-1 downto 59*8), w61 => Pw(41)(61*8-1 downto 60*8), w62 => Pw(41)(62*8-1 downto 61*8), w63 => Pw(41)(63*8-1 downto 62*8), w64 => Pw(41)(64*8-1 downto 63*8), 
w65 => Pw(41)( 65*8-1 downto  64*8), w66 => Pw(41)( 66*8-1 downto  65*8), w67 => Pw(41)( 67*8-1 downto  66*8), w68 => Pw(41)( 68*8-1 downto  67*8), w69 => Pw(41)( 69*8-1 downto  68*8), w70 => Pw(41)( 70*8-1 downto  69*8), w71 => Pw(41)( 71*8-1 downto  70*8), w72 => Pw(41)( 72*8-1 downto  71*8), 
w73 => Pw(41)( 73*8-1 downto  72*8), w74 => Pw(41)( 74*8-1 downto  73*8), w75 => Pw(41)( 75*8-1 downto  74*8), w76 => Pw(41)( 76*8-1 downto  75*8), w77 => Pw(41)( 77*8-1 downto  76*8), w78 => Pw(41)( 78*8-1 downto  77*8), w79 => Pw(41)( 79*8-1 downto  78*8), w80 => Pw(41)( 80*8-1 downto  79*8), 
w81 => Pw(41)( 81*8-1 downto  80*8), w82 => Pw(41)( 82*8-1 downto  81*8), w83 => Pw(41)( 83*8-1 downto  82*8), w84 => Pw(41)( 84*8-1 downto  83*8), w85 => Pw(41)( 85*8-1 downto  84*8), w86 => Pw(41)( 86*8-1 downto  85*8), w87 => Pw(41)( 87*8-1 downto  86*8), w88 => Pw(41)( 88*8-1 downto  87*8), 
w89 => Pw(41)( 89*8-1 downto  88*8), w90 => Pw(41)( 90*8-1 downto  89*8), w91 => Pw(41)( 91*8-1 downto  90*8), w92 => Pw(41)( 92*8-1 downto  91*8), w93 => Pw(41)( 93*8-1 downto  92*8), w94 => Pw(41)( 94*8-1 downto  93*8), w95 => Pw(41)( 95*8-1 downto  94*8), w96 => Pw(41)( 96*8-1 downto  95*8), 
w97 => Pw(41)( 97*8-1 downto  96*8), w98 => Pw(41)( 98*8-1 downto  97*8), w99 => Pw(41)( 99*8-1 downto  98*8), w100=> Pw(41)(100*8-1 downto  99*8), w101=> Pw(41)(101*8-1 downto 100*8), w102=> Pw(41)(102*8-1 downto 101*8), w103=> Pw(41)(103*8-1 downto 102*8), w104=> Pw(41)(104*8-1 downto 103*8), 
w105=> Pw(41)(105*8-1 downto 104*8), w106=> Pw(41)(106*8-1 downto 105*8), w107=> Pw(41)(107*8-1 downto 106*8), w108=> Pw(41)(108*8-1 downto 107*8), w109=> Pw(41)(109*8-1 downto 108*8), w110=> Pw(41)(110*8-1 downto 109*8), w111=> Pw(41)(111*8-1 downto 110*8), w112=> Pw(41)(112*8-1 downto 111*8), 
w113=> Pw(41)(113*8-1 downto 112*8), w114=> Pw(41)(114*8-1 downto 113*8), w115=> Pw(41)(115*8-1 downto 114*8), w116=> Pw(41)(116*8-1 downto 115*8), w117=> Pw(41)(117*8-1 downto 116*8), w118=> Pw(41)(118*8-1 downto 117*8), w119=> Pw(41)(119*8-1 downto 118*8), w120=> Pw(41)(120*8-1 downto 119*8), 
w121=> Pw(41)(121*8-1 downto 120*8), w122=> Pw(41)(122*8-1 downto 121*8), w123=> Pw(41)(123*8-1 downto 122*8), w124=> Pw(41)(124*8-1 downto 123*8), w125=> Pw(41)(125*8-1 downto 124*8), w126=> Pw(41)(126*8-1 downto 125*8), w127=> Pw(41)(127*8-1 downto 126*8), w128=> Pw(41)(128*8-1 downto 127*8), 

           d_out   => pca_d41_out   ,
           en_out  => open  ,
           sof_out => open );


PCA128_42_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(42)(     7 downto    0), w02 => Pw(42)( 2*8-1 downto    8), w03 => Pw(42)( 3*8-1 downto  2*8), w04 => Pw(42)( 4*8-1 downto  3*8), w05 => Pw(42)( 5*8-1 downto  4*8), w06 => Pw(42)( 6*8-1 downto  5*8), w07 => Pw(42)( 7*8-1 downto  6*8), w08 => Pw(42)( 8*8-1 downto  7*8),  
w09 => Pw(42)( 9*8-1 downto  8*8), w10 => Pw(42)(10*8-1 downto  9*8), w11 => Pw(42)(11*8-1 downto 10*8), w12 => Pw(42)(12*8-1 downto 11*8), w13 => Pw(42)(13*8-1 downto 12*8), w14 => Pw(42)(14*8-1 downto 13*8), w15 => Pw(42)(15*8-1 downto 14*8), w16 => Pw(42)(16*8-1 downto 15*8),  
w17 => Pw(42)(17*8-1 downto 16*8), w18 => Pw(42)(18*8-1 downto 17*8), w19 => Pw(42)(19*8-1 downto 18*8), w20 => Pw(42)(20*8-1 downto 19*8), w21 => Pw(42)(21*8-1 downto 20*8), w22 => Pw(42)(22*8-1 downto 21*8), w23 => Pw(42)(23*8-1 downto 22*8), w24 => Pw(42)(24*8-1 downto 23*8),  
w25 => Pw(42)(25*8-1 downto 24*8), w26 => Pw(42)(26*8-1 downto 25*8), w27 => Pw(42)(27*8-1 downto 26*8), w28 => Pw(42)(28*8-1 downto 27*8), w29 => Pw(42)(29*8-1 downto 28*8), w30 => Pw(42)(30*8-1 downto 29*8), w31 => Pw(42)(31*8-1 downto 30*8), w32 => Pw(42)(32*8-1 downto 31*8),  
w33 => Pw(42)(33*8-1 downto 32*8), w34 => Pw(42)(34*8-1 downto 33*8), w35 => Pw(42)(35*8-1 downto 34*8), w36 => Pw(42)(36*8-1 downto 35*8), w37 => Pw(42)(37*8-1 downto 36*8), w38 => Pw(42)(38*8-1 downto 37*8), w39 => Pw(42)(39*8-1 downto 38*8), w40 => Pw(42)(40*8-1 downto 39*8),  
w41 => Pw(42)(41*8-1 downto 40*8), w42 => Pw(42)(42*8-1 downto 41*8), w43 => Pw(42)(43*8-1 downto 42*8), w44 => Pw(42)(44*8-1 downto 43*8), w45 => Pw(42)(45*8-1 downto 44*8), w46 => Pw(42)(46*8-1 downto 45*8), w47 => Pw(42)(47*8-1 downto 46*8), w48 => Pw(42)(48*8-1 downto 47*8),  
w49 => Pw(42)(49*8-1 downto 48*8), w50 => Pw(42)(50*8-1 downto 49*8), w51 => Pw(42)(51*8-1 downto 50*8), w52 => Pw(42)(52*8-1 downto 51*8), w53 => Pw(42)(53*8-1 downto 52*8), w54 => Pw(42)(54*8-1 downto 53*8), w55 => Pw(42)(55*8-1 downto 54*8), w56 => Pw(42)(56*8-1 downto 55*8),  
w57 => Pw(42)(57*8-1 downto 56*8), w58 => Pw(42)(58*8-1 downto 57*8), w59 => Pw(42)(59*8-1 downto 58*8), w60 => Pw(42)(60*8-1 downto 59*8), w61 => Pw(42)(61*8-1 downto 60*8), w62 => Pw(42)(62*8-1 downto 61*8), w63 => Pw(42)(63*8-1 downto 62*8), w64 => Pw(42)(64*8-1 downto 63*8), 
w65 => Pw(42)( 65*8-1 downto  64*8), w66 => Pw(42)( 66*8-1 downto  65*8), w67 => Pw(42)( 67*8-1 downto  66*8), w68 => Pw(42)( 68*8-1 downto  67*8), w69 => Pw(42)( 69*8-1 downto  68*8), w70 => Pw(42)( 70*8-1 downto  69*8), w71 => Pw(42)( 71*8-1 downto  70*8), w72 => Pw(42)( 72*8-1 downto  71*8), 
w73 => Pw(42)( 73*8-1 downto  72*8), w74 => Pw(42)( 74*8-1 downto  73*8), w75 => Pw(42)( 75*8-1 downto  74*8), w76 => Pw(42)( 76*8-1 downto  75*8), w77 => Pw(42)( 77*8-1 downto  76*8), w78 => Pw(42)( 78*8-1 downto  77*8), w79 => Pw(42)( 79*8-1 downto  78*8), w80 => Pw(42)( 80*8-1 downto  79*8), 
w81 => Pw(42)( 81*8-1 downto  80*8), w82 => Pw(42)( 82*8-1 downto  81*8), w83 => Pw(42)( 83*8-1 downto  82*8), w84 => Pw(42)( 84*8-1 downto  83*8), w85 => Pw(42)( 85*8-1 downto  84*8), w86 => Pw(42)( 86*8-1 downto  85*8), w87 => Pw(42)( 87*8-1 downto  86*8), w88 => Pw(42)( 88*8-1 downto  87*8), 
w89 => Pw(42)( 89*8-1 downto  88*8), w90 => Pw(42)( 90*8-1 downto  89*8), w91 => Pw(42)( 91*8-1 downto  90*8), w92 => Pw(42)( 92*8-1 downto  91*8), w93 => Pw(42)( 93*8-1 downto  92*8), w94 => Pw(42)( 94*8-1 downto  93*8), w95 => Pw(42)( 95*8-1 downto  94*8), w96 => Pw(42)( 96*8-1 downto  95*8), 
w97 => Pw(42)( 97*8-1 downto  96*8), w98 => Pw(42)( 98*8-1 downto  97*8), w99 => Pw(42)( 99*8-1 downto  98*8), w100=> Pw(42)(100*8-1 downto  99*8), w101=> Pw(42)(101*8-1 downto 100*8), w102=> Pw(42)(102*8-1 downto 101*8), w103=> Pw(42)(103*8-1 downto 102*8), w104=> Pw(42)(104*8-1 downto 103*8), 
w105=> Pw(42)(105*8-1 downto 104*8), w106=> Pw(42)(106*8-1 downto 105*8), w107=> Pw(42)(107*8-1 downto 106*8), w108=> Pw(42)(108*8-1 downto 107*8), w109=> Pw(42)(109*8-1 downto 108*8), w110=> Pw(42)(110*8-1 downto 109*8), w111=> Pw(42)(111*8-1 downto 110*8), w112=> Pw(42)(112*8-1 downto 111*8), 
w113=> Pw(42)(113*8-1 downto 112*8), w114=> Pw(42)(114*8-1 downto 113*8), w115=> Pw(42)(115*8-1 downto 114*8), w116=> Pw(42)(116*8-1 downto 115*8), w117=> Pw(42)(117*8-1 downto 116*8), w118=> Pw(42)(118*8-1 downto 117*8), w119=> Pw(42)(119*8-1 downto 118*8), w120=> Pw(42)(120*8-1 downto 119*8), 
w121=> Pw(42)(121*8-1 downto 120*8), w122=> Pw(42)(122*8-1 downto 121*8), w123=> Pw(42)(123*8-1 downto 122*8), w124=> Pw(42)(124*8-1 downto 123*8), w125=> Pw(42)(125*8-1 downto 124*8), w126=> Pw(42)(126*8-1 downto 125*8), w127=> Pw(42)(127*8-1 downto 126*8), w128=> Pw(42)(128*8-1 downto 127*8), 

           d_out   => pca_d42_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_43_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(43)(     7 downto    0), w02 => Pw(43)( 2*8-1 downto    8), w03 => Pw(43)( 3*8-1 downto  2*8), w04 => Pw(43)( 4*8-1 downto  3*8), w05 => Pw(43)( 5*8-1 downto  4*8), w06 => Pw(43)( 6*8-1 downto  5*8), w07 => Pw(43)( 7*8-1 downto  6*8), w08 => Pw(43)( 8*8-1 downto  7*8),  
w09 => Pw(43)( 9*8-1 downto  8*8), w10 => Pw(43)(10*8-1 downto  9*8), w11 => Pw(43)(11*8-1 downto 10*8), w12 => Pw(43)(12*8-1 downto 11*8), w13 => Pw(43)(13*8-1 downto 12*8), w14 => Pw(43)(14*8-1 downto 13*8), w15 => Pw(43)(15*8-1 downto 14*8), w16 => Pw(43)(16*8-1 downto 15*8),  
w17 => Pw(43)(17*8-1 downto 16*8), w18 => Pw(43)(18*8-1 downto 17*8), w19 => Pw(43)(19*8-1 downto 18*8), w20 => Pw(43)(20*8-1 downto 19*8), w21 => Pw(43)(21*8-1 downto 20*8), w22 => Pw(43)(22*8-1 downto 21*8), w23 => Pw(43)(23*8-1 downto 22*8), w24 => Pw(43)(24*8-1 downto 23*8),  
w25 => Pw(43)(25*8-1 downto 24*8), w26 => Pw(43)(26*8-1 downto 25*8), w27 => Pw(43)(27*8-1 downto 26*8), w28 => Pw(43)(28*8-1 downto 27*8), w29 => Pw(43)(29*8-1 downto 28*8), w30 => Pw(43)(30*8-1 downto 29*8), w31 => Pw(43)(31*8-1 downto 30*8), w32 => Pw(43)(32*8-1 downto 31*8),  
w33 => Pw(43)(33*8-1 downto 32*8), w34 => Pw(43)(34*8-1 downto 33*8), w35 => Pw(43)(35*8-1 downto 34*8), w36 => Pw(43)(36*8-1 downto 35*8), w37 => Pw(43)(37*8-1 downto 36*8), w38 => Pw(43)(38*8-1 downto 37*8), w39 => Pw(43)(39*8-1 downto 38*8), w40 => Pw(43)(40*8-1 downto 39*8),  
w41 => Pw(43)(41*8-1 downto 40*8), w42 => Pw(43)(42*8-1 downto 41*8), w43 => Pw(43)(43*8-1 downto 42*8), w44 => Pw(43)(44*8-1 downto 43*8), w45 => Pw(43)(45*8-1 downto 44*8), w46 => Pw(43)(46*8-1 downto 45*8), w47 => Pw(43)(47*8-1 downto 46*8), w48 => Pw(43)(48*8-1 downto 47*8),  
w49 => Pw(43)(49*8-1 downto 48*8), w50 => Pw(43)(50*8-1 downto 49*8), w51 => Pw(43)(51*8-1 downto 50*8), w52 => Pw(43)(52*8-1 downto 51*8), w53 => Pw(43)(53*8-1 downto 52*8), w54 => Pw(43)(54*8-1 downto 53*8), w55 => Pw(43)(55*8-1 downto 54*8), w56 => Pw(43)(56*8-1 downto 55*8),  
w57 => Pw(43)(57*8-1 downto 56*8), w58 => Pw(43)(58*8-1 downto 57*8), w59 => Pw(43)(59*8-1 downto 58*8), w60 => Pw(43)(60*8-1 downto 59*8), w61 => Pw(43)(61*8-1 downto 60*8), w62 => Pw(43)(62*8-1 downto 61*8), w63 => Pw(43)(63*8-1 downto 62*8), w64 => Pw(43)(64*8-1 downto 63*8), 
w65 => Pw(43)( 65*8-1 downto  64*8), w66 => Pw(43)( 66*8-1 downto  65*8), w67 => Pw(43)( 67*8-1 downto  66*8), w68 => Pw(43)( 68*8-1 downto  67*8), w69 => Pw(43)( 69*8-1 downto  68*8), w70 => Pw(43)( 70*8-1 downto  69*8), w71 => Pw(43)( 71*8-1 downto  70*8), w72 => Pw(43)( 72*8-1 downto  71*8), 
w73 => Pw(43)( 73*8-1 downto  72*8), w74 => Pw(43)( 74*8-1 downto  73*8), w75 => Pw(43)( 75*8-1 downto  74*8), w76 => Pw(43)( 76*8-1 downto  75*8), w77 => Pw(43)( 77*8-1 downto  76*8), w78 => Pw(43)( 78*8-1 downto  77*8), w79 => Pw(43)( 79*8-1 downto  78*8), w80 => Pw(43)( 80*8-1 downto  79*8), 
w81 => Pw(43)( 81*8-1 downto  80*8), w82 => Pw(43)( 82*8-1 downto  81*8), w83 => Pw(43)( 83*8-1 downto  82*8), w84 => Pw(43)( 84*8-1 downto  83*8), w85 => Pw(43)( 85*8-1 downto  84*8), w86 => Pw(43)( 86*8-1 downto  85*8), w87 => Pw(43)( 87*8-1 downto  86*8), w88 => Pw(43)( 88*8-1 downto  87*8), 
w89 => Pw(43)( 89*8-1 downto  88*8), w90 => Pw(43)( 90*8-1 downto  89*8), w91 => Pw(43)( 91*8-1 downto  90*8), w92 => Pw(43)( 92*8-1 downto  91*8), w93 => Pw(43)( 93*8-1 downto  92*8), w94 => Pw(43)( 94*8-1 downto  93*8), w95 => Pw(43)( 95*8-1 downto  94*8), w96 => Pw(43)( 96*8-1 downto  95*8), 
w97 => Pw(43)( 97*8-1 downto  96*8), w98 => Pw(43)( 98*8-1 downto  97*8), w99 => Pw(43)( 99*8-1 downto  98*8), w100=> Pw(43)(100*8-1 downto  99*8), w101=> Pw(43)(101*8-1 downto 100*8), w102=> Pw(43)(102*8-1 downto 101*8), w103=> Pw(43)(103*8-1 downto 102*8), w104=> Pw(43)(104*8-1 downto 103*8), 
w105=> Pw(43)(105*8-1 downto 104*8), w106=> Pw(43)(106*8-1 downto 105*8), w107=> Pw(43)(107*8-1 downto 106*8), w108=> Pw(43)(108*8-1 downto 107*8), w109=> Pw(43)(109*8-1 downto 108*8), w110=> Pw(43)(110*8-1 downto 109*8), w111=> Pw(43)(111*8-1 downto 110*8), w112=> Pw(43)(112*8-1 downto 111*8), 
w113=> Pw(43)(113*8-1 downto 112*8), w114=> Pw(43)(114*8-1 downto 113*8), w115=> Pw(43)(115*8-1 downto 114*8), w116=> Pw(43)(116*8-1 downto 115*8), w117=> Pw(43)(117*8-1 downto 116*8), w118=> Pw(43)(118*8-1 downto 117*8), w119=> Pw(43)(119*8-1 downto 118*8), w120=> Pw(43)(120*8-1 downto 119*8), 
w121=> Pw(43)(121*8-1 downto 120*8), w122=> Pw(43)(122*8-1 downto 121*8), w123=> Pw(43)(123*8-1 downto 122*8), w124=> Pw(43)(124*8-1 downto 123*8), w125=> Pw(43)(125*8-1 downto 124*8), w126=> Pw(43)(126*8-1 downto 125*8), w127=> Pw(43)(127*8-1 downto 126*8), w128=> Pw(43)(128*8-1 downto 127*8), 

           d_out   => pca_d43_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_44_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(44)(     7 downto    0), w02 => Pw(44)( 2*8-1 downto    8), w03 => Pw(44)( 3*8-1 downto  2*8), w04 => Pw(44)( 4*8-1 downto  3*8), w05 => Pw(44)( 5*8-1 downto  4*8), w06 => Pw(44)( 6*8-1 downto  5*8), w07 => Pw(44)( 7*8-1 downto  6*8), w08 => Pw(44)( 8*8-1 downto  7*8),  
w09 => Pw(44)( 9*8-1 downto  8*8), w10 => Pw(44)(10*8-1 downto  9*8), w11 => Pw(44)(11*8-1 downto 10*8), w12 => Pw(44)(12*8-1 downto 11*8), w13 => Pw(44)(13*8-1 downto 12*8), w14 => Pw(44)(14*8-1 downto 13*8), w15 => Pw(44)(15*8-1 downto 14*8), w16 => Pw(44)(16*8-1 downto 15*8),  
w17 => Pw(44)(17*8-1 downto 16*8), w18 => Pw(44)(18*8-1 downto 17*8), w19 => Pw(44)(19*8-1 downto 18*8), w20 => Pw(44)(20*8-1 downto 19*8), w21 => Pw(44)(21*8-1 downto 20*8), w22 => Pw(44)(22*8-1 downto 21*8), w23 => Pw(44)(23*8-1 downto 22*8), w24 => Pw(44)(24*8-1 downto 23*8),  
w25 => Pw(44)(25*8-1 downto 24*8), w26 => Pw(44)(26*8-1 downto 25*8), w27 => Pw(44)(27*8-1 downto 26*8), w28 => Pw(44)(28*8-1 downto 27*8), w29 => Pw(44)(29*8-1 downto 28*8), w30 => Pw(44)(30*8-1 downto 29*8), w31 => Pw(44)(31*8-1 downto 30*8), w32 => Pw(44)(32*8-1 downto 31*8),  
w33 => Pw(44)(33*8-1 downto 32*8), w34 => Pw(44)(34*8-1 downto 33*8), w35 => Pw(44)(35*8-1 downto 34*8), w36 => Pw(44)(36*8-1 downto 35*8), w37 => Pw(44)(37*8-1 downto 36*8), w38 => Pw(44)(38*8-1 downto 37*8), w39 => Pw(44)(39*8-1 downto 38*8), w40 => Pw(44)(40*8-1 downto 39*8),  
w41 => Pw(44)(41*8-1 downto 40*8), w42 => Pw(44)(42*8-1 downto 41*8), w43 => Pw(44)(43*8-1 downto 42*8), w44 => Pw(44)(44*8-1 downto 43*8), w45 => Pw(44)(45*8-1 downto 44*8), w46 => Pw(44)(46*8-1 downto 45*8), w47 => Pw(44)(47*8-1 downto 46*8), w48 => Pw(44)(48*8-1 downto 47*8),  
w49 => Pw(44)(49*8-1 downto 48*8), w50 => Pw(44)(50*8-1 downto 49*8), w51 => Pw(44)(51*8-1 downto 50*8), w52 => Pw(44)(52*8-1 downto 51*8), w53 => Pw(44)(53*8-1 downto 52*8), w54 => Pw(44)(54*8-1 downto 53*8), w55 => Pw(44)(55*8-1 downto 54*8), w56 => Pw(44)(56*8-1 downto 55*8),  
w57 => Pw(44)(57*8-1 downto 56*8), w58 => Pw(44)(58*8-1 downto 57*8), w59 => Pw(44)(59*8-1 downto 58*8), w60 => Pw(44)(60*8-1 downto 59*8), w61 => Pw(44)(61*8-1 downto 60*8), w62 => Pw(44)(62*8-1 downto 61*8), w63 => Pw(44)(63*8-1 downto 62*8), w64 => Pw(44)(64*8-1 downto 63*8), 
w65 => Pw(44)( 65*8-1 downto  64*8), w66 => Pw(44)( 66*8-1 downto  65*8), w67 => Pw(44)( 67*8-1 downto  66*8), w68 => Pw(44)( 68*8-1 downto  67*8), w69 => Pw(44)( 69*8-1 downto  68*8), w70 => Pw(44)( 70*8-1 downto  69*8), w71 => Pw(44)( 71*8-1 downto  70*8), w72 => Pw(44)( 72*8-1 downto  71*8), 
w73 => Pw(44)( 73*8-1 downto  72*8), w74 => Pw(44)( 74*8-1 downto  73*8), w75 => Pw(44)( 75*8-1 downto  74*8), w76 => Pw(44)( 76*8-1 downto  75*8), w77 => Pw(44)( 77*8-1 downto  76*8), w78 => Pw(44)( 78*8-1 downto  77*8), w79 => Pw(44)( 79*8-1 downto  78*8), w80 => Pw(44)( 80*8-1 downto  79*8), 
w81 => Pw(44)( 81*8-1 downto  80*8), w82 => Pw(44)( 82*8-1 downto  81*8), w83 => Pw(44)( 83*8-1 downto  82*8), w84 => Pw(44)( 84*8-1 downto  83*8), w85 => Pw(44)( 85*8-1 downto  84*8), w86 => Pw(44)( 86*8-1 downto  85*8), w87 => Pw(44)( 87*8-1 downto  86*8), w88 => Pw(44)( 88*8-1 downto  87*8), 
w89 => Pw(44)( 89*8-1 downto  88*8), w90 => Pw(44)( 90*8-1 downto  89*8), w91 => Pw(44)( 91*8-1 downto  90*8), w92 => Pw(44)( 92*8-1 downto  91*8), w93 => Pw(44)( 93*8-1 downto  92*8), w94 => Pw(44)( 94*8-1 downto  93*8), w95 => Pw(44)( 95*8-1 downto  94*8), w96 => Pw(44)( 96*8-1 downto  95*8), 
w97 => Pw(44)( 97*8-1 downto  96*8), w98 => Pw(44)( 98*8-1 downto  97*8), w99 => Pw(44)( 99*8-1 downto  98*8), w100=> Pw(44)(100*8-1 downto  99*8), w101=> Pw(44)(101*8-1 downto 100*8), w102=> Pw(44)(102*8-1 downto 101*8), w103=> Pw(44)(103*8-1 downto 102*8), w104=> Pw(44)(104*8-1 downto 103*8), 
w105=> Pw(44)(105*8-1 downto 104*8), w106=> Pw(44)(106*8-1 downto 105*8), w107=> Pw(44)(107*8-1 downto 106*8), w108=> Pw(44)(108*8-1 downto 107*8), w109=> Pw(44)(109*8-1 downto 108*8), w110=> Pw(44)(110*8-1 downto 109*8), w111=> Pw(44)(111*8-1 downto 110*8), w112=> Pw(44)(112*8-1 downto 111*8), 
w113=> Pw(44)(113*8-1 downto 112*8), w114=> Pw(44)(114*8-1 downto 113*8), w115=> Pw(44)(115*8-1 downto 114*8), w116=> Pw(44)(116*8-1 downto 115*8), w117=> Pw(44)(117*8-1 downto 116*8), w118=> Pw(44)(118*8-1 downto 117*8), w119=> Pw(44)(119*8-1 downto 118*8), w120=> Pw(44)(120*8-1 downto 119*8), 
w121=> Pw(44)(121*8-1 downto 120*8), w122=> Pw(44)(122*8-1 downto 121*8), w123=> Pw(44)(123*8-1 downto 122*8), w124=> Pw(44)(124*8-1 downto 123*8), w125=> Pw(44)(125*8-1 downto 124*8), w126=> Pw(44)(126*8-1 downto 125*8), w127=> Pw(44)(127*8-1 downto 126*8), w128=> Pw(44)(128*8-1 downto 127*8), 

           d_out   => pca_d44_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_45_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(45)(     7 downto    0), w02 => Pw(45)( 2*8-1 downto    8), w03 => Pw(45)( 3*8-1 downto  2*8), w04 => Pw(45)( 4*8-1 downto  3*8), w05 => Pw(45)( 5*8-1 downto  4*8), w06 => Pw(45)( 6*8-1 downto  5*8), w07 => Pw(45)( 7*8-1 downto  6*8), w08 => Pw(45)( 8*8-1 downto  7*8),  
w09 => Pw(45)( 9*8-1 downto  8*8), w10 => Pw(45)(10*8-1 downto  9*8), w11 => Pw(45)(11*8-1 downto 10*8), w12 => Pw(45)(12*8-1 downto 11*8), w13 => Pw(45)(13*8-1 downto 12*8), w14 => Pw(45)(14*8-1 downto 13*8), w15 => Pw(45)(15*8-1 downto 14*8), w16 => Pw(45)(16*8-1 downto 15*8),  
w17 => Pw(45)(17*8-1 downto 16*8), w18 => Pw(45)(18*8-1 downto 17*8), w19 => Pw(45)(19*8-1 downto 18*8), w20 => Pw(45)(20*8-1 downto 19*8), w21 => Pw(45)(21*8-1 downto 20*8), w22 => Pw(45)(22*8-1 downto 21*8), w23 => Pw(45)(23*8-1 downto 22*8), w24 => Pw(45)(24*8-1 downto 23*8),  
w25 => Pw(45)(25*8-1 downto 24*8), w26 => Pw(45)(26*8-1 downto 25*8), w27 => Pw(45)(27*8-1 downto 26*8), w28 => Pw(45)(28*8-1 downto 27*8), w29 => Pw(45)(29*8-1 downto 28*8), w30 => Pw(45)(30*8-1 downto 29*8), w31 => Pw(45)(31*8-1 downto 30*8), w32 => Pw(45)(32*8-1 downto 31*8),  
w33 => Pw(45)(33*8-1 downto 32*8), w34 => Pw(45)(34*8-1 downto 33*8), w35 => Pw(45)(35*8-1 downto 34*8), w36 => Pw(45)(36*8-1 downto 35*8), w37 => Pw(45)(37*8-1 downto 36*8), w38 => Pw(45)(38*8-1 downto 37*8), w39 => Pw(45)(39*8-1 downto 38*8), w40 => Pw(45)(40*8-1 downto 39*8),  
w41 => Pw(45)(41*8-1 downto 40*8), w42 => Pw(45)(42*8-1 downto 41*8), w43 => Pw(45)(43*8-1 downto 42*8), w44 => Pw(45)(44*8-1 downto 43*8), w45 => Pw(45)(45*8-1 downto 44*8), w46 => Pw(45)(46*8-1 downto 45*8), w47 => Pw(45)(47*8-1 downto 46*8), w48 => Pw(45)(48*8-1 downto 47*8),  
w49 => Pw(45)(49*8-1 downto 48*8), w50 => Pw(45)(50*8-1 downto 49*8), w51 => Pw(45)(51*8-1 downto 50*8), w52 => Pw(45)(52*8-1 downto 51*8), w53 => Pw(45)(53*8-1 downto 52*8), w54 => Pw(45)(54*8-1 downto 53*8), w55 => Pw(45)(55*8-1 downto 54*8), w56 => Pw(45)(56*8-1 downto 55*8),  
w57 => Pw(45)(57*8-1 downto 56*8), w58 => Pw(45)(58*8-1 downto 57*8), w59 => Pw(45)(59*8-1 downto 58*8), w60 => Pw(45)(60*8-1 downto 59*8), w61 => Pw(45)(61*8-1 downto 60*8), w62 => Pw(45)(62*8-1 downto 61*8), w63 => Pw(45)(63*8-1 downto 62*8), w64 => Pw(45)(64*8-1 downto 63*8), 
w65 => Pw(45)( 65*8-1 downto  64*8), w66 => Pw(45)( 66*8-1 downto  65*8), w67 => Pw(45)( 67*8-1 downto  66*8), w68 => Pw(45)( 68*8-1 downto  67*8), w69 => Pw(45)( 69*8-1 downto  68*8), w70 => Pw(45)( 70*8-1 downto  69*8), w71 => Pw(45)( 71*8-1 downto  70*8), w72 => Pw(45)( 72*8-1 downto  71*8), 
w73 => Pw(45)( 73*8-1 downto  72*8), w74 => Pw(45)( 74*8-1 downto  73*8), w75 => Pw(45)( 75*8-1 downto  74*8), w76 => Pw(45)( 76*8-1 downto  75*8), w77 => Pw(45)( 77*8-1 downto  76*8), w78 => Pw(45)( 78*8-1 downto  77*8), w79 => Pw(45)( 79*8-1 downto  78*8), w80 => Pw(45)( 80*8-1 downto  79*8), 
w81 => Pw(45)( 81*8-1 downto  80*8), w82 => Pw(45)( 82*8-1 downto  81*8), w83 => Pw(45)( 83*8-1 downto  82*8), w84 => Pw(45)( 84*8-1 downto  83*8), w85 => Pw(45)( 85*8-1 downto  84*8), w86 => Pw(45)( 86*8-1 downto  85*8), w87 => Pw(45)( 87*8-1 downto  86*8), w88 => Pw(45)( 88*8-1 downto  87*8), 
w89 => Pw(45)( 89*8-1 downto  88*8), w90 => Pw(45)( 90*8-1 downto  89*8), w91 => Pw(45)( 91*8-1 downto  90*8), w92 => Pw(45)( 92*8-1 downto  91*8), w93 => Pw(45)( 93*8-1 downto  92*8), w94 => Pw(45)( 94*8-1 downto  93*8), w95 => Pw(45)( 95*8-1 downto  94*8), w96 => Pw(45)( 96*8-1 downto  95*8), 
w97 => Pw(45)( 97*8-1 downto  96*8), w98 => Pw(45)( 98*8-1 downto  97*8), w99 => Pw(45)( 99*8-1 downto  98*8), w100=> Pw(45)(100*8-1 downto  99*8), w101=> Pw(45)(101*8-1 downto 100*8), w102=> Pw(45)(102*8-1 downto 101*8), w103=> Pw(45)(103*8-1 downto 102*8), w104=> Pw(45)(104*8-1 downto 103*8), 
w105=> Pw(45)(105*8-1 downto 104*8), w106=> Pw(45)(106*8-1 downto 105*8), w107=> Pw(45)(107*8-1 downto 106*8), w108=> Pw(45)(108*8-1 downto 107*8), w109=> Pw(45)(109*8-1 downto 108*8), w110=> Pw(45)(110*8-1 downto 109*8), w111=> Pw(45)(111*8-1 downto 110*8), w112=> Pw(45)(112*8-1 downto 111*8), 
w113=> Pw(45)(113*8-1 downto 112*8), w114=> Pw(45)(114*8-1 downto 113*8), w115=> Pw(45)(115*8-1 downto 114*8), w116=> Pw(45)(116*8-1 downto 115*8), w117=> Pw(45)(117*8-1 downto 116*8), w118=> Pw(45)(118*8-1 downto 117*8), w119=> Pw(45)(119*8-1 downto 118*8), w120=> Pw(45)(120*8-1 downto 119*8), 
w121=> Pw(45)(121*8-1 downto 120*8), w122=> Pw(45)(122*8-1 downto 121*8), w123=> Pw(45)(123*8-1 downto 122*8), w124=> Pw(45)(124*8-1 downto 123*8), w125=> Pw(45)(125*8-1 downto 124*8), w126=> Pw(45)(126*8-1 downto 125*8), w127=> Pw(45)(127*8-1 downto 126*8), w128=> Pw(45)(128*8-1 downto 127*8), 

           d_out   => pca_d45_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_46_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(46)(     7 downto    0), w02 => Pw(46)( 2*8-1 downto    8), w03 => Pw(46)( 3*8-1 downto  2*8), w04 => Pw(46)( 4*8-1 downto  3*8), w05 => Pw(46)( 5*8-1 downto  4*8), w06 => Pw(46)( 6*8-1 downto  5*8), w07 => Pw(46)( 7*8-1 downto  6*8), w08 => Pw(46)( 8*8-1 downto  7*8),  
w09 => Pw(46)( 9*8-1 downto  8*8), w10 => Pw(46)(10*8-1 downto  9*8), w11 => Pw(46)(11*8-1 downto 10*8), w12 => Pw(46)(12*8-1 downto 11*8), w13 => Pw(46)(13*8-1 downto 12*8), w14 => Pw(46)(14*8-1 downto 13*8), w15 => Pw(46)(15*8-1 downto 14*8), w16 => Pw(46)(16*8-1 downto 15*8),  
w17 => Pw(46)(17*8-1 downto 16*8), w18 => Pw(46)(18*8-1 downto 17*8), w19 => Pw(46)(19*8-1 downto 18*8), w20 => Pw(46)(20*8-1 downto 19*8), w21 => Pw(46)(21*8-1 downto 20*8), w22 => Pw(46)(22*8-1 downto 21*8), w23 => Pw(46)(23*8-1 downto 22*8), w24 => Pw(46)(24*8-1 downto 23*8),  
w25 => Pw(46)(25*8-1 downto 24*8), w26 => Pw(46)(26*8-1 downto 25*8), w27 => Pw(46)(27*8-1 downto 26*8), w28 => Pw(46)(28*8-1 downto 27*8), w29 => Pw(46)(29*8-1 downto 28*8), w30 => Pw(46)(30*8-1 downto 29*8), w31 => Pw(46)(31*8-1 downto 30*8), w32 => Pw(46)(32*8-1 downto 31*8),  
w33 => Pw(46)(33*8-1 downto 32*8), w34 => Pw(46)(34*8-1 downto 33*8), w35 => Pw(46)(35*8-1 downto 34*8), w36 => Pw(46)(36*8-1 downto 35*8), w37 => Pw(46)(37*8-1 downto 36*8), w38 => Pw(46)(38*8-1 downto 37*8), w39 => Pw(46)(39*8-1 downto 38*8), w40 => Pw(46)(40*8-1 downto 39*8),  
w41 => Pw(46)(41*8-1 downto 40*8), w42 => Pw(46)(42*8-1 downto 41*8), w43 => Pw(46)(43*8-1 downto 42*8), w44 => Pw(46)(44*8-1 downto 43*8), w45 => Pw(46)(45*8-1 downto 44*8), w46 => Pw(46)(46*8-1 downto 45*8), w47 => Pw(46)(47*8-1 downto 46*8), w48 => Pw(46)(48*8-1 downto 47*8),  
w49 => Pw(46)(49*8-1 downto 48*8), w50 => Pw(46)(50*8-1 downto 49*8), w51 => Pw(46)(51*8-1 downto 50*8), w52 => Pw(46)(52*8-1 downto 51*8), w53 => Pw(46)(53*8-1 downto 52*8), w54 => Pw(46)(54*8-1 downto 53*8), w55 => Pw(46)(55*8-1 downto 54*8), w56 => Pw(46)(56*8-1 downto 55*8),  
w57 => Pw(46)(57*8-1 downto 56*8), w58 => Pw(46)(58*8-1 downto 57*8), w59 => Pw(46)(59*8-1 downto 58*8), w60 => Pw(46)(60*8-1 downto 59*8), w61 => Pw(46)(61*8-1 downto 60*8), w62 => Pw(46)(62*8-1 downto 61*8), w63 => Pw(46)(63*8-1 downto 62*8), w64 => Pw(46)(64*8-1 downto 63*8), 
w65 => Pw(46)( 65*8-1 downto  64*8), w66 => Pw(46)( 66*8-1 downto  65*8), w67 => Pw(46)( 67*8-1 downto  66*8), w68 => Pw(46)( 68*8-1 downto  67*8), w69 => Pw(46)( 69*8-1 downto  68*8), w70 => Pw(46)( 70*8-1 downto  69*8), w71 => Pw(46)( 71*8-1 downto  70*8), w72 => Pw(46)( 72*8-1 downto  71*8), 
w73 => Pw(46)( 73*8-1 downto  72*8), w74 => Pw(46)( 74*8-1 downto  73*8), w75 => Pw(46)( 75*8-1 downto  74*8), w76 => Pw(46)( 76*8-1 downto  75*8), w77 => Pw(46)( 77*8-1 downto  76*8), w78 => Pw(46)( 78*8-1 downto  77*8), w79 => Pw(46)( 79*8-1 downto  78*8), w80 => Pw(46)( 80*8-1 downto  79*8), 
w81 => Pw(46)( 81*8-1 downto  80*8), w82 => Pw(46)( 82*8-1 downto  81*8), w83 => Pw(46)( 83*8-1 downto  82*8), w84 => Pw(46)( 84*8-1 downto  83*8), w85 => Pw(46)( 85*8-1 downto  84*8), w86 => Pw(46)( 86*8-1 downto  85*8), w87 => Pw(46)( 87*8-1 downto  86*8), w88 => Pw(46)( 88*8-1 downto  87*8), 
w89 => Pw(46)( 89*8-1 downto  88*8), w90 => Pw(46)( 90*8-1 downto  89*8), w91 => Pw(46)( 91*8-1 downto  90*8), w92 => Pw(46)( 92*8-1 downto  91*8), w93 => Pw(46)( 93*8-1 downto  92*8), w94 => Pw(46)( 94*8-1 downto  93*8), w95 => Pw(46)( 95*8-1 downto  94*8), w96 => Pw(46)( 96*8-1 downto  95*8), 
w97 => Pw(46)( 97*8-1 downto  96*8), w98 => Pw(46)( 98*8-1 downto  97*8), w99 => Pw(46)( 99*8-1 downto  98*8), w100=> Pw(46)(100*8-1 downto  99*8), w101=> Pw(46)(101*8-1 downto 100*8), w102=> Pw(46)(102*8-1 downto 101*8), w103=> Pw(46)(103*8-1 downto 102*8), w104=> Pw(46)(104*8-1 downto 103*8), 
w105=> Pw(46)(105*8-1 downto 104*8), w106=> Pw(46)(106*8-1 downto 105*8), w107=> Pw(46)(107*8-1 downto 106*8), w108=> Pw(46)(108*8-1 downto 107*8), w109=> Pw(46)(109*8-1 downto 108*8), w110=> Pw(46)(110*8-1 downto 109*8), w111=> Pw(46)(111*8-1 downto 110*8), w112=> Pw(46)(112*8-1 downto 111*8), 
w113=> Pw(46)(113*8-1 downto 112*8), w114=> Pw(46)(114*8-1 downto 113*8), w115=> Pw(46)(115*8-1 downto 114*8), w116=> Pw(46)(116*8-1 downto 115*8), w117=> Pw(46)(117*8-1 downto 116*8), w118=> Pw(46)(118*8-1 downto 117*8), w119=> Pw(46)(119*8-1 downto 118*8), w120=> Pw(46)(120*8-1 downto 119*8), 
w121=> Pw(46)(121*8-1 downto 120*8), w122=> Pw(46)(122*8-1 downto 121*8), w123=> Pw(46)(123*8-1 downto 122*8), w124=> Pw(46)(124*8-1 downto 123*8), w125=> Pw(46)(125*8-1 downto 124*8), w126=> Pw(46)(126*8-1 downto 125*8), w127=> Pw(46)(127*8-1 downto 126*8), w128=> Pw(46)(128*8-1 downto 127*8), 

           d_out   => pca_d46_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_47_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(47)(     7 downto    0), w02 => Pw(47)( 2*8-1 downto    8), w03 => Pw(47)( 3*8-1 downto  2*8), w04 => Pw(47)( 4*8-1 downto  3*8), w05 => Pw(47)( 5*8-1 downto  4*8), w06 => Pw(47)( 6*8-1 downto  5*8), w07 => Pw(47)( 7*8-1 downto  6*8), w08 => Pw(47)( 8*8-1 downto  7*8),  
w09 => Pw(47)( 9*8-1 downto  8*8), w10 => Pw(47)(10*8-1 downto  9*8), w11 => Pw(47)(11*8-1 downto 10*8), w12 => Pw(47)(12*8-1 downto 11*8), w13 => Pw(47)(13*8-1 downto 12*8), w14 => Pw(47)(14*8-1 downto 13*8), w15 => Pw(47)(15*8-1 downto 14*8), w16 => Pw(47)(16*8-1 downto 15*8),  
w17 => Pw(47)(17*8-1 downto 16*8), w18 => Pw(47)(18*8-1 downto 17*8), w19 => Pw(47)(19*8-1 downto 18*8), w20 => Pw(47)(20*8-1 downto 19*8), w21 => Pw(47)(21*8-1 downto 20*8), w22 => Pw(47)(22*8-1 downto 21*8), w23 => Pw(47)(23*8-1 downto 22*8), w24 => Pw(47)(24*8-1 downto 23*8),  
w25 => Pw(47)(25*8-1 downto 24*8), w26 => Pw(47)(26*8-1 downto 25*8), w27 => Pw(47)(27*8-1 downto 26*8), w28 => Pw(47)(28*8-1 downto 27*8), w29 => Pw(47)(29*8-1 downto 28*8), w30 => Pw(47)(30*8-1 downto 29*8), w31 => Pw(47)(31*8-1 downto 30*8), w32 => Pw(47)(32*8-1 downto 31*8),  
w33 => Pw(47)(33*8-1 downto 32*8), w34 => Pw(47)(34*8-1 downto 33*8), w35 => Pw(47)(35*8-1 downto 34*8), w36 => Pw(47)(36*8-1 downto 35*8), w37 => Pw(47)(37*8-1 downto 36*8), w38 => Pw(47)(38*8-1 downto 37*8), w39 => Pw(47)(39*8-1 downto 38*8), w40 => Pw(47)(40*8-1 downto 39*8),  
w41 => Pw(47)(41*8-1 downto 40*8), w42 => Pw(47)(42*8-1 downto 41*8), w43 => Pw(47)(43*8-1 downto 42*8), w44 => Pw(47)(44*8-1 downto 43*8), w45 => Pw(47)(45*8-1 downto 44*8), w46 => Pw(47)(46*8-1 downto 45*8), w47 => Pw(47)(47*8-1 downto 46*8), w48 => Pw(47)(48*8-1 downto 47*8),  
w49 => Pw(47)(49*8-1 downto 48*8), w50 => Pw(47)(50*8-1 downto 49*8), w51 => Pw(47)(51*8-1 downto 50*8), w52 => Pw(47)(52*8-1 downto 51*8), w53 => Pw(47)(53*8-1 downto 52*8), w54 => Pw(47)(54*8-1 downto 53*8), w55 => Pw(47)(55*8-1 downto 54*8), w56 => Pw(47)(56*8-1 downto 55*8),  
w57 => Pw(47)(57*8-1 downto 56*8), w58 => Pw(47)(58*8-1 downto 57*8), w59 => Pw(47)(59*8-1 downto 58*8), w60 => Pw(47)(60*8-1 downto 59*8), w61 => Pw(47)(61*8-1 downto 60*8), w62 => Pw(47)(62*8-1 downto 61*8), w63 => Pw(47)(63*8-1 downto 62*8), w64 => Pw(47)(64*8-1 downto 63*8), 
w65 => Pw(47)( 65*8-1 downto  64*8), w66 => Pw(47)( 66*8-1 downto  65*8), w67 => Pw(47)( 67*8-1 downto  66*8), w68 => Pw(47)( 68*8-1 downto  67*8), w69 => Pw(47)( 69*8-1 downto  68*8), w70 => Pw(47)( 70*8-1 downto  69*8), w71 => Pw(47)( 71*8-1 downto  70*8), w72 => Pw(47)( 72*8-1 downto  71*8), 
w73 => Pw(47)( 73*8-1 downto  72*8), w74 => Pw(47)( 74*8-1 downto  73*8), w75 => Pw(47)( 75*8-1 downto  74*8), w76 => Pw(47)( 76*8-1 downto  75*8), w77 => Pw(47)( 77*8-1 downto  76*8), w78 => Pw(47)( 78*8-1 downto  77*8), w79 => Pw(47)( 79*8-1 downto  78*8), w80 => Pw(47)( 80*8-1 downto  79*8), 
w81 => Pw(47)( 81*8-1 downto  80*8), w82 => Pw(47)( 82*8-1 downto  81*8), w83 => Pw(47)( 83*8-1 downto  82*8), w84 => Pw(47)( 84*8-1 downto  83*8), w85 => Pw(47)( 85*8-1 downto  84*8), w86 => Pw(47)( 86*8-1 downto  85*8), w87 => Pw(47)( 87*8-1 downto  86*8), w88 => Pw(47)( 88*8-1 downto  87*8), 
w89 => Pw(47)( 89*8-1 downto  88*8), w90 => Pw(47)( 90*8-1 downto  89*8), w91 => Pw(47)( 91*8-1 downto  90*8), w92 => Pw(47)( 92*8-1 downto  91*8), w93 => Pw(47)( 93*8-1 downto  92*8), w94 => Pw(47)( 94*8-1 downto  93*8), w95 => Pw(47)( 95*8-1 downto  94*8), w96 => Pw(47)( 96*8-1 downto  95*8), 
w97 => Pw(47)( 97*8-1 downto  96*8), w98 => Pw(47)( 98*8-1 downto  97*8), w99 => Pw(47)( 99*8-1 downto  98*8), w100=> Pw(47)(100*8-1 downto  99*8), w101=> Pw(47)(101*8-1 downto 100*8), w102=> Pw(47)(102*8-1 downto 101*8), w103=> Pw(47)(103*8-1 downto 102*8), w104=> Pw(47)(104*8-1 downto 103*8), 
w105=> Pw(47)(105*8-1 downto 104*8), w106=> Pw(47)(106*8-1 downto 105*8), w107=> Pw(47)(107*8-1 downto 106*8), w108=> Pw(47)(108*8-1 downto 107*8), w109=> Pw(47)(109*8-1 downto 108*8), w110=> Pw(47)(110*8-1 downto 109*8), w111=> Pw(47)(111*8-1 downto 110*8), w112=> Pw(47)(112*8-1 downto 111*8), 
w113=> Pw(47)(113*8-1 downto 112*8), w114=> Pw(47)(114*8-1 downto 113*8), w115=> Pw(47)(115*8-1 downto 114*8), w116=> Pw(47)(116*8-1 downto 115*8), w117=> Pw(47)(117*8-1 downto 116*8), w118=> Pw(47)(118*8-1 downto 117*8), w119=> Pw(47)(119*8-1 downto 118*8), w120=> Pw(47)(120*8-1 downto 119*8), 
w121=> Pw(47)(121*8-1 downto 120*8), w122=> Pw(47)(122*8-1 downto 121*8), w123=> Pw(47)(123*8-1 downto 122*8), w124=> Pw(47)(124*8-1 downto 123*8), w125=> Pw(47)(125*8-1 downto 124*8), w126=> Pw(47)(126*8-1 downto 125*8), w127=> Pw(47)(127*8-1 downto 126*8), w128=> Pw(47)(128*8-1 downto 127*8), 

           d_out   => pca_d47_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_48_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(48)(     7 downto    0), w02 => Pw(48)( 2*8-1 downto    8), w03 => Pw(48)( 3*8-1 downto  2*8), w04 => Pw(48)( 4*8-1 downto  3*8), w05 => Pw(48)( 5*8-1 downto  4*8), w06 => Pw(48)( 6*8-1 downto  5*8), w07 => Pw(48)( 7*8-1 downto  6*8), w08 => Pw(48)( 8*8-1 downto  7*8),  
w09 => Pw(48)( 9*8-1 downto  8*8), w10 => Pw(48)(10*8-1 downto  9*8), w11 => Pw(48)(11*8-1 downto 10*8), w12 => Pw(48)(12*8-1 downto 11*8), w13 => Pw(48)(13*8-1 downto 12*8), w14 => Pw(48)(14*8-1 downto 13*8), w15 => Pw(48)(15*8-1 downto 14*8), w16 => Pw(48)(16*8-1 downto 15*8),  
w17 => Pw(48)(17*8-1 downto 16*8), w18 => Pw(48)(18*8-1 downto 17*8), w19 => Pw(48)(19*8-1 downto 18*8), w20 => Pw(48)(20*8-1 downto 19*8), w21 => Pw(48)(21*8-1 downto 20*8), w22 => Pw(48)(22*8-1 downto 21*8), w23 => Pw(48)(23*8-1 downto 22*8), w24 => Pw(48)(24*8-1 downto 23*8),  
w25 => Pw(48)(25*8-1 downto 24*8), w26 => Pw(48)(26*8-1 downto 25*8), w27 => Pw(48)(27*8-1 downto 26*8), w28 => Pw(48)(28*8-1 downto 27*8), w29 => Pw(48)(29*8-1 downto 28*8), w30 => Pw(48)(30*8-1 downto 29*8), w31 => Pw(48)(31*8-1 downto 30*8), w32 => Pw(48)(32*8-1 downto 31*8),  
w33 => Pw(48)(33*8-1 downto 32*8), w34 => Pw(48)(34*8-1 downto 33*8), w35 => Pw(48)(35*8-1 downto 34*8), w36 => Pw(48)(36*8-1 downto 35*8), w37 => Pw(48)(37*8-1 downto 36*8), w38 => Pw(48)(38*8-1 downto 37*8), w39 => Pw(48)(39*8-1 downto 38*8), w40 => Pw(48)(40*8-1 downto 39*8),  
w41 => Pw(48)(41*8-1 downto 40*8), w42 => Pw(48)(42*8-1 downto 41*8), w43 => Pw(48)(43*8-1 downto 42*8), w44 => Pw(48)(44*8-1 downto 43*8), w45 => Pw(48)(45*8-1 downto 44*8), w46 => Pw(48)(46*8-1 downto 45*8), w47 => Pw(48)(47*8-1 downto 46*8), w48 => Pw(48)(48*8-1 downto 47*8),  
w49 => Pw(48)(49*8-1 downto 48*8), w50 => Pw(48)(50*8-1 downto 49*8), w51 => Pw(48)(51*8-1 downto 50*8), w52 => Pw(48)(52*8-1 downto 51*8), w53 => Pw(48)(53*8-1 downto 52*8), w54 => Pw(48)(54*8-1 downto 53*8), w55 => Pw(48)(55*8-1 downto 54*8), w56 => Pw(48)(56*8-1 downto 55*8),  
w57 => Pw(48)(57*8-1 downto 56*8), w58 => Pw(48)(58*8-1 downto 57*8), w59 => Pw(48)(59*8-1 downto 58*8), w60 => Pw(48)(60*8-1 downto 59*8), w61 => Pw(48)(61*8-1 downto 60*8), w62 => Pw(48)(62*8-1 downto 61*8), w63 => Pw(48)(63*8-1 downto 62*8), w64 => Pw(48)(64*8-1 downto 63*8), 
w65 => Pw(48)( 65*8-1 downto  64*8), w66 => Pw(48)( 66*8-1 downto  65*8), w67 => Pw(48)( 67*8-1 downto  66*8), w68 => Pw(48)( 68*8-1 downto  67*8), w69 => Pw(48)( 69*8-1 downto  68*8), w70 => Pw(48)( 70*8-1 downto  69*8), w71 => Pw(48)( 71*8-1 downto  70*8), w72 => Pw(48)( 72*8-1 downto  71*8), 
w73 => Pw(48)( 73*8-1 downto  72*8), w74 => Pw(48)( 74*8-1 downto  73*8), w75 => Pw(48)( 75*8-1 downto  74*8), w76 => Pw(48)( 76*8-1 downto  75*8), w77 => Pw(48)( 77*8-1 downto  76*8), w78 => Pw(48)( 78*8-1 downto  77*8), w79 => Pw(48)( 79*8-1 downto  78*8), w80 => Pw(48)( 80*8-1 downto  79*8), 
w81 => Pw(48)( 81*8-1 downto  80*8), w82 => Pw(48)( 82*8-1 downto  81*8), w83 => Pw(48)( 83*8-1 downto  82*8), w84 => Pw(48)( 84*8-1 downto  83*8), w85 => Pw(48)( 85*8-1 downto  84*8), w86 => Pw(48)( 86*8-1 downto  85*8), w87 => Pw(48)( 87*8-1 downto  86*8), w88 => Pw(48)( 88*8-1 downto  87*8), 
w89 => Pw(48)( 89*8-1 downto  88*8), w90 => Pw(48)( 90*8-1 downto  89*8), w91 => Pw(48)( 91*8-1 downto  90*8), w92 => Pw(48)( 92*8-1 downto  91*8), w93 => Pw(48)( 93*8-1 downto  92*8), w94 => Pw(48)( 94*8-1 downto  93*8), w95 => Pw(48)( 95*8-1 downto  94*8), w96 => Pw(48)( 96*8-1 downto  95*8), 
w97 => Pw(48)( 97*8-1 downto  96*8), w98 => Pw(48)( 98*8-1 downto  97*8), w99 => Pw(48)( 99*8-1 downto  98*8), w100=> Pw(48)(100*8-1 downto  99*8), w101=> Pw(48)(101*8-1 downto 100*8), w102=> Pw(48)(102*8-1 downto 101*8), w103=> Pw(48)(103*8-1 downto 102*8), w104=> Pw(48)(104*8-1 downto 103*8), 
w105=> Pw(48)(105*8-1 downto 104*8), w106=> Pw(48)(106*8-1 downto 105*8), w107=> Pw(48)(107*8-1 downto 106*8), w108=> Pw(48)(108*8-1 downto 107*8), w109=> Pw(48)(109*8-1 downto 108*8), w110=> Pw(48)(110*8-1 downto 109*8), w111=> Pw(48)(111*8-1 downto 110*8), w112=> Pw(48)(112*8-1 downto 111*8), 
w113=> Pw(48)(113*8-1 downto 112*8), w114=> Pw(48)(114*8-1 downto 113*8), w115=> Pw(48)(115*8-1 downto 114*8), w116=> Pw(48)(116*8-1 downto 115*8), w117=> Pw(48)(117*8-1 downto 116*8), w118=> Pw(48)(118*8-1 downto 117*8), w119=> Pw(48)(119*8-1 downto 118*8), w120=> Pw(48)(120*8-1 downto 119*8), 
w121=> Pw(48)(121*8-1 downto 120*8), w122=> Pw(48)(122*8-1 downto 121*8), w123=> Pw(48)(123*8-1 downto 122*8), w124=> Pw(48)(124*8-1 downto 123*8), w125=> Pw(48)(125*8-1 downto 124*8), w126=> Pw(48)(126*8-1 downto 125*8), w127=> Pw(48)(127*8-1 downto 126*8), w128=> Pw(48)(128*8-1 downto 127*8), 

           d_out   => pca_d48_out   ,
           en_out  => open  ,
           sof_out => open );

  
  PCA128_49_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(49)(     7 downto    0), w02 => Pw(49)( 2*8-1 downto    8), w03 => Pw(49)( 3*8-1 downto  2*8), w04 => Pw(49)( 4*8-1 downto  3*8), w05 => Pw(49)( 5*8-1 downto  4*8), w06 => Pw(49)( 6*8-1 downto  5*8), w07 => Pw(49)( 7*8-1 downto  6*8), w08 => Pw(49)( 8*8-1 downto  7*8),  
w09 => Pw(49)( 9*8-1 downto  8*8), w10 => Pw(49)(10*8-1 downto  9*8), w11 => Pw(49)(11*8-1 downto 10*8), w12 => Pw(49)(12*8-1 downto 11*8), w13 => Pw(49)(13*8-1 downto 12*8), w14 => Pw(49)(14*8-1 downto 13*8), w15 => Pw(49)(15*8-1 downto 14*8), w16 => Pw(49)(16*8-1 downto 15*8),  
w17 => Pw(49)(17*8-1 downto 16*8), w18 => Pw(49)(18*8-1 downto 17*8), w19 => Pw(49)(19*8-1 downto 18*8), w20 => Pw(49)(20*8-1 downto 19*8), w21 => Pw(49)(21*8-1 downto 20*8), w22 => Pw(49)(22*8-1 downto 21*8), w23 => Pw(49)(23*8-1 downto 22*8), w24 => Pw(49)(24*8-1 downto 23*8),  
w25 => Pw(49)(25*8-1 downto 24*8), w26 => Pw(49)(26*8-1 downto 25*8), w27 => Pw(49)(27*8-1 downto 26*8), w28 => Pw(49)(28*8-1 downto 27*8), w29 => Pw(49)(29*8-1 downto 28*8), w30 => Pw(49)(30*8-1 downto 29*8), w31 => Pw(49)(31*8-1 downto 30*8), w32 => Pw(49)(32*8-1 downto 31*8),  
w33 => Pw(49)(33*8-1 downto 32*8), w34 => Pw(49)(34*8-1 downto 33*8), w35 => Pw(49)(35*8-1 downto 34*8), w36 => Pw(49)(36*8-1 downto 35*8), w37 => Pw(49)(37*8-1 downto 36*8), w38 => Pw(49)(38*8-1 downto 37*8), w39 => Pw(49)(39*8-1 downto 38*8), w40 => Pw(49)(40*8-1 downto 39*8),  
w41 => Pw(49)(41*8-1 downto 40*8), w42 => Pw(49)(42*8-1 downto 41*8), w43 => Pw(49)(43*8-1 downto 42*8), w44 => Pw(49)(44*8-1 downto 43*8), w45 => Pw(49)(45*8-1 downto 44*8), w46 => Pw(49)(46*8-1 downto 45*8), w47 => Pw(49)(47*8-1 downto 46*8), w48 => Pw(49)(48*8-1 downto 47*8),  
w49 => Pw(49)(49*8-1 downto 48*8), w50 => Pw(49)(50*8-1 downto 49*8), w51 => Pw(49)(51*8-1 downto 50*8), w52 => Pw(49)(52*8-1 downto 51*8), w53 => Pw(49)(53*8-1 downto 52*8), w54 => Pw(49)(54*8-1 downto 53*8), w55 => Pw(49)(55*8-1 downto 54*8), w56 => Pw(49)(56*8-1 downto 55*8),  
w57 => Pw(49)(57*8-1 downto 56*8), w58 => Pw(49)(58*8-1 downto 57*8), w59 => Pw(49)(59*8-1 downto 58*8), w60 => Pw(49)(60*8-1 downto 59*8), w61 => Pw(49)(61*8-1 downto 60*8), w62 => Pw(49)(62*8-1 downto 61*8), w63 => Pw(49)(63*8-1 downto 62*8), w64 => Pw(49)(64*8-1 downto 63*8), 
w65 => Pw(49)( 65*8-1 downto  64*8), w66 => Pw(49)( 66*8-1 downto  65*8), w67 => Pw(49)( 67*8-1 downto  66*8), w68 => Pw(49)( 68*8-1 downto  67*8), w69 => Pw(49)( 69*8-1 downto  68*8), w70 => Pw(49)( 70*8-1 downto  69*8), w71 => Pw(49)( 71*8-1 downto  70*8), w72 => Pw(49)( 72*8-1 downto  71*8), 
w73 => Pw(49)( 73*8-1 downto  72*8), w74 => Pw(49)( 74*8-1 downto  73*8), w75 => Pw(49)( 75*8-1 downto  74*8), w76 => Pw(49)( 76*8-1 downto  75*8), w77 => Pw(49)( 77*8-1 downto  76*8), w78 => Pw(49)( 78*8-1 downto  77*8), w79 => Pw(49)( 79*8-1 downto  78*8), w80 => Pw(49)( 80*8-1 downto  79*8), 
w81 => Pw(49)( 81*8-1 downto  80*8), w82 => Pw(49)( 82*8-1 downto  81*8), w83 => Pw(49)( 83*8-1 downto  82*8), w84 => Pw(49)( 84*8-1 downto  83*8), w85 => Pw(49)( 85*8-1 downto  84*8), w86 => Pw(49)( 86*8-1 downto  85*8), w87 => Pw(49)( 87*8-1 downto  86*8), w88 => Pw(49)( 88*8-1 downto  87*8), 
w89 => Pw(49)( 89*8-1 downto  88*8), w90 => Pw(49)( 90*8-1 downto  89*8), w91 => Pw(49)( 91*8-1 downto  90*8), w92 => Pw(49)( 92*8-1 downto  91*8), w93 => Pw(49)( 93*8-1 downto  92*8), w94 => Pw(49)( 94*8-1 downto  93*8), w95 => Pw(49)( 95*8-1 downto  94*8), w96 => Pw(49)( 96*8-1 downto  95*8), 
w97 => Pw(49)( 97*8-1 downto  96*8), w98 => Pw(49)( 98*8-1 downto  97*8), w99 => Pw(49)( 99*8-1 downto  98*8), w100=> Pw(49)(100*8-1 downto  99*8), w101=> Pw(49)(101*8-1 downto 100*8), w102=> Pw(49)(102*8-1 downto 101*8), w103=> Pw(49)(103*8-1 downto 102*8), w104=> Pw(49)(104*8-1 downto 103*8), 
w105=> Pw(49)(105*8-1 downto 104*8), w106=> Pw(49)(106*8-1 downto 105*8), w107=> Pw(49)(107*8-1 downto 106*8), w108=> Pw(49)(108*8-1 downto 107*8), w109=> Pw(49)(109*8-1 downto 108*8), w110=> Pw(49)(110*8-1 downto 109*8), w111=> Pw(49)(111*8-1 downto 110*8), w112=> Pw(49)(112*8-1 downto 111*8), 
w113=> Pw(49)(113*8-1 downto 112*8), w114=> Pw(49)(114*8-1 downto 113*8), w115=> Pw(49)(115*8-1 downto 114*8), w116=> Pw(49)(116*8-1 downto 115*8), w117=> Pw(49)(117*8-1 downto 116*8), w118=> Pw(49)(118*8-1 downto 117*8), w119=> Pw(49)(119*8-1 downto 118*8), w120=> Pw(49)(120*8-1 downto 119*8), 
w121=> Pw(49)(121*8-1 downto 120*8), w122=> Pw(49)(122*8-1 downto 121*8), w123=> Pw(49)(123*8-1 downto 122*8), w124=> Pw(49)(124*8-1 downto 123*8), w125=> Pw(49)(125*8-1 downto 124*8), w126=> Pw(49)(126*8-1 downto 125*8), w127=> Pw(49)(127*8-1 downto 126*8), w128=> Pw(49)(128*8-1 downto 127*8), 

           d_out   => pca_d49_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_50_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(50)(     7 downto    0), w02 => Pw(50)( 2*8-1 downto    8), w03 => Pw(50)( 3*8-1 downto  2*8), w04 => Pw(50)( 4*8-1 downto  3*8), w05 => Pw(50)( 5*8-1 downto  4*8), w06 => Pw(50)( 6*8-1 downto  5*8), w07 => Pw(50)( 7*8-1 downto  6*8), w08 => Pw(50)( 8*8-1 downto  7*8),  
w09 => Pw(50)( 9*8-1 downto  8*8), w10 => Pw(50)(10*8-1 downto  9*8), w11 => Pw(50)(11*8-1 downto 10*8), w12 => Pw(50)(12*8-1 downto 11*8), w13 => Pw(50)(13*8-1 downto 12*8), w14 => Pw(50)(14*8-1 downto 13*8), w15 => Pw(50)(15*8-1 downto 14*8), w16 => Pw(50)(16*8-1 downto 15*8),  
w17 => Pw(50)(17*8-1 downto 16*8), w18 => Pw(50)(18*8-1 downto 17*8), w19 => Pw(50)(19*8-1 downto 18*8), w20 => Pw(50)(20*8-1 downto 19*8), w21 => Pw(50)(21*8-1 downto 20*8), w22 => Pw(50)(22*8-1 downto 21*8), w23 => Pw(50)(23*8-1 downto 22*8), w24 => Pw(50)(24*8-1 downto 23*8),  
w25 => Pw(50)(25*8-1 downto 24*8), w26 => Pw(50)(26*8-1 downto 25*8), w27 => Pw(50)(27*8-1 downto 26*8), w28 => Pw(50)(28*8-1 downto 27*8), w29 => Pw(50)(29*8-1 downto 28*8), w30 => Pw(50)(30*8-1 downto 29*8), w31 => Pw(50)(31*8-1 downto 30*8), w32 => Pw(50)(32*8-1 downto 31*8),  
w33 => Pw(50)(33*8-1 downto 32*8), w34 => Pw(50)(34*8-1 downto 33*8), w35 => Pw(50)(35*8-1 downto 34*8), w36 => Pw(50)(36*8-1 downto 35*8), w37 => Pw(50)(37*8-1 downto 36*8), w38 => Pw(50)(38*8-1 downto 37*8), w39 => Pw(50)(39*8-1 downto 38*8), w40 => Pw(50)(40*8-1 downto 39*8),  
w41 => Pw(50)(41*8-1 downto 40*8), w42 => Pw(50)(42*8-1 downto 41*8), w43 => Pw(50)(43*8-1 downto 42*8), w44 => Pw(50)(44*8-1 downto 43*8), w45 => Pw(50)(45*8-1 downto 44*8), w46 => Pw(50)(46*8-1 downto 45*8), w47 => Pw(50)(47*8-1 downto 46*8), w48 => Pw(50)(48*8-1 downto 47*8),  
w49 => Pw(50)(49*8-1 downto 48*8), w50 => Pw(50)(50*8-1 downto 49*8), w51 => Pw(50)(51*8-1 downto 50*8), w52 => Pw(50)(52*8-1 downto 51*8), w53 => Pw(50)(53*8-1 downto 52*8), w54 => Pw(50)(54*8-1 downto 53*8), w55 => Pw(50)(55*8-1 downto 54*8), w56 => Pw(50)(56*8-1 downto 55*8),  
w57 => Pw(50)(57*8-1 downto 56*8), w58 => Pw(50)(58*8-1 downto 57*8), w59 => Pw(50)(59*8-1 downto 58*8), w60 => Pw(50)(60*8-1 downto 59*8), w61 => Pw(50)(61*8-1 downto 60*8), w62 => Pw(50)(62*8-1 downto 61*8), w63 => Pw(50)(63*8-1 downto 62*8), w64 => Pw(50)(64*8-1 downto 63*8), 
w65 => Pw(50)( 65*8-1 downto  64*8), w66 => Pw(50)( 66*8-1 downto  65*8), w67 => Pw(50)( 67*8-1 downto  66*8), w68 => Pw(50)( 68*8-1 downto  67*8), w69 => Pw(50)( 69*8-1 downto  68*8), w70 => Pw(50)( 70*8-1 downto  69*8), w71 => Pw(50)( 71*8-1 downto  70*8), w72 => Pw(50)( 72*8-1 downto  71*8), 
w73 => Pw(50)( 73*8-1 downto  72*8), w74 => Pw(50)( 74*8-1 downto  73*8), w75 => Pw(50)( 75*8-1 downto  74*8), w76 => Pw(50)( 76*8-1 downto  75*8), w77 => Pw(50)( 77*8-1 downto  76*8), w78 => Pw(50)( 78*8-1 downto  77*8), w79 => Pw(50)( 79*8-1 downto  78*8), w80 => Pw(50)( 80*8-1 downto  79*8), 
w81 => Pw(50)( 81*8-1 downto  80*8), w82 => Pw(50)( 82*8-1 downto  81*8), w83 => Pw(50)( 83*8-1 downto  82*8), w84 => Pw(50)( 84*8-1 downto  83*8), w85 => Pw(50)( 85*8-1 downto  84*8), w86 => Pw(50)( 86*8-1 downto  85*8), w87 => Pw(50)( 87*8-1 downto  86*8), w88 => Pw(50)( 88*8-1 downto  87*8), 
w89 => Pw(50)( 89*8-1 downto  88*8), w90 => Pw(50)( 90*8-1 downto  89*8), w91 => Pw(50)( 91*8-1 downto  90*8), w92 => Pw(50)( 92*8-1 downto  91*8), w93 => Pw(50)( 93*8-1 downto  92*8), w94 => Pw(50)( 94*8-1 downto  93*8), w95 => Pw(50)( 95*8-1 downto  94*8), w96 => Pw(50)( 96*8-1 downto  95*8), 
w97 => Pw(50)( 97*8-1 downto  96*8), w98 => Pw(50)( 98*8-1 downto  97*8), w99 => Pw(50)( 99*8-1 downto  98*8), w100=> Pw(50)(100*8-1 downto  99*8), w101=> Pw(50)(101*8-1 downto 100*8), w102=> Pw(50)(102*8-1 downto 101*8), w103=> Pw(50)(103*8-1 downto 102*8), w104=> Pw(50)(104*8-1 downto 103*8), 
w105=> Pw(50)(105*8-1 downto 104*8), w106=> Pw(50)(106*8-1 downto 105*8), w107=> Pw(50)(107*8-1 downto 106*8), w108=> Pw(50)(108*8-1 downto 107*8), w109=> Pw(50)(109*8-1 downto 108*8), w110=> Pw(50)(110*8-1 downto 109*8), w111=> Pw(50)(111*8-1 downto 110*8), w112=> Pw(50)(112*8-1 downto 111*8), 
w113=> Pw(50)(113*8-1 downto 112*8), w114=> Pw(50)(114*8-1 downto 113*8), w115=> Pw(50)(115*8-1 downto 114*8), w116=> Pw(50)(116*8-1 downto 115*8), w117=> Pw(50)(117*8-1 downto 116*8), w118=> Pw(50)(118*8-1 downto 117*8), w119=> Pw(50)(119*8-1 downto 118*8), w120=> Pw(50)(120*8-1 downto 119*8), 
w121=> Pw(50)(121*8-1 downto 120*8), w122=> Pw(50)(122*8-1 downto 121*8), w123=> Pw(50)(123*8-1 downto 122*8), w124=> Pw(50)(124*8-1 downto 123*8), w125=> Pw(50)(125*8-1 downto 124*8), w126=> Pw(50)(126*8-1 downto 125*8), w127=> Pw(50)(127*8-1 downto 126*8), w128=> Pw(50)(128*8-1 downto 127*8), 

           d_out   => pca_d50_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_51_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(51)(     7 downto    0), w02 => Pw(51)( 2*8-1 downto    8), w03 => Pw(51)( 3*8-1 downto  2*8), w04 => Pw(51)( 4*8-1 downto  3*8), w05 => Pw(51)( 5*8-1 downto  4*8), w06 => Pw(51)( 6*8-1 downto  5*8), w07 => Pw(51)( 7*8-1 downto  6*8), w08 => Pw(51)( 8*8-1 downto  7*8),  
w09 => Pw(51)( 9*8-1 downto  8*8), w10 => Pw(51)(10*8-1 downto  9*8), w11 => Pw(51)(11*8-1 downto 10*8), w12 => Pw(51)(12*8-1 downto 11*8), w13 => Pw(51)(13*8-1 downto 12*8), w14 => Pw(51)(14*8-1 downto 13*8), w15 => Pw(51)(15*8-1 downto 14*8), w16 => Pw(51)(16*8-1 downto 15*8),  
w17 => Pw(51)(17*8-1 downto 16*8), w18 => Pw(51)(18*8-1 downto 17*8), w19 => Pw(51)(19*8-1 downto 18*8), w20 => Pw(51)(20*8-1 downto 19*8), w21 => Pw(51)(21*8-1 downto 20*8), w22 => Pw(51)(22*8-1 downto 21*8), w23 => Pw(51)(23*8-1 downto 22*8), w24 => Pw(51)(24*8-1 downto 23*8),  
w25 => Pw(51)(25*8-1 downto 24*8), w26 => Pw(51)(26*8-1 downto 25*8), w27 => Pw(51)(27*8-1 downto 26*8), w28 => Pw(51)(28*8-1 downto 27*8), w29 => Pw(51)(29*8-1 downto 28*8), w30 => Pw(51)(30*8-1 downto 29*8), w31 => Pw(51)(31*8-1 downto 30*8), w32 => Pw(51)(32*8-1 downto 31*8),  
w33 => Pw(51)(33*8-1 downto 32*8), w34 => Pw(51)(34*8-1 downto 33*8), w35 => Pw(51)(35*8-1 downto 34*8), w36 => Pw(51)(36*8-1 downto 35*8), w37 => Pw(51)(37*8-1 downto 36*8), w38 => Pw(51)(38*8-1 downto 37*8), w39 => Pw(51)(39*8-1 downto 38*8), w40 => Pw(51)(40*8-1 downto 39*8),  
w41 => Pw(51)(41*8-1 downto 40*8), w42 => Pw(51)(42*8-1 downto 41*8), w43 => Pw(51)(43*8-1 downto 42*8), w44 => Pw(51)(44*8-1 downto 43*8), w45 => Pw(51)(45*8-1 downto 44*8), w46 => Pw(51)(46*8-1 downto 45*8), w47 => Pw(51)(47*8-1 downto 46*8), w48 => Pw(51)(48*8-1 downto 47*8),  
w49 => Pw(51)(49*8-1 downto 48*8), w50 => Pw(51)(50*8-1 downto 49*8), w51 => Pw(51)(51*8-1 downto 50*8), w52 => Pw(51)(52*8-1 downto 51*8), w53 => Pw(51)(53*8-1 downto 52*8), w54 => Pw(51)(54*8-1 downto 53*8), w55 => Pw(51)(55*8-1 downto 54*8), w56 => Pw(51)(56*8-1 downto 55*8),  
w57 => Pw(51)(57*8-1 downto 56*8), w58 => Pw(51)(58*8-1 downto 57*8), w59 => Pw(51)(59*8-1 downto 58*8), w60 => Pw(51)(60*8-1 downto 59*8), w61 => Pw(51)(61*8-1 downto 60*8), w62 => Pw(51)(62*8-1 downto 61*8), w63 => Pw(51)(63*8-1 downto 62*8), w64 => Pw(51)(64*8-1 downto 63*8), 
w65 => Pw(51)( 65*8-1 downto  64*8), w66 => Pw(51)( 66*8-1 downto  65*8), w67 => Pw(51)( 67*8-1 downto  66*8), w68 => Pw(51)( 68*8-1 downto  67*8), w69 => Pw(51)( 69*8-1 downto  68*8), w70 => Pw(51)( 70*8-1 downto  69*8), w71 => Pw(51)( 71*8-1 downto  70*8), w72 => Pw(51)( 72*8-1 downto  71*8), 
w73 => Pw(51)( 73*8-1 downto  72*8), w74 => Pw(51)( 74*8-1 downto  73*8), w75 => Pw(51)( 75*8-1 downto  74*8), w76 => Pw(51)( 76*8-1 downto  75*8), w77 => Pw(51)( 77*8-1 downto  76*8), w78 => Pw(51)( 78*8-1 downto  77*8), w79 => Pw(51)( 79*8-1 downto  78*8), w80 => Pw(51)( 80*8-1 downto  79*8), 
w81 => Pw(51)( 81*8-1 downto  80*8), w82 => Pw(51)( 82*8-1 downto  81*8), w83 => Pw(51)( 83*8-1 downto  82*8), w84 => Pw(51)( 84*8-1 downto  83*8), w85 => Pw(51)( 85*8-1 downto  84*8), w86 => Pw(51)( 86*8-1 downto  85*8), w87 => Pw(51)( 87*8-1 downto  86*8), w88 => Pw(51)( 88*8-1 downto  87*8), 
w89 => Pw(51)( 89*8-1 downto  88*8), w90 => Pw(51)( 90*8-1 downto  89*8), w91 => Pw(51)( 91*8-1 downto  90*8), w92 => Pw(51)( 92*8-1 downto  91*8), w93 => Pw(51)( 93*8-1 downto  92*8), w94 => Pw(51)( 94*8-1 downto  93*8), w95 => Pw(51)( 95*8-1 downto  94*8), w96 => Pw(51)( 96*8-1 downto  95*8), 
w97 => Pw(51)( 97*8-1 downto  96*8), w98 => Pw(51)( 98*8-1 downto  97*8), w99 => Pw(51)( 99*8-1 downto  98*8), w100=> Pw(51)(100*8-1 downto  99*8), w101=> Pw(51)(101*8-1 downto 100*8), w102=> Pw(51)(102*8-1 downto 101*8), w103=> Pw(51)(103*8-1 downto 102*8), w104=> Pw(51)(104*8-1 downto 103*8), 
w105=> Pw(51)(105*8-1 downto 104*8), w106=> Pw(51)(106*8-1 downto 105*8), w107=> Pw(51)(107*8-1 downto 106*8), w108=> Pw(51)(108*8-1 downto 107*8), w109=> Pw(51)(109*8-1 downto 108*8), w110=> Pw(51)(110*8-1 downto 109*8), w111=> Pw(51)(111*8-1 downto 110*8), w112=> Pw(51)(112*8-1 downto 111*8), 
w113=> Pw(51)(113*8-1 downto 112*8), w114=> Pw(51)(114*8-1 downto 113*8), w115=> Pw(51)(115*8-1 downto 114*8), w116=> Pw(51)(116*8-1 downto 115*8), w117=> Pw(51)(117*8-1 downto 116*8), w118=> Pw(51)(118*8-1 downto 117*8), w119=> Pw(51)(119*8-1 downto 118*8), w120=> Pw(51)(120*8-1 downto 119*8), 
w121=> Pw(51)(121*8-1 downto 120*8), w122=> Pw(51)(122*8-1 downto 121*8), w123=> Pw(51)(123*8-1 downto 122*8), w124=> Pw(51)(124*8-1 downto 123*8), w125=> Pw(51)(125*8-1 downto 124*8), w126=> Pw(51)(126*8-1 downto 125*8), w127=> Pw(51)(127*8-1 downto 126*8), w128=> Pw(51)(128*8-1 downto 127*8), 

           d_out   => pca_d51_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_52_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(52)(     7 downto    0), w02 => Pw(52)( 2*8-1 downto    8), w03 => Pw(52)( 3*8-1 downto  2*8), w04 => Pw(52)( 4*8-1 downto  3*8), w05 => Pw(52)( 5*8-1 downto  4*8), w06 => Pw(52)( 6*8-1 downto  5*8), w07 => Pw(52)( 7*8-1 downto  6*8), w08 => Pw(52)( 8*8-1 downto  7*8),  
w09 => Pw(52)( 9*8-1 downto  8*8), w10 => Pw(52)(10*8-1 downto  9*8), w11 => Pw(52)(11*8-1 downto 10*8), w12 => Pw(52)(12*8-1 downto 11*8), w13 => Pw(52)(13*8-1 downto 12*8), w14 => Pw(52)(14*8-1 downto 13*8), w15 => Pw(52)(15*8-1 downto 14*8), w16 => Pw(52)(16*8-1 downto 15*8),  
w17 => Pw(52)(17*8-1 downto 16*8), w18 => Pw(52)(18*8-1 downto 17*8), w19 => Pw(52)(19*8-1 downto 18*8), w20 => Pw(52)(20*8-1 downto 19*8), w21 => Pw(52)(21*8-1 downto 20*8), w22 => Pw(52)(22*8-1 downto 21*8), w23 => Pw(52)(23*8-1 downto 22*8), w24 => Pw(52)(24*8-1 downto 23*8),  
w25 => Pw(52)(25*8-1 downto 24*8), w26 => Pw(52)(26*8-1 downto 25*8), w27 => Pw(52)(27*8-1 downto 26*8), w28 => Pw(52)(28*8-1 downto 27*8), w29 => Pw(52)(29*8-1 downto 28*8), w30 => Pw(52)(30*8-1 downto 29*8), w31 => Pw(52)(31*8-1 downto 30*8), w32 => Pw(52)(32*8-1 downto 31*8),  
w33 => Pw(52)(33*8-1 downto 32*8), w34 => Pw(52)(34*8-1 downto 33*8), w35 => Pw(52)(35*8-1 downto 34*8), w36 => Pw(52)(36*8-1 downto 35*8), w37 => Pw(52)(37*8-1 downto 36*8), w38 => Pw(52)(38*8-1 downto 37*8), w39 => Pw(52)(39*8-1 downto 38*8), w40 => Pw(52)(40*8-1 downto 39*8),  
w41 => Pw(52)(41*8-1 downto 40*8), w42 => Pw(52)(42*8-1 downto 41*8), w43 => Pw(52)(43*8-1 downto 42*8), w44 => Pw(52)(44*8-1 downto 43*8), w45 => Pw(52)(45*8-1 downto 44*8), w46 => Pw(52)(46*8-1 downto 45*8), w47 => Pw(52)(47*8-1 downto 46*8), w48 => Pw(52)(48*8-1 downto 47*8),  
w49 => Pw(52)(49*8-1 downto 48*8), w50 => Pw(52)(50*8-1 downto 49*8), w51 => Pw(52)(51*8-1 downto 50*8), w52 => Pw(52)(52*8-1 downto 51*8), w53 => Pw(52)(53*8-1 downto 52*8), w54 => Pw(52)(54*8-1 downto 53*8), w55 => Pw(52)(55*8-1 downto 54*8), w56 => Pw(52)(56*8-1 downto 55*8),  
w57 => Pw(52)(57*8-1 downto 56*8), w58 => Pw(52)(58*8-1 downto 57*8), w59 => Pw(52)(59*8-1 downto 58*8), w60 => Pw(52)(60*8-1 downto 59*8), w61 => Pw(52)(61*8-1 downto 60*8), w62 => Pw(52)(62*8-1 downto 61*8), w63 => Pw(52)(63*8-1 downto 62*8), w64 => Pw(52)(64*8-1 downto 63*8), 
w65 => Pw(52)( 65*8-1 downto  64*8), w66 => Pw(52)( 66*8-1 downto  65*8), w67 => Pw(52)( 67*8-1 downto  66*8), w68 => Pw(52)( 68*8-1 downto  67*8), w69 => Pw(52)( 69*8-1 downto  68*8), w70 => Pw(52)( 70*8-1 downto  69*8), w71 => Pw(52)( 71*8-1 downto  70*8), w72 => Pw(52)( 72*8-1 downto  71*8), 
w73 => Pw(52)( 73*8-1 downto  72*8), w74 => Pw(52)( 74*8-1 downto  73*8), w75 => Pw(52)( 75*8-1 downto  74*8), w76 => Pw(52)( 76*8-1 downto  75*8), w77 => Pw(52)( 77*8-1 downto  76*8), w78 => Pw(52)( 78*8-1 downto  77*8), w79 => Pw(52)( 79*8-1 downto  78*8), w80 => Pw(52)( 80*8-1 downto  79*8), 
w81 => Pw(52)( 81*8-1 downto  80*8), w82 => Pw(52)( 82*8-1 downto  81*8), w83 => Pw(52)( 83*8-1 downto  82*8), w84 => Pw(52)( 84*8-1 downto  83*8), w85 => Pw(52)( 85*8-1 downto  84*8), w86 => Pw(52)( 86*8-1 downto  85*8), w87 => Pw(52)( 87*8-1 downto  86*8), w88 => Pw(52)( 88*8-1 downto  87*8), 
w89 => Pw(52)( 89*8-1 downto  88*8), w90 => Pw(52)( 90*8-1 downto  89*8), w91 => Pw(52)( 91*8-1 downto  90*8), w92 => Pw(52)( 92*8-1 downto  91*8), w93 => Pw(52)( 93*8-1 downto  92*8), w94 => Pw(52)( 94*8-1 downto  93*8), w95 => Pw(52)( 95*8-1 downto  94*8), w96 => Pw(52)( 96*8-1 downto  95*8), 
w97 => Pw(52)( 97*8-1 downto  96*8), w98 => Pw(52)( 98*8-1 downto  97*8), w99 => Pw(52)( 99*8-1 downto  98*8), w100=> Pw(52)(100*8-1 downto  99*8), w101=> Pw(52)(101*8-1 downto 100*8), w102=> Pw(52)(102*8-1 downto 101*8), w103=> Pw(52)(103*8-1 downto 102*8), w104=> Pw(52)(104*8-1 downto 103*8), 
w105=> Pw(52)(105*8-1 downto 104*8), w106=> Pw(52)(106*8-1 downto 105*8), w107=> Pw(52)(107*8-1 downto 106*8), w108=> Pw(52)(108*8-1 downto 107*8), w109=> Pw(52)(109*8-1 downto 108*8), w110=> Pw(52)(110*8-1 downto 109*8), w111=> Pw(52)(111*8-1 downto 110*8), w112=> Pw(52)(112*8-1 downto 111*8), 
w113=> Pw(52)(113*8-1 downto 112*8), w114=> Pw(52)(114*8-1 downto 113*8), w115=> Pw(52)(115*8-1 downto 114*8), w116=> Pw(52)(116*8-1 downto 115*8), w117=> Pw(52)(117*8-1 downto 116*8), w118=> Pw(52)(118*8-1 downto 117*8), w119=> Pw(52)(119*8-1 downto 118*8), w120=> Pw(52)(120*8-1 downto 119*8), 
w121=> Pw(52)(121*8-1 downto 120*8), w122=> Pw(52)(122*8-1 downto 121*8), w123=> Pw(52)(123*8-1 downto 122*8), w124=> Pw(52)(124*8-1 downto 123*8), w125=> Pw(52)(125*8-1 downto 124*8), w126=> Pw(52)(126*8-1 downto 125*8), w127=> Pw(52)(127*8-1 downto 126*8), w128=> Pw(52)(128*8-1 downto 127*8), 

           d_out   => pca_d52_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_53_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(53)(     7 downto    0), w02 => Pw(53)( 2*8-1 downto    8), w03 => Pw(53)( 3*8-1 downto  2*8), w04 => Pw(53)( 4*8-1 downto  3*8), w05 => Pw(53)( 5*8-1 downto  4*8), w06 => Pw(53)( 6*8-1 downto  5*8), w07 => Pw(53)( 7*8-1 downto  6*8), w08 => Pw(53)( 8*8-1 downto  7*8),  
w09 => Pw(53)( 9*8-1 downto  8*8), w10 => Pw(53)(10*8-1 downto  9*8), w11 => Pw(53)(11*8-1 downto 10*8), w12 => Pw(53)(12*8-1 downto 11*8), w13 => Pw(53)(13*8-1 downto 12*8), w14 => Pw(53)(14*8-1 downto 13*8), w15 => Pw(53)(15*8-1 downto 14*8), w16 => Pw(53)(16*8-1 downto 15*8),  
w17 => Pw(53)(17*8-1 downto 16*8), w18 => Pw(53)(18*8-1 downto 17*8), w19 => Pw(53)(19*8-1 downto 18*8), w20 => Pw(53)(20*8-1 downto 19*8), w21 => Pw(53)(21*8-1 downto 20*8), w22 => Pw(53)(22*8-1 downto 21*8), w23 => Pw(53)(23*8-1 downto 22*8), w24 => Pw(53)(24*8-1 downto 23*8),  
w25 => Pw(53)(25*8-1 downto 24*8), w26 => Pw(53)(26*8-1 downto 25*8), w27 => Pw(53)(27*8-1 downto 26*8), w28 => Pw(53)(28*8-1 downto 27*8), w29 => Pw(53)(29*8-1 downto 28*8), w30 => Pw(53)(30*8-1 downto 29*8), w31 => Pw(53)(31*8-1 downto 30*8), w32 => Pw(53)(32*8-1 downto 31*8),  
w33 => Pw(53)(33*8-1 downto 32*8), w34 => Pw(53)(34*8-1 downto 33*8), w35 => Pw(53)(35*8-1 downto 34*8), w36 => Pw(53)(36*8-1 downto 35*8), w37 => Pw(53)(37*8-1 downto 36*8), w38 => Pw(53)(38*8-1 downto 37*8), w39 => Pw(53)(39*8-1 downto 38*8), w40 => Pw(53)(40*8-1 downto 39*8),  
w41 => Pw(53)(41*8-1 downto 40*8), w42 => Pw(53)(42*8-1 downto 41*8), w43 => Pw(53)(43*8-1 downto 42*8), w44 => Pw(53)(44*8-1 downto 43*8), w45 => Pw(53)(45*8-1 downto 44*8), w46 => Pw(53)(46*8-1 downto 45*8), w47 => Pw(53)(47*8-1 downto 46*8), w48 => Pw(53)(48*8-1 downto 47*8),  
w49 => Pw(53)(49*8-1 downto 48*8), w50 => Pw(53)(50*8-1 downto 49*8), w51 => Pw(53)(51*8-1 downto 50*8), w52 => Pw(53)(52*8-1 downto 51*8), w53 => Pw(53)(53*8-1 downto 52*8), w54 => Pw(53)(54*8-1 downto 53*8), w55 => Pw(53)(55*8-1 downto 54*8), w56 => Pw(53)(56*8-1 downto 55*8),  
w57 => Pw(53)(57*8-1 downto 56*8), w58 => Pw(53)(58*8-1 downto 57*8), w59 => Pw(53)(59*8-1 downto 58*8), w60 => Pw(53)(60*8-1 downto 59*8), w61 => Pw(53)(61*8-1 downto 60*8), w62 => Pw(53)(62*8-1 downto 61*8), w63 => Pw(53)(63*8-1 downto 62*8), w64 => Pw(53)(64*8-1 downto 63*8), 
w65 => Pw(53)( 65*8-1 downto  64*8), w66 => Pw(53)( 66*8-1 downto  65*8), w67 => Pw(53)( 67*8-1 downto  66*8), w68 => Pw(53)( 68*8-1 downto  67*8), w69 => Pw(53)( 69*8-1 downto  68*8), w70 => Pw(53)( 70*8-1 downto  69*8), w71 => Pw(53)( 71*8-1 downto  70*8), w72 => Pw(53)( 72*8-1 downto  71*8), 
w73 => Pw(53)( 73*8-1 downto  72*8), w74 => Pw(53)( 74*8-1 downto  73*8), w75 => Pw(53)( 75*8-1 downto  74*8), w76 => Pw(53)( 76*8-1 downto  75*8), w77 => Pw(53)( 77*8-1 downto  76*8), w78 => Pw(53)( 78*8-1 downto  77*8), w79 => Pw(53)( 79*8-1 downto  78*8), w80 => Pw(53)( 80*8-1 downto  79*8), 
w81 => Pw(53)( 81*8-1 downto  80*8), w82 => Pw(53)( 82*8-1 downto  81*8), w83 => Pw(53)( 83*8-1 downto  82*8), w84 => Pw(53)( 84*8-1 downto  83*8), w85 => Pw(53)( 85*8-1 downto  84*8), w86 => Pw(53)( 86*8-1 downto  85*8), w87 => Pw(53)( 87*8-1 downto  86*8), w88 => Pw(53)( 88*8-1 downto  87*8), 
w89 => Pw(53)( 89*8-1 downto  88*8), w90 => Pw(53)( 90*8-1 downto  89*8), w91 => Pw(53)( 91*8-1 downto  90*8), w92 => Pw(53)( 92*8-1 downto  91*8), w93 => Pw(53)( 93*8-1 downto  92*8), w94 => Pw(53)( 94*8-1 downto  93*8), w95 => Pw(53)( 95*8-1 downto  94*8), w96 => Pw(53)( 96*8-1 downto  95*8), 
w97 => Pw(53)( 97*8-1 downto  96*8), w98 => Pw(53)( 98*8-1 downto  97*8), w99 => Pw(53)( 99*8-1 downto  98*8), w100=> Pw(53)(100*8-1 downto  99*8), w101=> Pw(53)(101*8-1 downto 100*8), w102=> Pw(53)(102*8-1 downto 101*8), w103=> Pw(53)(103*8-1 downto 102*8), w104=> Pw(53)(104*8-1 downto 103*8), 
w105=> Pw(53)(105*8-1 downto 104*8), w106=> Pw(53)(106*8-1 downto 105*8), w107=> Pw(53)(107*8-1 downto 106*8), w108=> Pw(53)(108*8-1 downto 107*8), w109=> Pw(53)(109*8-1 downto 108*8), w110=> Pw(53)(110*8-1 downto 109*8), w111=> Pw(53)(111*8-1 downto 110*8), w112=> Pw(53)(112*8-1 downto 111*8), 
w113=> Pw(53)(113*8-1 downto 112*8), w114=> Pw(53)(114*8-1 downto 113*8), w115=> Pw(53)(115*8-1 downto 114*8), w116=> Pw(53)(116*8-1 downto 115*8), w117=> Pw(53)(117*8-1 downto 116*8), w118=> Pw(53)(118*8-1 downto 117*8), w119=> Pw(53)(119*8-1 downto 118*8), w120=> Pw(53)(120*8-1 downto 119*8), 
w121=> Pw(53)(121*8-1 downto 120*8), w122=> Pw(53)(122*8-1 downto 121*8), w123=> Pw(53)(123*8-1 downto 122*8), w124=> Pw(53)(124*8-1 downto 123*8), w125=> Pw(53)(125*8-1 downto 124*8), w126=> Pw(53)(126*8-1 downto 125*8), w127=> Pw(53)(127*8-1 downto 126*8), w128=> Pw(53)(128*8-1 downto 127*8), 

           d_out   => pca_d53_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_54_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(54)(     7 downto    0), w02 => Pw(54)( 2*8-1 downto    8), w03 => Pw(54)( 3*8-1 downto  2*8), w04 => Pw(54)( 4*8-1 downto  3*8), w05 => Pw(54)( 5*8-1 downto  4*8), w06 => Pw(54)( 6*8-1 downto  5*8), w07 => Pw(54)( 7*8-1 downto  6*8), w08 => Pw(54)( 8*8-1 downto  7*8),  
w09 => Pw(54)( 9*8-1 downto  8*8), w10 => Pw(54)(10*8-1 downto  9*8), w11 => Pw(54)(11*8-1 downto 10*8), w12 => Pw(54)(12*8-1 downto 11*8), w13 => Pw(54)(13*8-1 downto 12*8), w14 => Pw(54)(14*8-1 downto 13*8), w15 => Pw(54)(15*8-1 downto 14*8), w16 => Pw(54)(16*8-1 downto 15*8),  
w17 => Pw(54)(17*8-1 downto 16*8), w18 => Pw(54)(18*8-1 downto 17*8), w19 => Pw(54)(19*8-1 downto 18*8), w20 => Pw(54)(20*8-1 downto 19*8), w21 => Pw(54)(21*8-1 downto 20*8), w22 => Pw(54)(22*8-1 downto 21*8), w23 => Pw(54)(23*8-1 downto 22*8), w24 => Pw(54)(24*8-1 downto 23*8),  
w25 => Pw(54)(25*8-1 downto 24*8), w26 => Pw(54)(26*8-1 downto 25*8), w27 => Pw(54)(27*8-1 downto 26*8), w28 => Pw(54)(28*8-1 downto 27*8), w29 => Pw(54)(29*8-1 downto 28*8), w30 => Pw(54)(30*8-1 downto 29*8), w31 => Pw(54)(31*8-1 downto 30*8), w32 => Pw(54)(32*8-1 downto 31*8),  
w33 => Pw(54)(33*8-1 downto 32*8), w34 => Pw(54)(34*8-1 downto 33*8), w35 => Pw(54)(35*8-1 downto 34*8), w36 => Pw(54)(36*8-1 downto 35*8), w37 => Pw(54)(37*8-1 downto 36*8), w38 => Pw(54)(38*8-1 downto 37*8), w39 => Pw(54)(39*8-1 downto 38*8), w40 => Pw(54)(40*8-1 downto 39*8),  
w41 => Pw(54)(41*8-1 downto 40*8), w42 => Pw(54)(42*8-1 downto 41*8), w43 => Pw(54)(43*8-1 downto 42*8), w44 => Pw(54)(44*8-1 downto 43*8), w45 => Pw(54)(45*8-1 downto 44*8), w46 => Pw(54)(46*8-1 downto 45*8), w47 => Pw(54)(47*8-1 downto 46*8), w48 => Pw(54)(48*8-1 downto 47*8),  
w49 => Pw(54)(49*8-1 downto 48*8), w50 => Pw(54)(50*8-1 downto 49*8), w51 => Pw(54)(51*8-1 downto 50*8), w52 => Pw(54)(52*8-1 downto 51*8), w53 => Pw(54)(53*8-1 downto 52*8), w54 => Pw(54)(54*8-1 downto 53*8), w55 => Pw(54)(55*8-1 downto 54*8), w56 => Pw(54)(56*8-1 downto 55*8),  
w57 => Pw(54)(57*8-1 downto 56*8), w58 => Pw(54)(58*8-1 downto 57*8), w59 => Pw(54)(59*8-1 downto 58*8), w60 => Pw(54)(60*8-1 downto 59*8), w61 => Pw(54)(61*8-1 downto 60*8), w62 => Pw(54)(62*8-1 downto 61*8), w63 => Pw(54)(63*8-1 downto 62*8), w64 => Pw(54)(64*8-1 downto 63*8), 
w65 => Pw(54)( 65*8-1 downto  64*8), w66 => Pw(54)( 66*8-1 downto  65*8), w67 => Pw(54)( 67*8-1 downto  66*8), w68 => Pw(54)( 68*8-1 downto  67*8), w69 => Pw(54)( 69*8-1 downto  68*8), w70 => Pw(54)( 70*8-1 downto  69*8), w71 => Pw(54)( 71*8-1 downto  70*8), w72 => Pw(54)( 72*8-1 downto  71*8), 
w73 => Pw(54)( 73*8-1 downto  72*8), w74 => Pw(54)( 74*8-1 downto  73*8), w75 => Pw(54)( 75*8-1 downto  74*8), w76 => Pw(54)( 76*8-1 downto  75*8), w77 => Pw(54)( 77*8-1 downto  76*8), w78 => Pw(54)( 78*8-1 downto  77*8), w79 => Pw(54)( 79*8-1 downto  78*8), w80 => Pw(54)( 80*8-1 downto  79*8), 
w81 => Pw(54)( 81*8-1 downto  80*8), w82 => Pw(54)( 82*8-1 downto  81*8), w83 => Pw(54)( 83*8-1 downto  82*8), w84 => Pw(54)( 84*8-1 downto  83*8), w85 => Pw(54)( 85*8-1 downto  84*8), w86 => Pw(54)( 86*8-1 downto  85*8), w87 => Pw(54)( 87*8-1 downto  86*8), w88 => Pw(54)( 88*8-1 downto  87*8), 
w89 => Pw(54)( 89*8-1 downto  88*8), w90 => Pw(54)( 90*8-1 downto  89*8), w91 => Pw(54)( 91*8-1 downto  90*8), w92 => Pw(54)( 92*8-1 downto  91*8), w93 => Pw(54)( 93*8-1 downto  92*8), w94 => Pw(54)( 94*8-1 downto  93*8), w95 => Pw(54)( 95*8-1 downto  94*8), w96 => Pw(54)( 96*8-1 downto  95*8), 
w97 => Pw(54)( 97*8-1 downto  96*8), w98 => Pw(54)( 98*8-1 downto  97*8), w99 => Pw(54)( 99*8-1 downto  98*8), w100=> Pw(54)(100*8-1 downto  99*8), w101=> Pw(54)(101*8-1 downto 100*8), w102=> Pw(54)(102*8-1 downto 101*8), w103=> Pw(54)(103*8-1 downto 102*8), w104=> Pw(54)(104*8-1 downto 103*8), 
w105=> Pw(54)(105*8-1 downto 104*8), w106=> Pw(54)(106*8-1 downto 105*8), w107=> Pw(54)(107*8-1 downto 106*8), w108=> Pw(54)(108*8-1 downto 107*8), w109=> Pw(54)(109*8-1 downto 108*8), w110=> Pw(54)(110*8-1 downto 109*8), w111=> Pw(54)(111*8-1 downto 110*8), w112=> Pw(54)(112*8-1 downto 111*8), 
w113=> Pw(54)(113*8-1 downto 112*8), w114=> Pw(54)(114*8-1 downto 113*8), w115=> Pw(54)(115*8-1 downto 114*8), w116=> Pw(54)(116*8-1 downto 115*8), w117=> Pw(54)(117*8-1 downto 116*8), w118=> Pw(54)(118*8-1 downto 117*8), w119=> Pw(54)(119*8-1 downto 118*8), w120=> Pw(54)(120*8-1 downto 119*8), 
w121=> Pw(54)(121*8-1 downto 120*8), w122=> Pw(54)(122*8-1 downto 121*8), w123=> Pw(54)(123*8-1 downto 122*8), w124=> Pw(54)(124*8-1 downto 123*8), w125=> Pw(54)(125*8-1 downto 124*8), w126=> Pw(54)(126*8-1 downto 125*8), w127=> Pw(54)(127*8-1 downto 126*8), w128=> Pw(54)(128*8-1 downto 127*8), 

           d_out   => pca_d54_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_55_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(55)(     7 downto    0), w02 => Pw(55)( 2*8-1 downto    8), w03 => Pw(55)( 3*8-1 downto  2*8), w04 => Pw(55)( 4*8-1 downto  3*8), w05 => Pw(55)( 5*8-1 downto  4*8), w06 => Pw(55)( 6*8-1 downto  5*8), w07 => Pw(55)( 7*8-1 downto  6*8), w08 => Pw(55)( 8*8-1 downto  7*8),  
w09 => Pw(55)( 9*8-1 downto  8*8), w10 => Pw(55)(10*8-1 downto  9*8), w11 => Pw(55)(11*8-1 downto 10*8), w12 => Pw(55)(12*8-1 downto 11*8), w13 => Pw(55)(13*8-1 downto 12*8), w14 => Pw(55)(14*8-1 downto 13*8), w15 => Pw(55)(15*8-1 downto 14*8), w16 => Pw(55)(16*8-1 downto 15*8),  
w17 => Pw(55)(17*8-1 downto 16*8), w18 => Pw(55)(18*8-1 downto 17*8), w19 => Pw(55)(19*8-1 downto 18*8), w20 => Pw(55)(20*8-1 downto 19*8), w21 => Pw(55)(21*8-1 downto 20*8), w22 => Pw(55)(22*8-1 downto 21*8), w23 => Pw(55)(23*8-1 downto 22*8), w24 => Pw(55)(24*8-1 downto 23*8),  
w25 => Pw(55)(25*8-1 downto 24*8), w26 => Pw(55)(26*8-1 downto 25*8), w27 => Pw(55)(27*8-1 downto 26*8), w28 => Pw(55)(28*8-1 downto 27*8), w29 => Pw(55)(29*8-1 downto 28*8), w30 => Pw(55)(30*8-1 downto 29*8), w31 => Pw(55)(31*8-1 downto 30*8), w32 => Pw(55)(32*8-1 downto 31*8),  
w33 => Pw(55)(33*8-1 downto 32*8), w34 => Pw(55)(34*8-1 downto 33*8), w35 => Pw(55)(35*8-1 downto 34*8), w36 => Pw(55)(36*8-1 downto 35*8), w37 => Pw(55)(37*8-1 downto 36*8), w38 => Pw(55)(38*8-1 downto 37*8), w39 => Pw(55)(39*8-1 downto 38*8), w40 => Pw(55)(40*8-1 downto 39*8),  
w41 => Pw(55)(41*8-1 downto 40*8), w42 => Pw(55)(42*8-1 downto 41*8), w43 => Pw(55)(43*8-1 downto 42*8), w44 => Pw(55)(44*8-1 downto 43*8), w45 => Pw(55)(45*8-1 downto 44*8), w46 => Pw(55)(46*8-1 downto 45*8), w47 => Pw(55)(47*8-1 downto 46*8), w48 => Pw(55)(48*8-1 downto 47*8),  
w49 => Pw(55)(49*8-1 downto 48*8), w50 => Pw(55)(50*8-1 downto 49*8), w51 => Pw(55)(51*8-1 downto 50*8), w52 => Pw(55)(52*8-1 downto 51*8), w53 => Pw(55)(53*8-1 downto 52*8), w54 => Pw(55)(54*8-1 downto 53*8), w55 => Pw(55)(55*8-1 downto 54*8), w56 => Pw(55)(56*8-1 downto 55*8),  
w57 => Pw(55)(57*8-1 downto 56*8), w58 => Pw(55)(58*8-1 downto 57*8), w59 => Pw(55)(59*8-1 downto 58*8), w60 => Pw(55)(60*8-1 downto 59*8), w61 => Pw(55)(61*8-1 downto 60*8), w62 => Pw(55)(62*8-1 downto 61*8), w63 => Pw(55)(63*8-1 downto 62*8), w64 => Pw(55)(64*8-1 downto 63*8), 
w65 => Pw(55)( 65*8-1 downto  64*8), w66 => Pw(55)( 66*8-1 downto  65*8), w67 => Pw(55)( 67*8-1 downto  66*8), w68 => Pw(55)( 68*8-1 downto  67*8), w69 => Pw(55)( 69*8-1 downto  68*8), w70 => Pw(55)( 70*8-1 downto  69*8), w71 => Pw(55)( 71*8-1 downto  70*8), w72 => Pw(55)( 72*8-1 downto  71*8), 
w73 => Pw(55)( 73*8-1 downto  72*8), w74 => Pw(55)( 74*8-1 downto  73*8), w75 => Pw(55)( 75*8-1 downto  74*8), w76 => Pw(55)( 76*8-1 downto  75*8), w77 => Pw(55)( 77*8-1 downto  76*8), w78 => Pw(55)( 78*8-1 downto  77*8), w79 => Pw(55)( 79*8-1 downto  78*8), w80 => Pw(55)( 80*8-1 downto  79*8), 
w81 => Pw(55)( 81*8-1 downto  80*8), w82 => Pw(55)( 82*8-1 downto  81*8), w83 => Pw(55)( 83*8-1 downto  82*8), w84 => Pw(55)( 84*8-1 downto  83*8), w85 => Pw(55)( 85*8-1 downto  84*8), w86 => Pw(55)( 86*8-1 downto  85*8), w87 => Pw(55)( 87*8-1 downto  86*8), w88 => Pw(55)( 88*8-1 downto  87*8), 
w89 => Pw(55)( 89*8-1 downto  88*8), w90 => Pw(55)( 90*8-1 downto  89*8), w91 => Pw(55)( 91*8-1 downto  90*8), w92 => Pw(55)( 92*8-1 downto  91*8), w93 => Pw(55)( 93*8-1 downto  92*8), w94 => Pw(55)( 94*8-1 downto  93*8), w95 => Pw(55)( 95*8-1 downto  94*8), w96 => Pw(55)( 96*8-1 downto  95*8), 
w97 => Pw(55)( 97*8-1 downto  96*8), w98 => Pw(55)( 98*8-1 downto  97*8), w99 => Pw(55)( 99*8-1 downto  98*8), w100=> Pw(55)(100*8-1 downto  99*8), w101=> Pw(55)(101*8-1 downto 100*8), w102=> Pw(55)(102*8-1 downto 101*8), w103=> Pw(55)(103*8-1 downto 102*8), w104=> Pw(55)(104*8-1 downto 103*8), 
w105=> Pw(55)(105*8-1 downto 104*8), w106=> Pw(55)(106*8-1 downto 105*8), w107=> Pw(55)(107*8-1 downto 106*8), w108=> Pw(55)(108*8-1 downto 107*8), w109=> Pw(55)(109*8-1 downto 108*8), w110=> Pw(55)(110*8-1 downto 109*8), w111=> Pw(55)(111*8-1 downto 110*8), w112=> Pw(55)(112*8-1 downto 111*8), 
w113=> Pw(55)(113*8-1 downto 112*8), w114=> Pw(55)(114*8-1 downto 113*8), w115=> Pw(55)(115*8-1 downto 114*8), w116=> Pw(55)(116*8-1 downto 115*8), w117=> Pw(55)(117*8-1 downto 116*8), w118=> Pw(55)(118*8-1 downto 117*8), w119=> Pw(55)(119*8-1 downto 118*8), w120=> Pw(55)(120*8-1 downto 119*8), 
w121=> Pw(55)(121*8-1 downto 120*8), w122=> Pw(55)(122*8-1 downto 121*8), w123=> Pw(55)(123*8-1 downto 122*8), w124=> Pw(55)(124*8-1 downto 123*8), w125=> Pw(55)(125*8-1 downto 124*8), w126=> Pw(55)(126*8-1 downto 125*8), w127=> Pw(55)(127*8-1 downto 126*8), w128=> Pw(55)(128*8-1 downto 127*8), 

           d_out   => pca_d55_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_56_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(56)(     7 downto    0), w02 => Pw(56)( 2*8-1 downto    8), w03 => Pw(56)( 3*8-1 downto  2*8), w04 => Pw(56)( 4*8-1 downto  3*8), w05 => Pw(56)( 5*8-1 downto  4*8), w06 => Pw(56)( 6*8-1 downto  5*8), w07 => Pw(56)( 7*8-1 downto  6*8), w08 => Pw(56)( 8*8-1 downto  7*8),  
w09 => Pw(56)( 9*8-1 downto  8*8), w10 => Pw(56)(10*8-1 downto  9*8), w11 => Pw(56)(11*8-1 downto 10*8), w12 => Pw(56)(12*8-1 downto 11*8), w13 => Pw(56)(13*8-1 downto 12*8), w14 => Pw(56)(14*8-1 downto 13*8), w15 => Pw(56)(15*8-1 downto 14*8), w16 => Pw(56)(16*8-1 downto 15*8),  
w17 => Pw(56)(17*8-1 downto 16*8), w18 => Pw(56)(18*8-1 downto 17*8), w19 => Pw(56)(19*8-1 downto 18*8), w20 => Pw(56)(20*8-1 downto 19*8), w21 => Pw(56)(21*8-1 downto 20*8), w22 => Pw(56)(22*8-1 downto 21*8), w23 => Pw(56)(23*8-1 downto 22*8), w24 => Pw(56)(24*8-1 downto 23*8),  
w25 => Pw(56)(25*8-1 downto 24*8), w26 => Pw(56)(26*8-1 downto 25*8), w27 => Pw(56)(27*8-1 downto 26*8), w28 => Pw(56)(28*8-1 downto 27*8), w29 => Pw(56)(29*8-1 downto 28*8), w30 => Pw(56)(30*8-1 downto 29*8), w31 => Pw(56)(31*8-1 downto 30*8), w32 => Pw(56)(32*8-1 downto 31*8),  
w33 => Pw(56)(33*8-1 downto 32*8), w34 => Pw(56)(34*8-1 downto 33*8), w35 => Pw(56)(35*8-1 downto 34*8), w36 => Pw(56)(36*8-1 downto 35*8), w37 => Pw(56)(37*8-1 downto 36*8), w38 => Pw(56)(38*8-1 downto 37*8), w39 => Pw(56)(39*8-1 downto 38*8), w40 => Pw(56)(40*8-1 downto 39*8),  
w41 => Pw(56)(41*8-1 downto 40*8), w42 => Pw(56)(42*8-1 downto 41*8), w43 => Pw(56)(43*8-1 downto 42*8), w44 => Pw(56)(44*8-1 downto 43*8), w45 => Pw(56)(45*8-1 downto 44*8), w46 => Pw(56)(46*8-1 downto 45*8), w47 => Pw(56)(47*8-1 downto 46*8), w48 => Pw(56)(48*8-1 downto 47*8),  
w49 => Pw(56)(49*8-1 downto 48*8), w50 => Pw(56)(50*8-1 downto 49*8), w51 => Pw(56)(51*8-1 downto 50*8), w52 => Pw(56)(52*8-1 downto 51*8), w53 => Pw(56)(53*8-1 downto 52*8), w54 => Pw(56)(54*8-1 downto 53*8), w55 => Pw(56)(55*8-1 downto 54*8), w56 => Pw(56)(56*8-1 downto 55*8),  
w57 => Pw(56)(57*8-1 downto 56*8), w58 => Pw(56)(58*8-1 downto 57*8), w59 => Pw(56)(59*8-1 downto 58*8), w60 => Pw(56)(60*8-1 downto 59*8), w61 => Pw(56)(61*8-1 downto 60*8), w62 => Pw(56)(62*8-1 downto 61*8), w63 => Pw(56)(63*8-1 downto 62*8), w64 => Pw(56)(64*8-1 downto 63*8), 
w65 => Pw(56)( 65*8-1 downto  64*8), w66 => Pw(56)( 66*8-1 downto  65*8), w67 => Pw(56)( 67*8-1 downto  66*8), w68 => Pw(56)( 68*8-1 downto  67*8), w69 => Pw(56)( 69*8-1 downto  68*8), w70 => Pw(56)( 70*8-1 downto  69*8), w71 => Pw(56)( 71*8-1 downto  70*8), w72 => Pw(56)( 72*8-1 downto  71*8), 
w73 => Pw(56)( 73*8-1 downto  72*8), w74 => Pw(56)( 74*8-1 downto  73*8), w75 => Pw(56)( 75*8-1 downto  74*8), w76 => Pw(56)( 76*8-1 downto  75*8), w77 => Pw(56)( 77*8-1 downto  76*8), w78 => Pw(56)( 78*8-1 downto  77*8), w79 => Pw(56)( 79*8-1 downto  78*8), w80 => Pw(56)( 80*8-1 downto  79*8), 
w81 => Pw(56)( 81*8-1 downto  80*8), w82 => Pw(56)( 82*8-1 downto  81*8), w83 => Pw(56)( 83*8-1 downto  82*8), w84 => Pw(56)( 84*8-1 downto  83*8), w85 => Pw(56)( 85*8-1 downto  84*8), w86 => Pw(56)( 86*8-1 downto  85*8), w87 => Pw(56)( 87*8-1 downto  86*8), w88 => Pw(56)( 88*8-1 downto  87*8), 
w89 => Pw(56)( 89*8-1 downto  88*8), w90 => Pw(56)( 90*8-1 downto  89*8), w91 => Pw(56)( 91*8-1 downto  90*8), w92 => Pw(56)( 92*8-1 downto  91*8), w93 => Pw(56)( 93*8-1 downto  92*8), w94 => Pw(56)( 94*8-1 downto  93*8), w95 => Pw(56)( 95*8-1 downto  94*8), w96 => Pw(56)( 96*8-1 downto  95*8), 
w97 => Pw(56)( 97*8-1 downto  96*8), w98 => Pw(56)( 98*8-1 downto  97*8), w99 => Pw(56)( 99*8-1 downto  98*8), w100=> Pw(56)(100*8-1 downto  99*8), w101=> Pw(56)(101*8-1 downto 100*8), w102=> Pw(56)(102*8-1 downto 101*8), w103=> Pw(56)(103*8-1 downto 102*8), w104=> Pw(56)(104*8-1 downto 103*8), 
w105=> Pw(56)(105*8-1 downto 104*8), w106=> Pw(56)(106*8-1 downto 105*8), w107=> Pw(56)(107*8-1 downto 106*8), w108=> Pw(56)(108*8-1 downto 107*8), w109=> Pw(56)(109*8-1 downto 108*8), w110=> Pw(56)(110*8-1 downto 109*8), w111=> Pw(56)(111*8-1 downto 110*8), w112=> Pw(56)(112*8-1 downto 111*8), 
w113=> Pw(56)(113*8-1 downto 112*8), w114=> Pw(56)(114*8-1 downto 113*8), w115=> Pw(56)(115*8-1 downto 114*8), w116=> Pw(56)(116*8-1 downto 115*8), w117=> Pw(56)(117*8-1 downto 116*8), w118=> Pw(56)(118*8-1 downto 117*8), w119=> Pw(56)(119*8-1 downto 118*8), w120=> Pw(56)(120*8-1 downto 119*8), 
w121=> Pw(56)(121*8-1 downto 120*8), w122=> Pw(56)(122*8-1 downto 121*8), w123=> Pw(56)(123*8-1 downto 122*8), w124=> Pw(56)(124*8-1 downto 123*8), w125=> Pw(56)(125*8-1 downto 124*8), w126=> Pw(56)(126*8-1 downto 125*8), w127=> Pw(56)(127*8-1 downto 126*8), w128=> Pw(56)(128*8-1 downto 127*8), 

           d_out   => pca_d56_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_57_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out, 

w01 => Pw(57)(     7 downto    0), w02 => Pw(57)( 2*8-1 downto    8), w03 => Pw(57)( 3*8-1 downto  2*8), w04 => Pw(57)( 4*8-1 downto  3*8), w05 => Pw(57)( 5*8-1 downto  4*8), w06 => Pw(57)( 6*8-1 downto  5*8), w07 => Pw(57)( 7*8-1 downto  6*8), w08 => Pw(57)( 8*8-1 downto  7*8),  
w09 => Pw(57)( 9*8-1 downto  8*8), w10 => Pw(57)(10*8-1 downto  9*8), w11 => Pw(57)(11*8-1 downto 10*8), w12 => Pw(57)(12*8-1 downto 11*8), w13 => Pw(57)(13*8-1 downto 12*8), w14 => Pw(57)(14*8-1 downto 13*8), w15 => Pw(57)(15*8-1 downto 14*8), w16 => Pw(57)(16*8-1 downto 15*8),  
w17 => Pw(57)(17*8-1 downto 16*8), w18 => Pw(57)(18*8-1 downto 17*8), w19 => Pw(57)(19*8-1 downto 18*8), w20 => Pw(57)(20*8-1 downto 19*8), w21 => Pw(57)(21*8-1 downto 20*8), w22 => Pw(57)(22*8-1 downto 21*8), w23 => Pw(57)(23*8-1 downto 22*8), w24 => Pw(57)(24*8-1 downto 23*8),  
w25 => Pw(57)(25*8-1 downto 24*8), w26 => Pw(57)(26*8-1 downto 25*8), w27 => Pw(57)(27*8-1 downto 26*8), w28 => Pw(57)(28*8-1 downto 27*8), w29 => Pw(57)(29*8-1 downto 28*8), w30 => Pw(57)(30*8-1 downto 29*8), w31 => Pw(57)(31*8-1 downto 30*8), w32 => Pw(57)(32*8-1 downto 31*8),  
w33 => Pw(57)(33*8-1 downto 32*8), w34 => Pw(57)(34*8-1 downto 33*8), w35 => Pw(57)(35*8-1 downto 34*8), w36 => Pw(57)(36*8-1 downto 35*8), w37 => Pw(57)(37*8-1 downto 36*8), w38 => Pw(57)(38*8-1 downto 37*8), w39 => Pw(57)(39*8-1 downto 38*8), w40 => Pw(57)(40*8-1 downto 39*8),  
w41 => Pw(57)(41*8-1 downto 40*8), w42 => Pw(57)(42*8-1 downto 41*8), w43 => Pw(57)(43*8-1 downto 42*8), w44 => Pw(57)(44*8-1 downto 43*8), w45 => Pw(57)(45*8-1 downto 44*8), w46 => Pw(57)(46*8-1 downto 45*8), w47 => Pw(57)(47*8-1 downto 46*8), w48 => Pw(57)(48*8-1 downto 47*8),  
w49 => Pw(57)(49*8-1 downto 48*8), w50 => Pw(57)(50*8-1 downto 49*8), w51 => Pw(57)(51*8-1 downto 50*8), w52 => Pw(57)(52*8-1 downto 51*8), w53 => Pw(57)(53*8-1 downto 52*8), w54 => Pw(57)(54*8-1 downto 53*8), w55 => Pw(57)(55*8-1 downto 54*8), w56 => Pw(57)(56*8-1 downto 55*8),  
w57 => Pw(57)(57*8-1 downto 56*8), w58 => Pw(57)(58*8-1 downto 57*8), w59 => Pw(57)(59*8-1 downto 58*8), w60 => Pw(57)(60*8-1 downto 59*8), w61 => Pw(57)(61*8-1 downto 60*8), w62 => Pw(57)(62*8-1 downto 61*8), w63 => Pw(57)(63*8-1 downto 62*8), w64 => Pw(57)(64*8-1 downto 63*8), 
w65 => Pw(57)( 65*8-1 downto  64*8), w66 => Pw(57)( 66*8-1 downto  65*8), w67 => Pw(57)( 67*8-1 downto  66*8), w68 => Pw(57)( 68*8-1 downto  67*8), w69 => Pw(57)( 69*8-1 downto  68*8), w70 => Pw(57)( 70*8-1 downto  69*8), w71 => Pw(57)( 71*8-1 downto  70*8), w72 => Pw(57)( 72*8-1 downto  71*8), 
w73 => Pw(57)( 73*8-1 downto  72*8), w74 => Pw(57)( 74*8-1 downto  73*8), w75 => Pw(57)( 75*8-1 downto  74*8), w76 => Pw(57)( 76*8-1 downto  75*8), w77 => Pw(57)( 77*8-1 downto  76*8), w78 => Pw(57)( 78*8-1 downto  77*8), w79 => Pw(57)( 79*8-1 downto  78*8), w80 => Pw(57)( 80*8-1 downto  79*8), 
w81 => Pw(57)( 81*8-1 downto  80*8), w82 => Pw(57)( 82*8-1 downto  81*8), w83 => Pw(57)( 83*8-1 downto  82*8), w84 => Pw(57)( 84*8-1 downto  83*8), w85 => Pw(57)( 85*8-1 downto  84*8), w86 => Pw(57)( 86*8-1 downto  85*8), w87 => Pw(57)( 87*8-1 downto  86*8), w88 => Pw(57)( 88*8-1 downto  87*8), 
w89 => Pw(57)( 89*8-1 downto  88*8), w90 => Pw(57)( 90*8-1 downto  89*8), w91 => Pw(57)( 91*8-1 downto  90*8), w92 => Pw(57)( 92*8-1 downto  91*8), w93 => Pw(57)( 93*8-1 downto  92*8), w94 => Pw(57)( 94*8-1 downto  93*8), w95 => Pw(57)( 95*8-1 downto  94*8), w96 => Pw(57)( 96*8-1 downto  95*8), 
w97 => Pw(57)( 97*8-1 downto  96*8), w98 => Pw(57)( 98*8-1 downto  97*8), w99 => Pw(57)( 99*8-1 downto  98*8), w100=> Pw(57)(100*8-1 downto  99*8), w101=> Pw(57)(101*8-1 downto 100*8), w102=> Pw(57)(102*8-1 downto 101*8), w103=> Pw(57)(103*8-1 downto 102*8), w104=> Pw(57)(104*8-1 downto 103*8), 
w105=> Pw(57)(105*8-1 downto 104*8), w106=> Pw(57)(106*8-1 downto 105*8), w107=> Pw(57)(107*8-1 downto 106*8), w108=> Pw(57)(108*8-1 downto 107*8), w109=> Pw(57)(109*8-1 downto 108*8), w110=> Pw(57)(110*8-1 downto 109*8), w111=> Pw(57)(111*8-1 downto 110*8), w112=> Pw(57)(112*8-1 downto 111*8), 
w113=> Pw(57)(113*8-1 downto 112*8), w114=> Pw(57)(114*8-1 downto 113*8), w115=> Pw(57)(115*8-1 downto 114*8), w116=> Pw(57)(116*8-1 downto 115*8), w117=> Pw(57)(117*8-1 downto 116*8), w118=> Pw(57)(118*8-1 downto 117*8), w119=> Pw(57)(119*8-1 downto 118*8), w120=> Pw(57)(120*8-1 downto 119*8), 
w121=> Pw(57)(121*8-1 downto 120*8), w122=> Pw(57)(122*8-1 downto 121*8), w123=> Pw(57)(123*8-1 downto 122*8), w124=> Pw(57)(124*8-1 downto 123*8), w125=> Pw(57)(125*8-1 downto 124*8), w126=> Pw(57)(126*8-1 downto 125*8), w127=> Pw(57)(127*8-1 downto 126*8), w128=> Pw(57)(128*8-1 downto 127*8), 

           d_out   => pca_d57_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_58_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out, 

w01 => Pw(58)(     7 downto    0), w02 => Pw(58)( 2*8-1 downto    8), w03 => Pw(58)( 3*8-1 downto  2*8), w04 => Pw(58)( 4*8-1 downto  3*8), w05 => Pw(58)( 5*8-1 downto  4*8), w06 => Pw(58)( 6*8-1 downto  5*8), w07 => Pw(58)( 7*8-1 downto  6*8), w08 => Pw(58)( 8*8-1 downto  7*8),  
w09 => Pw(58)( 9*8-1 downto  8*8), w10 => Pw(58)(10*8-1 downto  9*8), w11 => Pw(58)(11*8-1 downto 10*8), w12 => Pw(58)(12*8-1 downto 11*8), w13 => Pw(58)(13*8-1 downto 12*8), w14 => Pw(58)(14*8-1 downto 13*8), w15 => Pw(58)(15*8-1 downto 14*8), w16 => Pw(58)(16*8-1 downto 15*8),  
w17 => Pw(58)(17*8-1 downto 16*8), w18 => Pw(58)(18*8-1 downto 17*8), w19 => Pw(58)(19*8-1 downto 18*8), w20 => Pw(58)(20*8-1 downto 19*8), w21 => Pw(58)(21*8-1 downto 20*8), w22 => Pw(58)(22*8-1 downto 21*8), w23 => Pw(58)(23*8-1 downto 22*8), w24 => Pw(58)(24*8-1 downto 23*8),  
w25 => Pw(58)(25*8-1 downto 24*8), w26 => Pw(58)(26*8-1 downto 25*8), w27 => Pw(58)(27*8-1 downto 26*8), w28 => Pw(58)(28*8-1 downto 27*8), w29 => Pw(58)(29*8-1 downto 28*8), w30 => Pw(58)(30*8-1 downto 29*8), w31 => Pw(58)(31*8-1 downto 30*8), w32 => Pw(58)(32*8-1 downto 31*8),  
w33 => Pw(58)(33*8-1 downto 32*8), w34 => Pw(58)(34*8-1 downto 33*8), w35 => Pw(58)(35*8-1 downto 34*8), w36 => Pw(58)(36*8-1 downto 35*8), w37 => Pw(58)(37*8-1 downto 36*8), w38 => Pw(58)(38*8-1 downto 37*8), w39 => Pw(58)(39*8-1 downto 38*8), w40 => Pw(58)(40*8-1 downto 39*8),  
w41 => Pw(58)(41*8-1 downto 40*8), w42 => Pw(58)(42*8-1 downto 41*8), w43 => Pw(58)(43*8-1 downto 42*8), w44 => Pw(58)(44*8-1 downto 43*8), w45 => Pw(58)(45*8-1 downto 44*8), w46 => Pw(58)(46*8-1 downto 45*8), w47 => Pw(58)(47*8-1 downto 46*8), w48 => Pw(58)(48*8-1 downto 47*8),  
w49 => Pw(58)(49*8-1 downto 48*8), w50 => Pw(58)(50*8-1 downto 49*8), w51 => Pw(58)(51*8-1 downto 50*8), w52 => Pw(58)(52*8-1 downto 51*8), w53 => Pw(58)(53*8-1 downto 52*8), w54 => Pw(58)(54*8-1 downto 53*8), w55 => Pw(58)(55*8-1 downto 54*8), w56 => Pw(58)(56*8-1 downto 55*8),  
w57 => Pw(58)(57*8-1 downto 56*8), w58 => Pw(58)(58*8-1 downto 57*8), w59 => Pw(58)(59*8-1 downto 58*8), w60 => Pw(58)(60*8-1 downto 59*8), w61 => Pw(58)(61*8-1 downto 60*8), w62 => Pw(58)(62*8-1 downto 61*8), w63 => Pw(58)(63*8-1 downto 62*8), w64 => Pw(58)(64*8-1 downto 63*8), 
w65 => Pw(58)( 65*8-1 downto  64*8), w66 => Pw(58)( 66*8-1 downto  65*8), w67 => Pw(58)( 67*8-1 downto  66*8), w68 => Pw(58)( 68*8-1 downto  67*8), w69 => Pw(58)( 69*8-1 downto  68*8), w70 => Pw(58)( 70*8-1 downto  69*8), w71 => Pw(58)( 71*8-1 downto  70*8), w72 => Pw(58)( 72*8-1 downto  71*8), 
w73 => Pw(58)( 73*8-1 downto  72*8), w74 => Pw(58)( 74*8-1 downto  73*8), w75 => Pw(58)( 75*8-1 downto  74*8), w76 => Pw(58)( 76*8-1 downto  75*8), w77 => Pw(58)( 77*8-1 downto  76*8), w78 => Pw(58)( 78*8-1 downto  77*8), w79 => Pw(58)( 79*8-1 downto  78*8), w80 => Pw(58)( 80*8-1 downto  79*8), 
w81 => Pw(58)( 81*8-1 downto  80*8), w82 => Pw(58)( 82*8-1 downto  81*8), w83 => Pw(58)( 83*8-1 downto  82*8), w84 => Pw(58)( 84*8-1 downto  83*8), w85 => Pw(58)( 85*8-1 downto  84*8), w86 => Pw(58)( 86*8-1 downto  85*8), w87 => Pw(58)( 87*8-1 downto  86*8), w88 => Pw(58)( 88*8-1 downto  87*8), 
w89 => Pw(58)( 89*8-1 downto  88*8), w90 => Pw(58)( 90*8-1 downto  89*8), w91 => Pw(58)( 91*8-1 downto  90*8), w92 => Pw(58)( 92*8-1 downto  91*8), w93 => Pw(58)( 93*8-1 downto  92*8), w94 => Pw(58)( 94*8-1 downto  93*8), w95 => Pw(58)( 95*8-1 downto  94*8), w96 => Pw(58)( 96*8-1 downto  95*8), 
w97 => Pw(58)( 97*8-1 downto  96*8), w98 => Pw(58)( 98*8-1 downto  97*8), w99 => Pw(58)( 99*8-1 downto  98*8), w100=> Pw(58)(100*8-1 downto  99*8), w101=> Pw(58)(101*8-1 downto 100*8), w102=> Pw(58)(102*8-1 downto 101*8), w103=> Pw(58)(103*8-1 downto 102*8), w104=> Pw(58)(104*8-1 downto 103*8), 
w105=> Pw(58)(105*8-1 downto 104*8), w106=> Pw(58)(106*8-1 downto 105*8), w107=> Pw(58)(107*8-1 downto 106*8), w108=> Pw(58)(108*8-1 downto 107*8), w109=> Pw(58)(109*8-1 downto 108*8), w110=> Pw(58)(110*8-1 downto 109*8), w111=> Pw(58)(111*8-1 downto 110*8), w112=> Pw(58)(112*8-1 downto 111*8), 
w113=> Pw(58)(113*8-1 downto 112*8), w114=> Pw(58)(114*8-1 downto 113*8), w115=> Pw(58)(115*8-1 downto 114*8), w116=> Pw(58)(116*8-1 downto 115*8), w117=> Pw(58)(117*8-1 downto 116*8), w118=> Pw(58)(118*8-1 downto 117*8), w119=> Pw(58)(119*8-1 downto 118*8), w120=> Pw(58)(120*8-1 downto 119*8), 
w121=> Pw(58)(121*8-1 downto 120*8), w122=> Pw(58)(122*8-1 downto 121*8), w123=> Pw(58)(123*8-1 downto 122*8), w124=> Pw(58)(124*8-1 downto 123*8), w125=> Pw(58)(125*8-1 downto 124*8), w126=> Pw(58)(126*8-1 downto 125*8), w127=> Pw(58)(127*8-1 downto 126*8), w128=> Pw(58)(128*8-1 downto 127*8), 

           d_out   => pca_d58_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_59_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(59)(     7 downto    0), w02 => Pw(59)( 2*8-1 downto    8), w03 => Pw(59)( 3*8-1 downto  2*8), w04 => Pw(59)( 4*8-1 downto  3*8), w05 => Pw(59)( 5*8-1 downto  4*8), w06 => Pw(59)( 6*8-1 downto  5*8), w07 => Pw(59)( 7*8-1 downto  6*8), w08 => Pw(59)( 8*8-1 downto  7*8),  
w09 => Pw(59)( 9*8-1 downto  8*8), w10 => Pw(59)(10*8-1 downto  9*8), w11 => Pw(59)(11*8-1 downto 10*8), w12 => Pw(59)(12*8-1 downto 11*8), w13 => Pw(59)(13*8-1 downto 12*8), w14 => Pw(59)(14*8-1 downto 13*8), w15 => Pw(59)(15*8-1 downto 14*8), w16 => Pw(59)(16*8-1 downto 15*8),  
w17 => Pw(59)(17*8-1 downto 16*8), w18 => Pw(59)(18*8-1 downto 17*8), w19 => Pw(59)(19*8-1 downto 18*8), w20 => Pw(59)(20*8-1 downto 19*8), w21 => Pw(59)(21*8-1 downto 20*8), w22 => Pw(59)(22*8-1 downto 21*8), w23 => Pw(59)(23*8-1 downto 22*8), w24 => Pw(59)(24*8-1 downto 23*8),  
w25 => Pw(59)(25*8-1 downto 24*8), w26 => Pw(59)(26*8-1 downto 25*8), w27 => Pw(59)(27*8-1 downto 26*8), w28 => Pw(59)(28*8-1 downto 27*8), w29 => Pw(59)(29*8-1 downto 28*8), w30 => Pw(59)(30*8-1 downto 29*8), w31 => Pw(59)(31*8-1 downto 30*8), w32 => Pw(59)(32*8-1 downto 31*8),  
w33 => Pw(59)(33*8-1 downto 32*8), w34 => Pw(59)(34*8-1 downto 33*8), w35 => Pw(59)(35*8-1 downto 34*8), w36 => Pw(59)(36*8-1 downto 35*8), w37 => Pw(59)(37*8-1 downto 36*8), w38 => Pw(59)(38*8-1 downto 37*8), w39 => Pw(59)(39*8-1 downto 38*8), w40 => Pw(59)(40*8-1 downto 39*8),  
w41 => Pw(59)(41*8-1 downto 40*8), w42 => Pw(59)(42*8-1 downto 41*8), w43 => Pw(59)(43*8-1 downto 42*8), w44 => Pw(59)(44*8-1 downto 43*8), w45 => Pw(59)(45*8-1 downto 44*8), w46 => Pw(59)(46*8-1 downto 45*8), w47 => Pw(59)(47*8-1 downto 46*8), w48 => Pw(59)(48*8-1 downto 47*8),  
w49 => Pw(59)(49*8-1 downto 48*8), w50 => Pw(59)(50*8-1 downto 49*8), w51 => Pw(59)(51*8-1 downto 50*8), w52 => Pw(59)(52*8-1 downto 51*8), w53 => Pw(59)(53*8-1 downto 52*8), w54 => Pw(59)(54*8-1 downto 53*8), w55 => Pw(59)(55*8-1 downto 54*8), w56 => Pw(59)(56*8-1 downto 55*8),  
w57 => Pw(59)(57*8-1 downto 56*8), w58 => Pw(59)(58*8-1 downto 57*8), w59 => Pw(59)(59*8-1 downto 58*8), w60 => Pw(59)(60*8-1 downto 59*8), w61 => Pw(59)(61*8-1 downto 60*8), w62 => Pw(59)(62*8-1 downto 61*8), w63 => Pw(59)(63*8-1 downto 62*8), w64 => Pw(59)(64*8-1 downto 63*8), 
w65 => Pw(59)( 65*8-1 downto  64*8), w66 => Pw(59)( 66*8-1 downto  65*8), w67 => Pw(59)( 67*8-1 downto  66*8), w68 => Pw(59)( 68*8-1 downto  67*8), w69 => Pw(59)( 69*8-1 downto  68*8), w70 => Pw(59)( 70*8-1 downto  69*8), w71 => Pw(59)( 71*8-1 downto  70*8), w72 => Pw(59)( 72*8-1 downto  71*8), 
w73 => Pw(59)( 73*8-1 downto  72*8), w74 => Pw(59)( 74*8-1 downto  73*8), w75 => Pw(59)( 75*8-1 downto  74*8), w76 => Pw(59)( 76*8-1 downto  75*8), w77 => Pw(59)( 77*8-1 downto  76*8), w78 => Pw(59)( 78*8-1 downto  77*8), w79 => Pw(59)( 79*8-1 downto  78*8), w80 => Pw(59)( 80*8-1 downto  79*8), 
w81 => Pw(59)( 81*8-1 downto  80*8), w82 => Pw(59)( 82*8-1 downto  81*8), w83 => Pw(59)( 83*8-1 downto  82*8), w84 => Pw(59)( 84*8-1 downto  83*8), w85 => Pw(59)( 85*8-1 downto  84*8), w86 => Pw(59)( 86*8-1 downto  85*8), w87 => Pw(59)( 87*8-1 downto  86*8), w88 => Pw(59)( 88*8-1 downto  87*8), 
w89 => Pw(59)( 89*8-1 downto  88*8), w90 => Pw(59)( 90*8-1 downto  89*8), w91 => Pw(59)( 91*8-1 downto  90*8), w92 => Pw(59)( 92*8-1 downto  91*8), w93 => Pw(59)( 93*8-1 downto  92*8), w94 => Pw(59)( 94*8-1 downto  93*8), w95 => Pw(59)( 95*8-1 downto  94*8), w96 => Pw(59)( 96*8-1 downto  95*8), 
w97 => Pw(59)( 97*8-1 downto  96*8), w98 => Pw(59)( 98*8-1 downto  97*8), w99 => Pw(59)( 99*8-1 downto  98*8), w100=> Pw(59)(100*8-1 downto  99*8), w101=> Pw(59)(101*8-1 downto 100*8), w102=> Pw(59)(102*8-1 downto 101*8), w103=> Pw(59)(103*8-1 downto 102*8), w104=> Pw(59)(104*8-1 downto 103*8), 
w105=> Pw(59)(105*8-1 downto 104*8), w106=> Pw(59)(106*8-1 downto 105*8), w107=> Pw(59)(107*8-1 downto 106*8), w108=> Pw(59)(108*8-1 downto 107*8), w109=> Pw(59)(109*8-1 downto 108*8), w110=> Pw(59)(110*8-1 downto 109*8), w111=> Pw(59)(111*8-1 downto 110*8), w112=> Pw(59)(112*8-1 downto 111*8), 
w113=> Pw(59)(113*8-1 downto 112*8), w114=> Pw(59)(114*8-1 downto 113*8), w115=> Pw(59)(115*8-1 downto 114*8), w116=> Pw(59)(116*8-1 downto 115*8), w117=> Pw(59)(117*8-1 downto 116*8), w118=> Pw(59)(118*8-1 downto 117*8), w119=> Pw(59)(119*8-1 downto 118*8), w120=> Pw(59)(120*8-1 downto 119*8), 
w121=> Pw(59)(121*8-1 downto 120*8), w122=> Pw(59)(122*8-1 downto 121*8), w123=> Pw(59)(123*8-1 downto 122*8), w124=> Pw(59)(124*8-1 downto 123*8), w125=> Pw(59)(125*8-1 downto 124*8), w126=> Pw(59)(126*8-1 downto 125*8), w127=> Pw(59)(127*8-1 downto 126*8), w128=> Pw(59)(128*8-1 downto 127*8), 

           d_out   => pca_d59_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_60_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(60)(     7 downto    0), w02 => Pw(60)( 2*8-1 downto    8), w03 => Pw(60)( 3*8-1 downto  2*8), w04 => Pw(60)( 4*8-1 downto  3*8), w05 => Pw(60)( 5*8-1 downto  4*8), w06 => Pw(60)( 6*8-1 downto  5*8), w07 => Pw(60)( 7*8-1 downto  6*8), w08 => Pw(60)( 8*8-1 downto  7*8),  
w09 => Pw(60)( 9*8-1 downto  8*8), w10 => Pw(60)(10*8-1 downto  9*8), w11 => Pw(60)(11*8-1 downto 10*8), w12 => Pw(60)(12*8-1 downto 11*8), w13 => Pw(60)(13*8-1 downto 12*8), w14 => Pw(60)(14*8-1 downto 13*8), w15 => Pw(60)(15*8-1 downto 14*8), w16 => Pw(60)(16*8-1 downto 15*8),  
w17 => Pw(60)(17*8-1 downto 16*8), w18 => Pw(60)(18*8-1 downto 17*8), w19 => Pw(60)(19*8-1 downto 18*8), w20 => Pw(60)(20*8-1 downto 19*8), w21 => Pw(60)(21*8-1 downto 20*8), w22 => Pw(60)(22*8-1 downto 21*8), w23 => Pw(60)(23*8-1 downto 22*8), w24 => Pw(60)(24*8-1 downto 23*8),  
w25 => Pw(60)(25*8-1 downto 24*8), w26 => Pw(60)(26*8-1 downto 25*8), w27 => Pw(60)(27*8-1 downto 26*8), w28 => Pw(60)(28*8-1 downto 27*8), w29 => Pw(60)(29*8-1 downto 28*8), w30 => Pw(60)(30*8-1 downto 29*8), w31 => Pw(60)(31*8-1 downto 30*8), w32 => Pw(60)(32*8-1 downto 31*8),  
w33 => Pw(60)(33*8-1 downto 32*8), w34 => Pw(60)(34*8-1 downto 33*8), w35 => Pw(60)(35*8-1 downto 34*8), w36 => Pw(60)(36*8-1 downto 35*8), w37 => Pw(60)(37*8-1 downto 36*8), w38 => Pw(60)(38*8-1 downto 37*8), w39 => Pw(60)(39*8-1 downto 38*8), w40 => Pw(60)(40*8-1 downto 39*8),  
w41 => Pw(60)(41*8-1 downto 40*8), w42 => Pw(60)(42*8-1 downto 41*8), w43 => Pw(60)(43*8-1 downto 42*8), w44 => Pw(60)(44*8-1 downto 43*8), w45 => Pw(60)(45*8-1 downto 44*8), w46 => Pw(60)(46*8-1 downto 45*8), w47 => Pw(60)(47*8-1 downto 46*8), w48 => Pw(60)(48*8-1 downto 47*8),  
w49 => Pw(60)(49*8-1 downto 48*8), w50 => Pw(60)(50*8-1 downto 49*8), w51 => Pw(60)(51*8-1 downto 50*8), w52 => Pw(60)(52*8-1 downto 51*8), w53 => Pw(60)(53*8-1 downto 52*8), w54 => Pw(60)(54*8-1 downto 53*8), w55 => Pw(60)(55*8-1 downto 54*8), w56 => Pw(60)(56*8-1 downto 55*8),  
w57 => Pw(60)(57*8-1 downto 56*8), w58 => Pw(60)(58*8-1 downto 57*8), w59 => Pw(60)(59*8-1 downto 58*8), w60 => Pw(60)(60*8-1 downto 59*8), w61 => Pw(60)(61*8-1 downto 60*8), w62 => Pw(60)(62*8-1 downto 61*8), w63 => Pw(60)(63*8-1 downto 62*8), w64 => Pw(60)(64*8-1 downto 63*8), 
w65 => Pw(60)( 65*8-1 downto  64*8), w66 => Pw(60)( 66*8-1 downto  65*8), w67 => Pw(60)( 67*8-1 downto  66*8), w68 => Pw(60)( 68*8-1 downto  67*8), w69 => Pw(60)( 69*8-1 downto  68*8), w70 => Pw(60)( 70*8-1 downto  69*8), w71 => Pw(60)( 71*8-1 downto  70*8), w72 => Pw(60)( 72*8-1 downto  71*8), 
w73 => Pw(60)( 73*8-1 downto  72*8), w74 => Pw(60)( 74*8-1 downto  73*8), w75 => Pw(60)( 75*8-1 downto  74*8), w76 => Pw(60)( 76*8-1 downto  75*8), w77 => Pw(60)( 77*8-1 downto  76*8), w78 => Pw(60)( 78*8-1 downto  77*8), w79 => Pw(60)( 79*8-1 downto  78*8), w80 => Pw(60)( 80*8-1 downto  79*8), 
w81 => Pw(60)( 81*8-1 downto  80*8), w82 => Pw(60)( 82*8-1 downto  81*8), w83 => Pw(60)( 83*8-1 downto  82*8), w84 => Pw(60)( 84*8-1 downto  83*8), w85 => Pw(60)( 85*8-1 downto  84*8), w86 => Pw(60)( 86*8-1 downto  85*8), w87 => Pw(60)( 87*8-1 downto  86*8), w88 => Pw(60)( 88*8-1 downto  87*8), 
w89 => Pw(60)( 89*8-1 downto  88*8), w90 => Pw(60)( 90*8-1 downto  89*8), w91 => Pw(60)( 91*8-1 downto  90*8), w92 => Pw(60)( 92*8-1 downto  91*8), w93 => Pw(60)( 93*8-1 downto  92*8), w94 => Pw(60)( 94*8-1 downto  93*8), w95 => Pw(60)( 95*8-1 downto  94*8), w96 => Pw(60)( 96*8-1 downto  95*8), 
w97 => Pw(60)( 97*8-1 downto  96*8), w98 => Pw(60)( 98*8-1 downto  97*8), w99 => Pw(60)( 99*8-1 downto  98*8), w100=> Pw(60)(100*8-1 downto  99*8), w101=> Pw(60)(101*8-1 downto 100*8), w102=> Pw(60)(102*8-1 downto 101*8), w103=> Pw(60)(103*8-1 downto 102*8), w104=> Pw(60)(104*8-1 downto 103*8), 
w105=> Pw(60)(105*8-1 downto 104*8), w106=> Pw(60)(106*8-1 downto 105*8), w107=> Pw(60)(107*8-1 downto 106*8), w108=> Pw(60)(108*8-1 downto 107*8), w109=> Pw(60)(109*8-1 downto 108*8), w110=> Pw(60)(110*8-1 downto 109*8), w111=> Pw(60)(111*8-1 downto 110*8), w112=> Pw(60)(112*8-1 downto 111*8), 
w113=> Pw(60)(113*8-1 downto 112*8), w114=> Pw(60)(114*8-1 downto 113*8), w115=> Pw(60)(115*8-1 downto 114*8), w116=> Pw(60)(116*8-1 downto 115*8), w117=> Pw(60)(117*8-1 downto 116*8), w118=> Pw(60)(118*8-1 downto 117*8), w119=> Pw(60)(119*8-1 downto 118*8), w120=> Pw(60)(120*8-1 downto 119*8), 
w121=> Pw(60)(121*8-1 downto 120*8), w122=> Pw(60)(122*8-1 downto 121*8), w123=> Pw(60)(123*8-1 downto 122*8), w124=> Pw(60)(124*8-1 downto 123*8), w125=> Pw(60)(125*8-1 downto 124*8), w126=> Pw(60)(126*8-1 downto 125*8), w127=> Pw(60)(127*8-1 downto 126*8), w128=> Pw(60)(128*8-1 downto 127*8), 

           d_out   => pca_d60_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_61_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(61)(     7 downto    0), w02 => Pw(61)( 2*8-1 downto    8), w03 => Pw(61)( 3*8-1 downto  2*8), w04 => Pw(61)( 4*8-1 downto  3*8), w05 => Pw(61)( 5*8-1 downto  4*8), w06 => Pw(61)( 6*8-1 downto  5*8), w07 => Pw(61)( 7*8-1 downto  6*8), w08 => Pw(61)( 8*8-1 downto  7*8),  
w09 => Pw(61)( 9*8-1 downto  8*8), w10 => Pw(61)(10*8-1 downto  9*8), w11 => Pw(61)(11*8-1 downto 10*8), w12 => Pw(61)(12*8-1 downto 11*8), w13 => Pw(61)(13*8-1 downto 12*8), w14 => Pw(61)(14*8-1 downto 13*8), w15 => Pw(61)(15*8-1 downto 14*8), w16 => Pw(61)(16*8-1 downto 15*8),  
w17 => Pw(61)(17*8-1 downto 16*8), w18 => Pw(61)(18*8-1 downto 17*8), w19 => Pw(61)(19*8-1 downto 18*8), w20 => Pw(61)(20*8-1 downto 19*8), w21 => Pw(61)(21*8-1 downto 20*8), w22 => Pw(61)(22*8-1 downto 21*8), w23 => Pw(61)(23*8-1 downto 22*8), w24 => Pw(61)(24*8-1 downto 23*8),  
w25 => Pw(61)(25*8-1 downto 24*8), w26 => Pw(61)(26*8-1 downto 25*8), w27 => Pw(61)(27*8-1 downto 26*8), w28 => Pw(61)(28*8-1 downto 27*8), w29 => Pw(61)(29*8-1 downto 28*8), w30 => Pw(61)(30*8-1 downto 29*8), w31 => Pw(61)(31*8-1 downto 30*8), w32 => Pw(61)(32*8-1 downto 31*8),  
w33 => Pw(61)(33*8-1 downto 32*8), w34 => Pw(61)(34*8-1 downto 33*8), w35 => Pw(61)(35*8-1 downto 34*8), w36 => Pw(61)(36*8-1 downto 35*8), w37 => Pw(61)(37*8-1 downto 36*8), w38 => Pw(61)(38*8-1 downto 37*8), w39 => Pw(61)(39*8-1 downto 38*8), w40 => Pw(61)(40*8-1 downto 39*8),  
w41 => Pw(61)(41*8-1 downto 40*8), w42 => Pw(61)(42*8-1 downto 41*8), w43 => Pw(61)(43*8-1 downto 42*8), w44 => Pw(61)(44*8-1 downto 43*8), w45 => Pw(61)(45*8-1 downto 44*8), w46 => Pw(61)(46*8-1 downto 45*8), w47 => Pw(61)(47*8-1 downto 46*8), w48 => Pw(61)(48*8-1 downto 47*8),  
w49 => Pw(61)(49*8-1 downto 48*8), w50 => Pw(61)(50*8-1 downto 49*8), w51 => Pw(61)(51*8-1 downto 50*8), w52 => Pw(61)(52*8-1 downto 51*8), w53 => Pw(61)(53*8-1 downto 52*8), w54 => Pw(61)(54*8-1 downto 53*8), w55 => Pw(61)(55*8-1 downto 54*8), w56 => Pw(61)(56*8-1 downto 55*8),  
w57 => Pw(61)(57*8-1 downto 56*8), w58 => Pw(61)(58*8-1 downto 57*8), w59 => Pw(61)(59*8-1 downto 58*8), w60 => Pw(61)(60*8-1 downto 59*8), w61 => Pw(61)(61*8-1 downto 60*8), w62 => Pw(61)(62*8-1 downto 61*8), w63 => Pw(61)(63*8-1 downto 62*8), w64 => Pw(61)(64*8-1 downto 63*8), 
w65 => Pw(61)( 65*8-1 downto  64*8), w66 => Pw(61)( 66*8-1 downto  65*8), w67 => Pw(61)( 67*8-1 downto  66*8), w68 => Pw(61)( 68*8-1 downto  67*8), w69 => Pw(61)( 69*8-1 downto  68*8), w70 => Pw(61)( 70*8-1 downto  69*8), w71 => Pw(61)( 71*8-1 downto  70*8), w72 => Pw(61)( 72*8-1 downto  71*8), 
w73 => Pw(61)( 73*8-1 downto  72*8), w74 => Pw(61)( 74*8-1 downto  73*8), w75 => Pw(61)( 75*8-1 downto  74*8), w76 => Pw(61)( 76*8-1 downto  75*8), w77 => Pw(61)( 77*8-1 downto  76*8), w78 => Pw(61)( 78*8-1 downto  77*8), w79 => Pw(61)( 79*8-1 downto  78*8), w80 => Pw(61)( 80*8-1 downto  79*8), 
w81 => Pw(61)( 81*8-1 downto  80*8), w82 => Pw(61)( 82*8-1 downto  81*8), w83 => Pw(61)( 83*8-1 downto  82*8), w84 => Pw(61)( 84*8-1 downto  83*8), w85 => Pw(61)( 85*8-1 downto  84*8), w86 => Pw(61)( 86*8-1 downto  85*8), w87 => Pw(61)( 87*8-1 downto  86*8), w88 => Pw(61)( 88*8-1 downto  87*8), 
w89 => Pw(61)( 89*8-1 downto  88*8), w90 => Pw(61)( 90*8-1 downto  89*8), w91 => Pw(61)( 91*8-1 downto  90*8), w92 => Pw(61)( 92*8-1 downto  91*8), w93 => Pw(61)( 93*8-1 downto  92*8), w94 => Pw(61)( 94*8-1 downto  93*8), w95 => Pw(61)( 95*8-1 downto  94*8), w96 => Pw(61)( 96*8-1 downto  95*8), 
w97 => Pw(61)( 97*8-1 downto  96*8), w98 => Pw(61)( 98*8-1 downto  97*8), w99 => Pw(61)( 99*8-1 downto  98*8), w100=> Pw(61)(100*8-1 downto  99*8), w101=> Pw(61)(101*8-1 downto 100*8), w102=> Pw(61)(102*8-1 downto 101*8), w103=> Pw(61)(103*8-1 downto 102*8), w104=> Pw(61)(104*8-1 downto 103*8), 
w105=> Pw(61)(105*8-1 downto 104*8), w106=> Pw(61)(106*8-1 downto 105*8), w107=> Pw(61)(107*8-1 downto 106*8), w108=> Pw(61)(108*8-1 downto 107*8), w109=> Pw(61)(109*8-1 downto 108*8), w110=> Pw(61)(110*8-1 downto 109*8), w111=> Pw(61)(111*8-1 downto 110*8), w112=> Pw(61)(112*8-1 downto 111*8), 
w113=> Pw(61)(113*8-1 downto 112*8), w114=> Pw(61)(114*8-1 downto 113*8), w115=> Pw(61)(115*8-1 downto 114*8), w116=> Pw(61)(116*8-1 downto 115*8), w117=> Pw(61)(117*8-1 downto 116*8), w118=> Pw(61)(118*8-1 downto 117*8), w119=> Pw(61)(119*8-1 downto 118*8), w120=> Pw(61)(120*8-1 downto 119*8), 
w121=> Pw(61)(121*8-1 downto 120*8), w122=> Pw(61)(122*8-1 downto 121*8), w123=> Pw(61)(123*8-1 downto 122*8), w124=> Pw(61)(124*8-1 downto 123*8), w125=> Pw(61)(125*8-1 downto 124*8), w126=> Pw(61)(126*8-1 downto 125*8), w127=> Pw(61)(127*8-1 downto 126*8), w128=> Pw(61)(128*8-1 downto 127*8), 

           d_out   => pca_d61_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_62_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(62)(     7 downto    0), w02 => Pw(62)( 2*8-1 downto    8), w03 => Pw(62)( 3*8-1 downto  2*8), w04 => Pw(62)( 4*8-1 downto  3*8), w05 => Pw(62)( 5*8-1 downto  4*8), w06 => Pw(62)( 6*8-1 downto  5*8), w07 => Pw(62)( 7*8-1 downto  6*8), w08 => Pw(62)( 8*8-1 downto  7*8),  
w09 => Pw(62)( 9*8-1 downto  8*8), w10 => Pw(62)(10*8-1 downto  9*8), w11 => Pw(62)(11*8-1 downto 10*8), w12 => Pw(62)(12*8-1 downto 11*8), w13 => Pw(62)(13*8-1 downto 12*8), w14 => Pw(62)(14*8-1 downto 13*8), w15 => Pw(62)(15*8-1 downto 14*8), w16 => Pw(62)(16*8-1 downto 15*8),  
w17 => Pw(62)(17*8-1 downto 16*8), w18 => Pw(62)(18*8-1 downto 17*8), w19 => Pw(62)(19*8-1 downto 18*8), w20 => Pw(62)(20*8-1 downto 19*8), w21 => Pw(62)(21*8-1 downto 20*8), w22 => Pw(62)(22*8-1 downto 21*8), w23 => Pw(62)(23*8-1 downto 22*8), w24 => Pw(62)(24*8-1 downto 23*8),  
w25 => Pw(62)(25*8-1 downto 24*8), w26 => Pw(62)(26*8-1 downto 25*8), w27 => Pw(62)(27*8-1 downto 26*8), w28 => Pw(62)(28*8-1 downto 27*8), w29 => Pw(62)(29*8-1 downto 28*8), w30 => Pw(62)(30*8-1 downto 29*8), w31 => Pw(62)(31*8-1 downto 30*8), w32 => Pw(62)(32*8-1 downto 31*8),  
w33 => Pw(62)(33*8-1 downto 32*8), w34 => Pw(62)(34*8-1 downto 33*8), w35 => Pw(62)(35*8-1 downto 34*8), w36 => Pw(62)(36*8-1 downto 35*8), w37 => Pw(62)(37*8-1 downto 36*8), w38 => Pw(62)(38*8-1 downto 37*8), w39 => Pw(62)(39*8-1 downto 38*8), w40 => Pw(62)(40*8-1 downto 39*8),  
w41 => Pw(62)(41*8-1 downto 40*8), w42 => Pw(62)(42*8-1 downto 41*8), w43 => Pw(62)(43*8-1 downto 42*8), w44 => Pw(62)(44*8-1 downto 43*8), w45 => Pw(62)(45*8-1 downto 44*8), w46 => Pw(62)(46*8-1 downto 45*8), w47 => Pw(62)(47*8-1 downto 46*8), w48 => Pw(62)(48*8-1 downto 47*8),  
w49 => Pw(62)(49*8-1 downto 48*8), w50 => Pw(62)(50*8-1 downto 49*8), w51 => Pw(62)(51*8-1 downto 50*8), w52 => Pw(62)(52*8-1 downto 51*8), w53 => Pw(62)(53*8-1 downto 52*8), w54 => Pw(62)(54*8-1 downto 53*8), w55 => Pw(62)(55*8-1 downto 54*8), w56 => Pw(62)(56*8-1 downto 55*8),  
w57 => Pw(62)(57*8-1 downto 56*8), w58 => Pw(62)(58*8-1 downto 57*8), w59 => Pw(62)(59*8-1 downto 58*8), w60 => Pw(62)(60*8-1 downto 59*8), w61 => Pw(62)(61*8-1 downto 60*8), w62 => Pw(62)(62*8-1 downto 61*8), w63 => Pw(62)(63*8-1 downto 62*8), w64 => Pw(62)(64*8-1 downto 63*8), 
w65 => Pw(62)( 65*8-1 downto  64*8), w66 => Pw(62)( 66*8-1 downto  65*8), w67 => Pw(62)( 67*8-1 downto  66*8), w68 => Pw(62)( 68*8-1 downto  67*8), w69 => Pw(62)( 69*8-1 downto  68*8), w70 => Pw(62)( 70*8-1 downto  69*8), w71 => Pw(62)( 71*8-1 downto  70*8), w72 => Pw(62)( 72*8-1 downto  71*8), 
w73 => Pw(62)( 73*8-1 downto  72*8), w74 => Pw(62)( 74*8-1 downto  73*8), w75 => Pw(62)( 75*8-1 downto  74*8), w76 => Pw(62)( 76*8-1 downto  75*8), w77 => Pw(62)( 77*8-1 downto  76*8), w78 => Pw(62)( 78*8-1 downto  77*8), w79 => Pw(62)( 79*8-1 downto  78*8), w80 => Pw(62)( 80*8-1 downto  79*8), 
w81 => Pw(62)( 81*8-1 downto  80*8), w82 => Pw(62)( 82*8-1 downto  81*8), w83 => Pw(62)( 83*8-1 downto  82*8), w84 => Pw(62)( 84*8-1 downto  83*8), w85 => Pw(62)( 85*8-1 downto  84*8), w86 => Pw(62)( 86*8-1 downto  85*8), w87 => Pw(62)( 87*8-1 downto  86*8), w88 => Pw(62)( 88*8-1 downto  87*8), 
w89 => Pw(62)( 89*8-1 downto  88*8), w90 => Pw(62)( 90*8-1 downto  89*8), w91 => Pw(62)( 91*8-1 downto  90*8), w92 => Pw(62)( 92*8-1 downto  91*8), w93 => Pw(62)( 93*8-1 downto  92*8), w94 => Pw(62)( 94*8-1 downto  93*8), w95 => Pw(62)( 95*8-1 downto  94*8), w96 => Pw(62)( 96*8-1 downto  95*8), 
w97 => Pw(62)( 97*8-1 downto  96*8), w98 => Pw(62)( 98*8-1 downto  97*8), w99 => Pw(62)( 99*8-1 downto  98*8), w100=> Pw(62)(100*8-1 downto  99*8), w101=> Pw(62)(101*8-1 downto 100*8), w102=> Pw(62)(102*8-1 downto 101*8), w103=> Pw(62)(103*8-1 downto 102*8), w104=> Pw(62)(104*8-1 downto 103*8), 
w105=> Pw(62)(105*8-1 downto 104*8), w106=> Pw(62)(106*8-1 downto 105*8), w107=> Pw(62)(107*8-1 downto 106*8), w108=> Pw(62)(108*8-1 downto 107*8), w109=> Pw(62)(109*8-1 downto 108*8), w110=> Pw(62)(110*8-1 downto 109*8), w111=> Pw(62)(111*8-1 downto 110*8), w112=> Pw(62)(112*8-1 downto 111*8), 
w113=> Pw(62)(113*8-1 downto 112*8), w114=> Pw(62)(114*8-1 downto 113*8), w115=> Pw(62)(115*8-1 downto 114*8), w116=> Pw(62)(116*8-1 downto 115*8), w117=> Pw(62)(117*8-1 downto 116*8), w118=> Pw(62)(118*8-1 downto 117*8), w119=> Pw(62)(119*8-1 downto 118*8), w120=> Pw(62)(120*8-1 downto 119*8), 
w121=> Pw(62)(121*8-1 downto 120*8), w122=> Pw(62)(122*8-1 downto 121*8), w123=> Pw(62)(123*8-1 downto 122*8), w124=> Pw(62)(124*8-1 downto 123*8), w125=> Pw(62)(125*8-1 downto 124*8), w126=> Pw(62)(126*8-1 downto 125*8), w127=> Pw(62)(127*8-1 downto 126*8), w128=> Pw(62)(128*8-1 downto 127*8), 

           d_out   => pca_d62_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_63_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,  

w01 => Pw(63)(     7 downto    0), w02 => Pw(63)( 2*8-1 downto    8), w03 => Pw(63)( 3*8-1 downto  2*8), w04 => Pw(63)( 4*8-1 downto  3*8), w05 => Pw(63)( 5*8-1 downto  4*8), w06 => Pw(63)( 6*8-1 downto  5*8), w07 => Pw(63)( 7*8-1 downto  6*8), w08 => Pw(63)( 8*8-1 downto  7*8),  
w09 => Pw(63)( 9*8-1 downto  8*8), w10 => Pw(63)(10*8-1 downto  9*8), w11 => Pw(63)(11*8-1 downto 10*8), w12 => Pw(63)(12*8-1 downto 11*8), w13 => Pw(63)(13*8-1 downto 12*8), w14 => Pw(63)(14*8-1 downto 13*8), w15 => Pw(63)(15*8-1 downto 14*8), w16 => Pw(63)(16*8-1 downto 15*8),  
w17 => Pw(63)(17*8-1 downto 16*8), w18 => Pw(63)(18*8-1 downto 17*8), w19 => Pw(63)(19*8-1 downto 18*8), w20 => Pw(63)(20*8-1 downto 19*8), w21 => Pw(63)(21*8-1 downto 20*8), w22 => Pw(63)(22*8-1 downto 21*8), w23 => Pw(63)(23*8-1 downto 22*8), w24 => Pw(63)(24*8-1 downto 23*8),  
w25 => Pw(63)(25*8-1 downto 24*8), w26 => Pw(63)(26*8-1 downto 25*8), w27 => Pw(63)(27*8-1 downto 26*8), w28 => Pw(63)(28*8-1 downto 27*8), w29 => Pw(63)(29*8-1 downto 28*8), w30 => Pw(63)(30*8-1 downto 29*8), w31 => Pw(63)(31*8-1 downto 30*8), w32 => Pw(63)(32*8-1 downto 31*8),  
w33 => Pw(63)(33*8-1 downto 32*8), w34 => Pw(63)(34*8-1 downto 33*8), w35 => Pw(63)(35*8-1 downto 34*8), w36 => Pw(63)(36*8-1 downto 35*8), w37 => Pw(63)(37*8-1 downto 36*8), w38 => Pw(63)(38*8-1 downto 37*8), w39 => Pw(63)(39*8-1 downto 38*8), w40 => Pw(63)(40*8-1 downto 39*8),  
w41 => Pw(63)(41*8-1 downto 40*8), w42 => Pw(63)(42*8-1 downto 41*8), w43 => Pw(63)(43*8-1 downto 42*8), w44 => Pw(63)(44*8-1 downto 43*8), w45 => Pw(63)(45*8-1 downto 44*8), w46 => Pw(63)(46*8-1 downto 45*8), w47 => Pw(63)(47*8-1 downto 46*8), w48 => Pw(63)(48*8-1 downto 47*8),  
w49 => Pw(63)(49*8-1 downto 48*8), w50 => Pw(63)(50*8-1 downto 49*8), w51 => Pw(63)(51*8-1 downto 50*8), w52 => Pw(63)(52*8-1 downto 51*8), w53 => Pw(63)(53*8-1 downto 52*8), w54 => Pw(63)(54*8-1 downto 53*8), w55 => Pw(63)(55*8-1 downto 54*8), w56 => Pw(63)(56*8-1 downto 55*8),  
w57 => Pw(63)(57*8-1 downto 56*8), w58 => Pw(63)(58*8-1 downto 57*8), w59 => Pw(63)(59*8-1 downto 58*8), w60 => Pw(63)(60*8-1 downto 59*8), w61 => Pw(63)(61*8-1 downto 60*8), w62 => Pw(63)(62*8-1 downto 61*8), w63 => Pw(63)(63*8-1 downto 62*8), w64 => Pw(63)(64*8-1 downto 63*8), 
w65 => Pw(63)( 65*8-1 downto  64*8), w66 => Pw(63)( 66*8-1 downto  65*8), w67 => Pw(63)( 67*8-1 downto  66*8), w68 => Pw(63)( 68*8-1 downto  67*8), w69 => Pw(63)( 69*8-1 downto  68*8), w70 => Pw(63)( 70*8-1 downto  69*8), w71 => Pw(63)( 71*8-1 downto  70*8), w72 => Pw(63)( 72*8-1 downto  71*8), 
w73 => Pw(63)( 73*8-1 downto  72*8), w74 => Pw(63)( 74*8-1 downto  73*8), w75 => Pw(63)( 75*8-1 downto  74*8), w76 => Pw(63)( 76*8-1 downto  75*8), w77 => Pw(63)( 77*8-1 downto  76*8), w78 => Pw(63)( 78*8-1 downto  77*8), w79 => Pw(63)( 79*8-1 downto  78*8), w80 => Pw(63)( 80*8-1 downto  79*8), 
w81 => Pw(63)( 81*8-1 downto  80*8), w82 => Pw(63)( 82*8-1 downto  81*8), w83 => Pw(63)( 83*8-1 downto  82*8), w84 => Pw(63)( 84*8-1 downto  83*8), w85 => Pw(63)( 85*8-1 downto  84*8), w86 => Pw(63)( 86*8-1 downto  85*8), w87 => Pw(63)( 87*8-1 downto  86*8), w88 => Pw(63)( 88*8-1 downto  87*8), 
w89 => Pw(63)( 89*8-1 downto  88*8), w90 => Pw(63)( 90*8-1 downto  89*8), w91 => Pw(63)( 91*8-1 downto  90*8), w92 => Pw(63)( 92*8-1 downto  91*8), w93 => Pw(63)( 93*8-1 downto  92*8), w94 => Pw(63)( 94*8-1 downto  93*8), w95 => Pw(63)( 95*8-1 downto  94*8), w96 => Pw(63)( 96*8-1 downto  95*8), 
w97 => Pw(63)( 97*8-1 downto  96*8), w98 => Pw(63)( 98*8-1 downto  97*8), w99 => Pw(63)( 99*8-1 downto  98*8), w100=> Pw(63)(100*8-1 downto  99*8), w101=> Pw(63)(101*8-1 downto 100*8), w102=> Pw(63)(102*8-1 downto 101*8), w103=> Pw(63)(103*8-1 downto 102*8), w104=> Pw(63)(104*8-1 downto 103*8), 
w105=> Pw(63)(105*8-1 downto 104*8), w106=> Pw(63)(106*8-1 downto 105*8), w107=> Pw(63)(107*8-1 downto 106*8), w108=> Pw(63)(108*8-1 downto 107*8), w109=> Pw(63)(109*8-1 downto 108*8), w110=> Pw(63)(110*8-1 downto 109*8), w111=> Pw(63)(111*8-1 downto 110*8), w112=> Pw(63)(112*8-1 downto 111*8), 
w113=> Pw(63)(113*8-1 downto 112*8), w114=> Pw(63)(114*8-1 downto 113*8), w115=> Pw(63)(115*8-1 downto 114*8), w116=> Pw(63)(116*8-1 downto 115*8), w117=> Pw(63)(117*8-1 downto 116*8), w118=> Pw(63)(118*8-1 downto 117*8), w119=> Pw(63)(119*8-1 downto 118*8), w120=> Pw(63)(120*8-1 downto 119*8), 
w121=> Pw(63)(121*8-1 downto 120*8), w122=> Pw(63)(122*8-1 downto 121*8), w123=> Pw(63)(123*8-1 downto 122*8), w124=> Pw(63)(124*8-1 downto 123*8), w125=> Pw(63)(125*8-1 downto 124*8), w126=> Pw(63)(126*8-1 downto 125*8), w127=> Pw(63)(127*8-1 downto 126*8), w128=> Pw(63)(128*8-1 downto 127*8), 

           d_out   => pca_d63_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_64_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(64)(     7 downto    0),   w02 => Pw(64)( 2*8-1 downto    8),   w03 => Pw(64)( 3*8-1 downto  2*8),   w04 => Pw(64)( 4*8-1 downto  3*8),   w05 => Pw(64)( 5*8-1 downto  4*8),   w06 => Pw(64)( 6*8-1 downto  5*8),   w07 => Pw(64)( 7*8-1 downto  6*8),   w08 => Pw(64)( 8*8-1 downto  7*8),  
w09 => Pw(64)( 9*8-1 downto  8*8),   w10 => Pw(64)(10*8-1 downto  9*8),   w11 => Pw(64)(11*8-1 downto 10*8),   w12 => Pw(64)(12*8-1 downto 11*8),   w13 => Pw(64)(13*8-1 downto 12*8),   w14 => Pw(64)(14*8-1 downto 13*8),   w15 => Pw(64)(15*8-1 downto 14*8),   w16 => Pw(64)(16*8-1 downto 15*8),  
w17 => Pw(64)(17*8-1 downto 16*8),   w18 => Pw(64)(18*8-1 downto 17*8),   w19 => Pw(64)(19*8-1 downto 18*8),   w20 => Pw(64)(20*8-1 downto 19*8),   w21 => Pw(64)(21*8-1 downto 20*8),   w22 => Pw(64)(22*8-1 downto 21*8),   w23 => Pw(64)(23*8-1 downto 22*8),   w24 => Pw(64)(24*8-1 downto 23*8),  
w25 => Pw(64)(25*8-1 downto 24*8),   w26 => Pw(64)(26*8-1 downto 25*8),   w27 => Pw(64)(27*8-1 downto 26*8),   w28 => Pw(64)(28*8-1 downto 27*8),   w29 => Pw(64)(29*8-1 downto 28*8),   w30 => Pw(64)(30*8-1 downto 29*8),   w31 => Pw(64)(31*8-1 downto 30*8),   w32 => Pw(64)(32*8-1 downto 31*8),  
w33 => Pw(64)(33*8-1 downto 32*8),   w34 => Pw(64)(34*8-1 downto 33*8),   w35 => Pw(64)(35*8-1 downto 34*8),   w36 => Pw(64)(36*8-1 downto 35*8),   w37 => Pw(64)(37*8-1 downto 36*8),   w38 => Pw(64)(38*8-1 downto 37*8),   w39 => Pw(64)(39*8-1 downto 38*8),   w40 => Pw(64)(40*8-1 downto 39*8),  
w41 => Pw(64)(41*8-1 downto 40*8),   w42 => Pw(64)(42*8-1 downto 41*8),   w43 => Pw(64)(43*8-1 downto 42*8),   w44 => Pw(64)(44*8-1 downto 43*8),   w45 => Pw(64)(45*8-1 downto 44*8),   w46 => Pw(64)(46*8-1 downto 45*8),   w47 => Pw(64)(47*8-1 downto 46*8),   w48 => Pw(64)(48*8-1 downto 47*8),  
w49 => Pw(64)(49*8-1 downto 48*8),   w50 => Pw(64)(50*8-1 downto 49*8),   w51 => Pw(64)(51*8-1 downto 50*8),   w52 => Pw(64)(52*8-1 downto 51*8),   w53 => Pw(64)(53*8-1 downto 52*8),   w54 => Pw(64)(54*8-1 downto 53*8),   w55 => Pw(64)(55*8-1 downto 54*8),   w56 => Pw(64)(56*8-1 downto 55*8),  
w57 => Pw(64)(57*8-1 downto 56*8),   w58 => Pw(64)(58*8-1 downto 57*8),   w59 => Pw(64)(59*8-1 downto 58*8),   w60 => Pw(64)(60*8-1 downto 59*8),   w61 => Pw(64)(61*8-1 downto 60*8),   w62 => Pw(64)(62*8-1 downto 61*8),   w63 => Pw(64)(63*8-1 downto 62*8),   w64 => Pw(64)(64*8-1 downto 63*8), 
w65 => Pw(64)( 65*8-1 downto  64*8), w66 => Pw(64)( 66*8-1 downto  65*8), w67 => Pw(64)( 67*8-1 downto  66*8), w68 => Pw(64)( 68*8-1 downto  67*8), w69 => Pw(64)( 69*8-1 downto  68*8), w70 => Pw(64)( 70*8-1 downto  69*8), w71 => Pw(64)( 71*8-1 downto  70*8), w72 => Pw(64)( 72*8-1 downto  71*8), 
w73 => Pw(64)( 73*8-1 downto  72*8), w74 => Pw(64)( 74*8-1 downto  73*8), w75 => Pw(64)( 75*8-1 downto  74*8), w76 => Pw(64)( 76*8-1 downto  75*8), w77 => Pw(64)( 77*8-1 downto  76*8), w78 => Pw(64)( 78*8-1 downto  77*8), w79 => Pw(64)( 79*8-1 downto  78*8), w80 => Pw(64)( 80*8-1 downto  79*8), 
w81 => Pw(64)( 81*8-1 downto  80*8), w82 => Pw(64)( 82*8-1 downto  81*8), w83 => Pw(64)( 83*8-1 downto  82*8), w84 => Pw(64)( 84*8-1 downto  83*8), w85 => Pw(64)( 85*8-1 downto  84*8), w86 => Pw(64)( 86*8-1 downto  85*8), w87 => Pw(64)( 87*8-1 downto  86*8), w88 => Pw(64)( 88*8-1 downto  87*8), 
w89 => Pw(64)( 89*8-1 downto  88*8), w90 => Pw(64)( 90*8-1 downto  89*8), w91 => Pw(64)( 91*8-1 downto  90*8), w92 => Pw(64)( 92*8-1 downto  91*8), w93 => Pw(64)( 93*8-1 downto  92*8), w94 => Pw(64)( 94*8-1 downto  93*8), w95 => Pw(64)( 95*8-1 downto  94*8), w96 => Pw(64)( 96*8-1 downto  95*8), 
w97 => Pw(64)( 97*8-1 downto  96*8), w98 => Pw(64)( 98*8-1 downto  97*8), w99 => Pw(64)( 99*8-1 downto  98*8), w100=> Pw(64)(100*8-1 downto  99*8), w101=> Pw(64)(101*8-1 downto 100*8), w102=> Pw(64)(102*8-1 downto 101*8), w103=> Pw(64)(103*8-1 downto 102*8), w104=> Pw(64)(104*8-1 downto 103*8), 
w105=> Pw(64)(105*8-1 downto 104*8), w106=> Pw(64)(106*8-1 downto 105*8), w107=> Pw(64)(107*8-1 downto 106*8), w108=> Pw(64)(108*8-1 downto 107*8), w109=> Pw(64)(109*8-1 downto 108*8), w110=> Pw(64)(110*8-1 downto 109*8), w111=> Pw(64)(111*8-1 downto 110*8), w112=> Pw(64)(112*8-1 downto 111*8), 
w113=> Pw(64)(113*8-1 downto 112*8), w114=> Pw(64)(114*8-1 downto 113*8), w115=> Pw(64)(115*8-1 downto 114*8), w116=> Pw(64)(116*8-1 downto 115*8), w117=> Pw(64)(117*8-1 downto 116*8), w118=> Pw(64)(118*8-1 downto 117*8), w119=> Pw(64)(119*8-1 downto 118*8), w120=> Pw(64)(120*8-1 downto 119*8), 
w121=> Pw(64)(121*8-1 downto 120*8), w122=> Pw(64)(122*8-1 downto 121*8), w123=> Pw(64)(123*8-1 downto 122*8), w124=> Pw(64)(124*8-1 downto 123*8), w125=> Pw(64)(125*8-1 downto 124*8), w126=> Pw(64)(126*8-1 downto 125*8), w127=> Pw(64)(127*8-1 downto 126*8), w128=> Pw(64)(128*8-1 downto 127*8), 
           d_out   => pca_d64_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_65_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(65)(     7 downto    0),   w02 => Pw(65)( 2*8-1 downto    8),   w03 => Pw(65)( 3*8-1 downto  2*8),   w04 => Pw(65)( 4*8-1 downto  3*8),   w05 => Pw(65)( 5*8-1 downto  4*8),   w06 => Pw(65)( 6*8-1 downto  5*8),   w07 => Pw(65)( 7*8-1 downto  6*8),   w08 => Pw(65)( 8*8-1 downto  7*8),  
w09 => Pw(65)( 9*8-1 downto  8*8),   w10 => Pw(65)(10*8-1 downto  9*8),   w11 => Pw(65)(11*8-1 downto 10*8),   w12 => Pw(65)(12*8-1 downto 11*8),   w13 => Pw(65)(13*8-1 downto 12*8),   w14 => Pw(65)(14*8-1 downto 13*8),   w15 => Pw(65)(15*8-1 downto 14*8),   w16 => Pw(65)(16*8-1 downto 15*8),  
w17 => Pw(65)(17*8-1 downto 16*8),   w18 => Pw(65)(18*8-1 downto 17*8),   w19 => Pw(65)(19*8-1 downto 18*8),   w20 => Pw(65)(20*8-1 downto 19*8),   w21 => Pw(65)(21*8-1 downto 20*8),   w22 => Pw(65)(22*8-1 downto 21*8),   w23 => Pw(65)(23*8-1 downto 22*8),   w24 => Pw(65)(24*8-1 downto 23*8),  
w25 => Pw(65)(25*8-1 downto 24*8),   w26 => Pw(65)(26*8-1 downto 25*8),   w27 => Pw(65)(27*8-1 downto 26*8),   w28 => Pw(65)(28*8-1 downto 27*8),   w29 => Pw(65)(29*8-1 downto 28*8),   w30 => Pw(65)(30*8-1 downto 29*8),   w31 => Pw(65)(31*8-1 downto 30*8),   w32 => Pw(65)(32*8-1 downto 31*8),  
w33 => Pw(65)(33*8-1 downto 32*8),   w34 => Pw(65)(34*8-1 downto 33*8),   w35 => Pw(65)(35*8-1 downto 34*8),   w36 => Pw(65)(36*8-1 downto 35*8),   w37 => Pw(65)(37*8-1 downto 36*8),   w38 => Pw(65)(38*8-1 downto 37*8),   w39 => Pw(65)(39*8-1 downto 38*8),   w40 => Pw(65)(40*8-1 downto 39*8),  
w41 => Pw(65)(41*8-1 downto 40*8),   w42 => Pw(65)(42*8-1 downto 41*8),   w43 => Pw(65)(43*8-1 downto 42*8),   w44 => Pw(65)(44*8-1 downto 43*8),   w45 => Pw(65)(45*8-1 downto 44*8),   w46 => Pw(65)(46*8-1 downto 45*8),   w47 => Pw(65)(47*8-1 downto 46*8),   w48 => Pw(65)(48*8-1 downto 47*8),  
w49 => Pw(65)(49*8-1 downto 48*8),   w50 => Pw(65)(50*8-1 downto 49*8),   w51 => Pw(65)(51*8-1 downto 50*8),   w52 => Pw(65)(52*8-1 downto 51*8),   w53 => Pw(65)(53*8-1 downto 52*8),   w54 => Pw(65)(54*8-1 downto 53*8),   w55 => Pw(65)(55*8-1 downto 54*8),   w56 => Pw(65)(56*8-1 downto 55*8),  
w57 => Pw(65)(57*8-1 downto 56*8),   w58 => Pw(65)(58*8-1 downto 57*8),   w59 => Pw(65)(59*8-1 downto 58*8),   w60 => Pw(65)(60*8-1 downto 59*8),   w61 => Pw(65)(61*8-1 downto 60*8),   w62 => Pw(65)(62*8-1 downto 61*8),   w63 => Pw(65)(63*8-1 downto 62*8),   w64 => Pw(65)(64*8-1 downto 63*8), 
w65 => Pw(65)( 65*8-1 downto  64*8), w66 => Pw(65)( 66*8-1 downto  65*8), w67 => Pw(65)( 67*8-1 downto  66*8), w68 => Pw(65)( 68*8-1 downto  67*8), w69 => Pw(65)( 69*8-1 downto  68*8), w70 => Pw(65)( 70*8-1 downto  69*8), w71 => Pw(65)( 71*8-1 downto  70*8), w72 => Pw(65)( 72*8-1 downto  71*8), 
w73 => Pw(65)( 73*8-1 downto  72*8), w74 => Pw(65)( 74*8-1 downto  73*8), w75 => Pw(65)( 75*8-1 downto  74*8), w76 => Pw(65)( 76*8-1 downto  75*8), w77 => Pw(65)( 77*8-1 downto  76*8), w78 => Pw(65)( 78*8-1 downto  77*8), w79 => Pw(65)( 79*8-1 downto  78*8), w80 => Pw(65)( 80*8-1 downto  79*8), 
w81 => Pw(65)( 81*8-1 downto  80*8), w82 => Pw(65)( 82*8-1 downto  81*8), w83 => Pw(65)( 83*8-1 downto  82*8), w84 => Pw(65)( 84*8-1 downto  83*8), w85 => Pw(65)( 85*8-1 downto  84*8), w86 => Pw(65)( 86*8-1 downto  85*8), w87 => Pw(65)( 87*8-1 downto  86*8), w88 => Pw(65)( 88*8-1 downto  87*8), 
w89 => Pw(65)( 89*8-1 downto  88*8), w90 => Pw(65)( 90*8-1 downto  89*8), w91 => Pw(65)( 91*8-1 downto  90*8), w92 => Pw(65)( 92*8-1 downto  91*8), w93 => Pw(65)( 93*8-1 downto  92*8), w94 => Pw(65)( 94*8-1 downto  93*8), w95 => Pw(65)( 95*8-1 downto  94*8), w96 => Pw(65)( 96*8-1 downto  95*8), 
w97 => Pw(65)( 97*8-1 downto  96*8), w98 => Pw(65)( 98*8-1 downto  97*8), w99 => Pw(65)( 99*8-1 downto  98*8), w100=> Pw(65)(100*8-1 downto  99*8), w101=> Pw(65)(101*8-1 downto 100*8), w102=> Pw(65)(102*8-1 downto 101*8), w103=> Pw(65)(103*8-1 downto 102*8), w104=> Pw(65)(104*8-1 downto 103*8), 
w105=> Pw(65)(105*8-1 downto 104*8), w106=> Pw(65)(106*8-1 downto 105*8), w107=> Pw(65)(107*8-1 downto 106*8), w108=> Pw(65)(108*8-1 downto 107*8), w109=> Pw(65)(109*8-1 downto 108*8), w110=> Pw(65)(110*8-1 downto 109*8), w111=> Pw(65)(111*8-1 downto 110*8), w112=> Pw(65)(112*8-1 downto 111*8), 
w113=> Pw(65)(113*8-1 downto 112*8), w114=> Pw(65)(114*8-1 downto 113*8), w115=> Pw(65)(115*8-1 downto 114*8), w116=> Pw(65)(116*8-1 downto 115*8), w117=> Pw(65)(117*8-1 downto 116*8), w118=> Pw(65)(118*8-1 downto 117*8), w119=> Pw(65)(119*8-1 downto 118*8), w120=> Pw(65)(120*8-1 downto 119*8), 
w121=> Pw(65)(121*8-1 downto 120*8), w122=> Pw(65)(122*8-1 downto 121*8), w123=> Pw(65)(123*8-1 downto 122*8), w124=> Pw(65)(124*8-1 downto 123*8), w125=> Pw(65)(125*8-1 downto 124*8), w126=> Pw(65)(126*8-1 downto 125*8), w127=> Pw(65)(127*8-1 downto 126*8), w128=> Pw(65)(128*8-1 downto 127*8), 
           d_out   => pca_d65_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_66_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(66)(     7 downto    0),   w02 => Pw(66)( 2*8-1 downto    8),   w03 => Pw(66)( 3*8-1 downto  2*8),   w04 => Pw(66)( 4*8-1 downto  3*8),   w05 => Pw(66)( 5*8-1 downto  4*8),   w06 => Pw(66)( 6*8-1 downto  5*8),   w07 => Pw(66)( 7*8-1 downto  6*8),   w08 => Pw(66)( 8*8-1 downto  7*8),  
w09 => Pw(66)( 9*8-1 downto  8*8),   w10 => Pw(66)(10*8-1 downto  9*8),   w11 => Pw(66)(11*8-1 downto 10*8),   w12 => Pw(66)(12*8-1 downto 11*8),   w13 => Pw(66)(13*8-1 downto 12*8),   w14 => Pw(66)(14*8-1 downto 13*8),   w15 => Pw(66)(15*8-1 downto 14*8),   w16 => Pw(66)(16*8-1 downto 15*8),  
w17 => Pw(66)(17*8-1 downto 16*8),   w18 => Pw(66)(18*8-1 downto 17*8),   w19 => Pw(66)(19*8-1 downto 18*8),   w20 => Pw(66)(20*8-1 downto 19*8),   w21 => Pw(66)(21*8-1 downto 20*8),   w22 => Pw(66)(22*8-1 downto 21*8),   w23 => Pw(66)(23*8-1 downto 22*8),   w24 => Pw(66)(24*8-1 downto 23*8),  
w25 => Pw(66)(25*8-1 downto 24*8),   w26 => Pw(66)(26*8-1 downto 25*8),   w27 => Pw(66)(27*8-1 downto 26*8),   w28 => Pw(66)(28*8-1 downto 27*8),   w29 => Pw(66)(29*8-1 downto 28*8),   w30 => Pw(66)(30*8-1 downto 29*8),   w31 => Pw(66)(31*8-1 downto 30*8),   w32 => Pw(66)(32*8-1 downto 31*8),  
w33 => Pw(66)(33*8-1 downto 32*8),   w34 => Pw(66)(34*8-1 downto 33*8),   w35 => Pw(66)(35*8-1 downto 34*8),   w36 => Pw(66)(36*8-1 downto 35*8),   w37 => Pw(66)(37*8-1 downto 36*8),   w38 => Pw(66)(38*8-1 downto 37*8),   w39 => Pw(66)(39*8-1 downto 38*8),   w40 => Pw(66)(40*8-1 downto 39*8),  
w41 => Pw(66)(41*8-1 downto 40*8),   w42 => Pw(66)(42*8-1 downto 41*8),   w43 => Pw(66)(43*8-1 downto 42*8),   w44 => Pw(66)(44*8-1 downto 43*8),   w45 => Pw(66)(45*8-1 downto 44*8),   w46 => Pw(66)(46*8-1 downto 45*8),   w47 => Pw(66)(47*8-1 downto 46*8),   w48 => Pw(66)(48*8-1 downto 47*8),  
w49 => Pw(66)(49*8-1 downto 48*8),   w50 => Pw(66)(50*8-1 downto 49*8),   w51 => Pw(66)(51*8-1 downto 50*8),   w52 => Pw(66)(52*8-1 downto 51*8),   w53 => Pw(66)(53*8-1 downto 52*8),   w54 => Pw(66)(54*8-1 downto 53*8),   w55 => Pw(66)(55*8-1 downto 54*8),   w56 => Pw(66)(56*8-1 downto 55*8),  
w57 => Pw(66)(57*8-1 downto 56*8),   w58 => Pw(66)(58*8-1 downto 57*8),   w59 => Pw(66)(59*8-1 downto 58*8),   w60 => Pw(66)(60*8-1 downto 59*8),   w61 => Pw(66)(61*8-1 downto 60*8),   w62 => Pw(66)(62*8-1 downto 61*8),   w63 => Pw(66)(63*8-1 downto 62*8),   w64 => Pw(66)(64*8-1 downto 63*8), 
w65 => Pw(66)( 65*8-1 downto  64*8), w66 => Pw(66)( 66*8-1 downto  65*8), w67 => Pw(66)( 67*8-1 downto  66*8), w68 => Pw(66)( 68*8-1 downto  67*8), w69 => Pw(66)( 69*8-1 downto  68*8), w70 => Pw(66)( 70*8-1 downto  69*8), w71 => Pw(66)( 71*8-1 downto  70*8), w72 => Pw(66)( 72*8-1 downto  71*8), 
w73 => Pw(66)( 73*8-1 downto  72*8), w74 => Pw(66)( 74*8-1 downto  73*8), w75 => Pw(66)( 75*8-1 downto  74*8), w76 => Pw(66)( 76*8-1 downto  75*8), w77 => Pw(66)( 77*8-1 downto  76*8), w78 => Pw(66)( 78*8-1 downto  77*8), w79 => Pw(66)( 79*8-1 downto  78*8), w80 => Pw(66)( 80*8-1 downto  79*8), 
w81 => Pw(66)( 81*8-1 downto  80*8), w82 => Pw(66)( 82*8-1 downto  81*8), w83 => Pw(66)( 83*8-1 downto  82*8), w84 => Pw(66)( 84*8-1 downto  83*8), w85 => Pw(66)( 85*8-1 downto  84*8), w86 => Pw(66)( 86*8-1 downto  85*8), w87 => Pw(66)( 87*8-1 downto  86*8), w88 => Pw(66)( 88*8-1 downto  87*8), 
w89 => Pw(66)( 89*8-1 downto  88*8), w90 => Pw(66)( 90*8-1 downto  89*8), w91 => Pw(66)( 91*8-1 downto  90*8), w92 => Pw(66)( 92*8-1 downto  91*8), w93 => Pw(66)( 93*8-1 downto  92*8), w94 => Pw(66)( 94*8-1 downto  93*8), w95 => Pw(66)( 95*8-1 downto  94*8), w96 => Pw(66)( 96*8-1 downto  95*8), 
w97 => Pw(66)( 97*8-1 downto  96*8), w98 => Pw(66)( 98*8-1 downto  97*8), w99 => Pw(66)( 99*8-1 downto  98*8), w100=> Pw(66)(100*8-1 downto  99*8), w101=> Pw(66)(101*8-1 downto 100*8), w102=> Pw(66)(102*8-1 downto 101*8), w103=> Pw(66)(103*8-1 downto 102*8), w104=> Pw(66)(104*8-1 downto 103*8), 
w105=> Pw(66)(105*8-1 downto 104*8), w106=> Pw(66)(106*8-1 downto 105*8), w107=> Pw(66)(107*8-1 downto 106*8), w108=> Pw(66)(108*8-1 downto 107*8), w109=> Pw(66)(109*8-1 downto 108*8), w110=> Pw(66)(110*8-1 downto 109*8), w111=> Pw(66)(111*8-1 downto 110*8), w112=> Pw(66)(112*8-1 downto 111*8), 
w113=> Pw(66)(113*8-1 downto 112*8), w114=> Pw(66)(114*8-1 downto 113*8), w115=> Pw(66)(115*8-1 downto 114*8), w116=> Pw(66)(116*8-1 downto 115*8), w117=> Pw(66)(117*8-1 downto 116*8), w118=> Pw(66)(118*8-1 downto 117*8), w119=> Pw(66)(119*8-1 downto 118*8), w120=> Pw(66)(120*8-1 downto 119*8), 
w121=> Pw(66)(121*8-1 downto 120*8), w122=> Pw(66)(122*8-1 downto 121*8), w123=> Pw(66)(123*8-1 downto 122*8), w124=> Pw(66)(124*8-1 downto 123*8), w125=> Pw(66)(125*8-1 downto 124*8), w126=> Pw(66)(126*8-1 downto 125*8), w127=> Pw(66)(127*8-1 downto 126*8), w128=> Pw(66)(128*8-1 downto 127*8), 
           d_out   => pca_d66_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_67_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(67)(     7 downto    0),   w02 => Pw(67)( 2*8-1 downto    8),   w03 => Pw(67)( 3*8-1 downto  2*8),   w04 => Pw(67)( 4*8-1 downto  3*8),   w05 => Pw(67)( 5*8-1 downto  4*8),   w06 => Pw(67)( 6*8-1 downto  5*8),   w07 => Pw(67)( 7*8-1 downto  6*8),   w08 => Pw(67)( 8*8-1 downto  7*8),  
w09 => Pw(67)( 9*8-1 downto  8*8),   w10 => Pw(67)(10*8-1 downto  9*8),   w11 => Pw(67)(11*8-1 downto 10*8),   w12 => Pw(67)(12*8-1 downto 11*8),   w13 => Pw(67)(13*8-1 downto 12*8),   w14 => Pw(67)(14*8-1 downto 13*8),   w15 => Pw(67)(15*8-1 downto 14*8),   w16 => Pw(67)(16*8-1 downto 15*8),  
w17 => Pw(67)(17*8-1 downto 16*8),   w18 => Pw(67)(18*8-1 downto 17*8),   w19 => Pw(67)(19*8-1 downto 18*8),   w20 => Pw(67)(20*8-1 downto 19*8),   w21 => Pw(67)(21*8-1 downto 20*8),   w22 => Pw(67)(22*8-1 downto 21*8),   w23 => Pw(67)(23*8-1 downto 22*8),   w24 => Pw(67)(24*8-1 downto 23*8),  
w25 => Pw(67)(25*8-1 downto 24*8),   w26 => Pw(67)(26*8-1 downto 25*8),   w27 => Pw(67)(27*8-1 downto 26*8),   w28 => Pw(67)(28*8-1 downto 27*8),   w29 => Pw(67)(29*8-1 downto 28*8),   w30 => Pw(67)(30*8-1 downto 29*8),   w31 => Pw(67)(31*8-1 downto 30*8),   w32 => Pw(67)(32*8-1 downto 31*8),  
w33 => Pw(67)(33*8-1 downto 32*8),   w34 => Pw(67)(34*8-1 downto 33*8),   w35 => Pw(67)(35*8-1 downto 34*8),   w36 => Pw(67)(36*8-1 downto 35*8),   w37 => Pw(67)(37*8-1 downto 36*8),   w38 => Pw(67)(38*8-1 downto 37*8),   w39 => Pw(67)(39*8-1 downto 38*8),   w40 => Pw(67)(40*8-1 downto 39*8),  
w41 => Pw(67)(41*8-1 downto 40*8),   w42 => Pw(67)(42*8-1 downto 41*8),   w43 => Pw(67)(43*8-1 downto 42*8),   w44 => Pw(67)(44*8-1 downto 43*8),   w45 => Pw(67)(45*8-1 downto 44*8),   w46 => Pw(67)(46*8-1 downto 45*8),   w47 => Pw(67)(47*8-1 downto 46*8),   w48 => Pw(67)(48*8-1 downto 47*8),  
w49 => Pw(67)(49*8-1 downto 48*8),   w50 => Pw(67)(50*8-1 downto 49*8),   w51 => Pw(67)(51*8-1 downto 50*8),   w52 => Pw(67)(52*8-1 downto 51*8),   w53 => Pw(67)(53*8-1 downto 52*8),   w54 => Pw(67)(54*8-1 downto 53*8),   w55 => Pw(67)(55*8-1 downto 54*8),   w56 => Pw(67)(56*8-1 downto 55*8),  
w57 => Pw(67)(57*8-1 downto 56*8),   w58 => Pw(67)(58*8-1 downto 57*8),   w59 => Pw(67)(59*8-1 downto 58*8),   w60 => Pw(67)(60*8-1 downto 59*8),   w61 => Pw(67)(61*8-1 downto 60*8),   w62 => Pw(67)(62*8-1 downto 61*8),   w63 => Pw(67)(63*8-1 downto 62*8),   w64 => Pw(67)(64*8-1 downto 63*8), 
w65 => Pw(67)( 65*8-1 downto  64*8), w66 => Pw(67)( 66*8-1 downto  65*8), w67 => Pw(67)( 67*8-1 downto  66*8), w68 => Pw(67)( 68*8-1 downto  67*8), w69 => Pw(67)( 69*8-1 downto  68*8), w70 => Pw(67)( 70*8-1 downto  69*8), w71 => Pw(67)( 71*8-1 downto  70*8), w72 => Pw(67)( 72*8-1 downto  71*8), 
w73 => Pw(67)( 73*8-1 downto  72*8), w74 => Pw(67)( 74*8-1 downto  73*8), w75 => Pw(67)( 75*8-1 downto  74*8), w76 => Pw(67)( 76*8-1 downto  75*8), w77 => Pw(67)( 77*8-1 downto  76*8), w78 => Pw(67)( 78*8-1 downto  77*8), w79 => Pw(67)( 79*8-1 downto  78*8), w80 => Pw(67)( 80*8-1 downto  79*8), 
w81 => Pw(67)( 81*8-1 downto  80*8), w82 => Pw(67)( 82*8-1 downto  81*8), w83 => Pw(67)( 83*8-1 downto  82*8), w84 => Pw(67)( 84*8-1 downto  83*8), w85 => Pw(67)( 85*8-1 downto  84*8), w86 => Pw(67)( 86*8-1 downto  85*8), w87 => Pw(67)( 87*8-1 downto  86*8), w88 => Pw(67)( 88*8-1 downto  87*8), 
w89 => Pw(67)( 89*8-1 downto  88*8), w90 => Pw(67)( 90*8-1 downto  89*8), w91 => Pw(67)( 91*8-1 downto  90*8), w92 => Pw(67)( 92*8-1 downto  91*8), w93 => Pw(67)( 93*8-1 downto  92*8), w94 => Pw(67)( 94*8-1 downto  93*8), w95 => Pw(67)( 95*8-1 downto  94*8), w96 => Pw(67)( 96*8-1 downto  95*8), 
w97 => Pw(67)( 97*8-1 downto  96*8), w98 => Pw(67)( 98*8-1 downto  97*8), w99 => Pw(67)( 99*8-1 downto  98*8), w100=> Pw(67)(100*8-1 downto  99*8), w101=> Pw(67)(101*8-1 downto 100*8), w102=> Pw(67)(102*8-1 downto 101*8), w103=> Pw(67)(103*8-1 downto 102*8), w104=> Pw(67)(104*8-1 downto 103*8), 
w105=> Pw(67)(105*8-1 downto 104*8), w106=> Pw(67)(106*8-1 downto 105*8), w107=> Pw(67)(107*8-1 downto 106*8), w108=> Pw(67)(108*8-1 downto 107*8), w109=> Pw(67)(109*8-1 downto 108*8), w110=> Pw(67)(110*8-1 downto 109*8), w111=> Pw(67)(111*8-1 downto 110*8), w112=> Pw(67)(112*8-1 downto 111*8), 
w113=> Pw(67)(113*8-1 downto 112*8), w114=> Pw(67)(114*8-1 downto 113*8), w115=> Pw(67)(115*8-1 downto 114*8), w116=> Pw(67)(116*8-1 downto 115*8), w117=> Pw(67)(117*8-1 downto 116*8), w118=> Pw(67)(118*8-1 downto 117*8), w119=> Pw(67)(119*8-1 downto 118*8), w120=> Pw(67)(120*8-1 downto 119*8), 
w121=> Pw(67)(121*8-1 downto 120*8), w122=> Pw(67)(122*8-1 downto 121*8), w123=> Pw(67)(123*8-1 downto 122*8), w124=> Pw(67)(124*8-1 downto 123*8), w125=> Pw(67)(125*8-1 downto 124*8), w126=> Pw(67)(126*8-1 downto 125*8), w127=> Pw(67)(127*8-1 downto 126*8), w128=> Pw(67)(128*8-1 downto 127*8), 
           d_out   => pca_d67_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_68_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(68)(     7 downto    0),   w02 => Pw(68)( 2*8-1 downto    8),   w03 => Pw(68)( 3*8-1 downto  2*8),   w04 => Pw(68)( 4*8-1 downto  3*8),   w05 => Pw(68)( 5*8-1 downto  4*8),   w06 => Pw(68)( 6*8-1 downto  5*8),   w07 => Pw(68)( 7*8-1 downto  6*8),   w08 => Pw(68)( 8*8-1 downto  7*8),  
w09 => Pw(68)( 9*8-1 downto  8*8),   w10 => Pw(68)(10*8-1 downto  9*8),   w11 => Pw(68)(11*8-1 downto 10*8),   w12 => Pw(68)(12*8-1 downto 11*8),   w13 => Pw(68)(13*8-1 downto 12*8),   w14 => Pw(68)(14*8-1 downto 13*8),   w15 => Pw(68)(15*8-1 downto 14*8),   w16 => Pw(68)(16*8-1 downto 15*8),  
w17 => Pw(68)(17*8-1 downto 16*8),   w18 => Pw(68)(18*8-1 downto 17*8),   w19 => Pw(68)(19*8-1 downto 18*8),   w20 => Pw(68)(20*8-1 downto 19*8),   w21 => Pw(68)(21*8-1 downto 20*8),   w22 => Pw(68)(22*8-1 downto 21*8),   w23 => Pw(68)(23*8-1 downto 22*8),   w24 => Pw(68)(24*8-1 downto 23*8),  
w25 => Pw(68)(25*8-1 downto 24*8),   w26 => Pw(68)(26*8-1 downto 25*8),   w27 => Pw(68)(27*8-1 downto 26*8),   w28 => Pw(68)(28*8-1 downto 27*8),   w29 => Pw(68)(29*8-1 downto 28*8),   w30 => Pw(68)(30*8-1 downto 29*8),   w31 => Pw(68)(31*8-1 downto 30*8),   w32 => Pw(68)(32*8-1 downto 31*8),  
w33 => Pw(68)(33*8-1 downto 32*8),   w34 => Pw(68)(34*8-1 downto 33*8),   w35 => Pw(68)(35*8-1 downto 34*8),   w36 => Pw(68)(36*8-1 downto 35*8),   w37 => Pw(68)(37*8-1 downto 36*8),   w38 => Pw(68)(38*8-1 downto 37*8),   w39 => Pw(68)(39*8-1 downto 38*8),   w40 => Pw(68)(40*8-1 downto 39*8),  
w41 => Pw(68)(41*8-1 downto 40*8),   w42 => Pw(68)(42*8-1 downto 41*8),   w43 => Pw(68)(43*8-1 downto 42*8),   w44 => Pw(68)(44*8-1 downto 43*8),   w45 => Pw(68)(45*8-1 downto 44*8),   w46 => Pw(68)(46*8-1 downto 45*8),   w47 => Pw(68)(47*8-1 downto 46*8),   w48 => Pw(68)(48*8-1 downto 47*8),  
w49 => Pw(68)(49*8-1 downto 48*8),   w50 => Pw(68)(50*8-1 downto 49*8),   w51 => Pw(68)(51*8-1 downto 50*8),   w52 => Pw(68)(52*8-1 downto 51*8),   w53 => Pw(68)(53*8-1 downto 52*8),   w54 => Pw(68)(54*8-1 downto 53*8),   w55 => Pw(68)(55*8-1 downto 54*8),   w56 => Pw(68)(56*8-1 downto 55*8),  
w57 => Pw(68)(57*8-1 downto 56*8),   w58 => Pw(68)(58*8-1 downto 57*8),   w59 => Pw(68)(59*8-1 downto 58*8),   w60 => Pw(68)(60*8-1 downto 59*8),   w61 => Pw(68)(61*8-1 downto 60*8),   w62 => Pw(68)(62*8-1 downto 61*8),   w63 => Pw(68)(63*8-1 downto 62*8),   w64 => Pw(68)(64*8-1 downto 63*8), 
w65 => Pw(68)( 65*8-1 downto  64*8), w66 => Pw(68)( 66*8-1 downto  65*8), w67 => Pw(68)( 67*8-1 downto  66*8), w68 => Pw(68)( 68*8-1 downto  67*8), w69 => Pw(68)( 69*8-1 downto  68*8), w70 => Pw(68)( 70*8-1 downto  69*8), w71 => Pw(68)( 71*8-1 downto  70*8), w72 => Pw(68)( 72*8-1 downto  71*8), 
w73 => Pw(68)( 73*8-1 downto  72*8), w74 => Pw(68)( 74*8-1 downto  73*8), w75 => Pw(68)( 75*8-1 downto  74*8), w76 => Pw(68)( 76*8-1 downto  75*8), w77 => Pw(68)( 77*8-1 downto  76*8), w78 => Pw(68)( 78*8-1 downto  77*8), w79 => Pw(68)( 79*8-1 downto  78*8), w80 => Pw(68)( 80*8-1 downto  79*8), 
w81 => Pw(68)( 81*8-1 downto  80*8), w82 => Pw(68)( 82*8-1 downto  81*8), w83 => Pw(68)( 83*8-1 downto  82*8), w84 => Pw(68)( 84*8-1 downto  83*8), w85 => Pw(68)( 85*8-1 downto  84*8), w86 => Pw(68)( 86*8-1 downto  85*8), w87 => Pw(68)( 87*8-1 downto  86*8), w88 => Pw(68)( 88*8-1 downto  87*8), 
w89 => Pw(68)( 89*8-1 downto  88*8), w90 => Pw(68)( 90*8-1 downto  89*8), w91 => Pw(68)( 91*8-1 downto  90*8), w92 => Pw(68)( 92*8-1 downto  91*8), w93 => Pw(68)( 93*8-1 downto  92*8), w94 => Pw(68)( 94*8-1 downto  93*8), w95 => Pw(68)( 95*8-1 downto  94*8), w96 => Pw(68)( 96*8-1 downto  95*8), 
w97 => Pw(68)( 97*8-1 downto  96*8), w98 => Pw(68)( 98*8-1 downto  97*8), w99 => Pw(68)( 99*8-1 downto  98*8), w100=> Pw(68)(100*8-1 downto  99*8), w101=> Pw(68)(101*8-1 downto 100*8), w102=> Pw(68)(102*8-1 downto 101*8), w103=> Pw(68)(103*8-1 downto 102*8), w104=> Pw(68)(104*8-1 downto 103*8), 
w105=> Pw(68)(105*8-1 downto 104*8), w106=> Pw(68)(106*8-1 downto 105*8), w107=> Pw(68)(107*8-1 downto 106*8), w108=> Pw(68)(108*8-1 downto 107*8), w109=> Pw(68)(109*8-1 downto 108*8), w110=> Pw(68)(110*8-1 downto 109*8), w111=> Pw(68)(111*8-1 downto 110*8), w112=> Pw(68)(112*8-1 downto 111*8), 
w113=> Pw(68)(113*8-1 downto 112*8), w114=> Pw(68)(114*8-1 downto 113*8), w115=> Pw(68)(115*8-1 downto 114*8), w116=> Pw(68)(116*8-1 downto 115*8), w117=> Pw(68)(117*8-1 downto 116*8), w118=> Pw(68)(118*8-1 downto 117*8), w119=> Pw(68)(119*8-1 downto 118*8), w120=> Pw(68)(120*8-1 downto 119*8), 
w121=> Pw(68)(121*8-1 downto 120*8), w122=> Pw(68)(122*8-1 downto 121*8), w123=> Pw(68)(123*8-1 downto 122*8), w124=> Pw(68)(124*8-1 downto 123*8), w125=> Pw(68)(125*8-1 downto 124*8), w126=> Pw(68)(126*8-1 downto 125*8), w127=> Pw(68)(127*8-1 downto 126*8), w128=> Pw(68)(128*8-1 downto 127*8), 
           d_out   => pca_d68_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_69_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(69)(     7 downto    0),   w02 => Pw(69)( 2*8-1 downto    8),   w03 => Pw(69)( 3*8-1 downto  2*8),   w04 => Pw(69)( 4*8-1 downto  3*8),   w05 => Pw(69)( 5*8-1 downto  4*8),   w06 => Pw(69)( 6*8-1 downto  5*8),   w07 => Pw(69)( 7*8-1 downto  6*8),   w08 => Pw(69)( 8*8-1 downto  7*8),  
w09 => Pw(69)( 9*8-1 downto  8*8),   w10 => Pw(69)(10*8-1 downto  9*8),   w11 => Pw(69)(11*8-1 downto 10*8),   w12 => Pw(69)(12*8-1 downto 11*8),   w13 => Pw(69)(13*8-1 downto 12*8),   w14 => Pw(69)(14*8-1 downto 13*8),   w15 => Pw(69)(15*8-1 downto 14*8),   w16 => Pw(69)(16*8-1 downto 15*8),  
w17 => Pw(69)(17*8-1 downto 16*8),   w18 => Pw(69)(18*8-1 downto 17*8),   w19 => Pw(69)(19*8-1 downto 18*8),   w20 => Pw(69)(20*8-1 downto 19*8),   w21 => Pw(69)(21*8-1 downto 20*8),   w22 => Pw(69)(22*8-1 downto 21*8),   w23 => Pw(69)(23*8-1 downto 22*8),   w24 => Pw(69)(24*8-1 downto 23*8),  
w25 => Pw(69)(25*8-1 downto 24*8),   w26 => Pw(69)(26*8-1 downto 25*8),   w27 => Pw(69)(27*8-1 downto 26*8),   w28 => Pw(69)(28*8-1 downto 27*8),   w29 => Pw(69)(29*8-1 downto 28*8),   w30 => Pw(69)(30*8-1 downto 29*8),   w31 => Pw(69)(31*8-1 downto 30*8),   w32 => Pw(69)(32*8-1 downto 31*8),  
w33 => Pw(69)(33*8-1 downto 32*8),   w34 => Pw(69)(34*8-1 downto 33*8),   w35 => Pw(69)(35*8-1 downto 34*8),   w36 => Pw(69)(36*8-1 downto 35*8),   w37 => Pw(69)(37*8-1 downto 36*8),   w38 => Pw(69)(38*8-1 downto 37*8),   w39 => Pw(69)(39*8-1 downto 38*8),   w40 => Pw(69)(40*8-1 downto 39*8),  
w41 => Pw(69)(41*8-1 downto 40*8),   w42 => Pw(69)(42*8-1 downto 41*8),   w43 => Pw(69)(43*8-1 downto 42*8),   w44 => Pw(69)(44*8-1 downto 43*8),   w45 => Pw(69)(45*8-1 downto 44*8),   w46 => Pw(69)(46*8-1 downto 45*8),   w47 => Pw(69)(47*8-1 downto 46*8),   w48 => Pw(69)(48*8-1 downto 47*8),  
w49 => Pw(69)(49*8-1 downto 48*8),   w50 => Pw(69)(50*8-1 downto 49*8),   w51 => Pw(69)(51*8-1 downto 50*8),   w52 => Pw(69)(52*8-1 downto 51*8),   w53 => Pw(69)(53*8-1 downto 52*8),   w54 => Pw(69)(54*8-1 downto 53*8),   w55 => Pw(69)(55*8-1 downto 54*8),   w56 => Pw(69)(56*8-1 downto 55*8),  
w57 => Pw(69)(57*8-1 downto 56*8),   w58 => Pw(69)(58*8-1 downto 57*8),   w59 => Pw(69)(59*8-1 downto 58*8),   w60 => Pw(69)(60*8-1 downto 59*8),   w61 => Pw(69)(61*8-1 downto 60*8),   w62 => Pw(69)(62*8-1 downto 61*8),   w63 => Pw(69)(63*8-1 downto 62*8),   w64 => Pw(69)(64*8-1 downto 63*8), 
w65 => Pw(69)( 65*8-1 downto  64*8), w66 => Pw(69)( 66*8-1 downto  65*8), w67 => Pw(69)( 67*8-1 downto  66*8), w68 => Pw(69)( 68*8-1 downto  67*8), w69 => Pw(69)( 69*8-1 downto  68*8), w70 => Pw(69)( 70*8-1 downto  69*8), w71 => Pw(69)( 71*8-1 downto  70*8), w72 => Pw(69)( 72*8-1 downto  71*8), 
w73 => Pw(69)( 73*8-1 downto  72*8), w74 => Pw(69)( 74*8-1 downto  73*8), w75 => Pw(69)( 75*8-1 downto  74*8), w76 => Pw(69)( 76*8-1 downto  75*8), w77 => Pw(69)( 77*8-1 downto  76*8), w78 => Pw(69)( 78*8-1 downto  77*8), w79 => Pw(69)( 79*8-1 downto  78*8), w80 => Pw(69)( 80*8-1 downto  79*8), 
w81 => Pw(69)( 81*8-1 downto  80*8), w82 => Pw(69)( 82*8-1 downto  81*8), w83 => Pw(69)( 83*8-1 downto  82*8), w84 => Pw(69)( 84*8-1 downto  83*8), w85 => Pw(69)( 85*8-1 downto  84*8), w86 => Pw(69)( 86*8-1 downto  85*8), w87 => Pw(69)( 87*8-1 downto  86*8), w88 => Pw(69)( 88*8-1 downto  87*8), 
w89 => Pw(69)( 89*8-1 downto  88*8), w90 => Pw(69)( 90*8-1 downto  89*8), w91 => Pw(69)( 91*8-1 downto  90*8), w92 => Pw(69)( 92*8-1 downto  91*8), w93 => Pw(69)( 93*8-1 downto  92*8), w94 => Pw(69)( 94*8-1 downto  93*8), w95 => Pw(69)( 95*8-1 downto  94*8), w96 => Pw(69)( 96*8-1 downto  95*8), 
w97 => Pw(69)( 97*8-1 downto  96*8), w98 => Pw(69)( 98*8-1 downto  97*8), w99 => Pw(69)( 99*8-1 downto  98*8), w100=> Pw(69)(100*8-1 downto  99*8), w101=> Pw(69)(101*8-1 downto 100*8), w102=> Pw(69)(102*8-1 downto 101*8), w103=> Pw(69)(103*8-1 downto 102*8), w104=> Pw(69)(104*8-1 downto 103*8), 
w105=> Pw(69)(105*8-1 downto 104*8), w106=> Pw(69)(106*8-1 downto 105*8), w107=> Pw(69)(107*8-1 downto 106*8), w108=> Pw(69)(108*8-1 downto 107*8), w109=> Pw(69)(109*8-1 downto 108*8), w110=> Pw(69)(110*8-1 downto 109*8), w111=> Pw(69)(111*8-1 downto 110*8), w112=> Pw(69)(112*8-1 downto 111*8), 
w113=> Pw(69)(113*8-1 downto 112*8), w114=> Pw(69)(114*8-1 downto 113*8), w115=> Pw(69)(115*8-1 downto 114*8), w116=> Pw(69)(116*8-1 downto 115*8), w117=> Pw(69)(117*8-1 downto 116*8), w118=> Pw(69)(118*8-1 downto 117*8), w119=> Pw(69)(119*8-1 downto 118*8), w120=> Pw(69)(120*8-1 downto 119*8), 
w121=> Pw(69)(121*8-1 downto 120*8), w122=> Pw(69)(122*8-1 downto 121*8), w123=> Pw(69)(123*8-1 downto 122*8), w124=> Pw(69)(124*8-1 downto 123*8), w125=> Pw(69)(125*8-1 downto 124*8), w126=> Pw(69)(126*8-1 downto 125*8), w127=> Pw(69)(127*8-1 downto 126*8), w128=> Pw(69)(128*8-1 downto 127*8), 
           d_out   => pca_d69_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_70_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(70)(     7 downto    0),   w02 => Pw(70)( 2*8-1 downto    8),   w03 => Pw(70)( 3*8-1 downto  2*8),   w04 => Pw(70)( 4*8-1 downto  3*8),   w05 => Pw(70)( 5*8-1 downto  4*8),   w06 => Pw(70)( 6*8-1 downto  5*8),   w07 => Pw(70)( 7*8-1 downto  6*8),   w08 => Pw(70)( 8*8-1 downto  7*8),  
w09 => Pw(70)( 9*8-1 downto  8*8),   w10 => Pw(70)(10*8-1 downto  9*8),   w11 => Pw(70)(11*8-1 downto 10*8),   w12 => Pw(70)(12*8-1 downto 11*8),   w13 => Pw(70)(13*8-1 downto 12*8),   w14 => Pw(70)(14*8-1 downto 13*8),   w15 => Pw(70)(15*8-1 downto 14*8),   w16 => Pw(70)(16*8-1 downto 15*8),  
w17 => Pw(70)(17*8-1 downto 16*8),   w18 => Pw(70)(18*8-1 downto 17*8),   w19 => Pw(70)(19*8-1 downto 18*8),   w20 => Pw(70)(20*8-1 downto 19*8),   w21 => Pw(70)(21*8-1 downto 20*8),   w22 => Pw(70)(22*8-1 downto 21*8),   w23 => Pw(70)(23*8-1 downto 22*8),   w24 => Pw(70)(24*8-1 downto 23*8),  
w25 => Pw(70)(25*8-1 downto 24*8),   w26 => Pw(70)(26*8-1 downto 25*8),   w27 => Pw(70)(27*8-1 downto 26*8),   w28 => Pw(70)(28*8-1 downto 27*8),   w29 => Pw(70)(29*8-1 downto 28*8),   w30 => Pw(70)(30*8-1 downto 29*8),   w31 => Pw(70)(31*8-1 downto 30*8),   w32 => Pw(70)(32*8-1 downto 31*8),  
w33 => Pw(70)(33*8-1 downto 32*8),   w34 => Pw(70)(34*8-1 downto 33*8),   w35 => Pw(70)(35*8-1 downto 34*8),   w36 => Pw(70)(36*8-1 downto 35*8),   w37 => Pw(70)(37*8-1 downto 36*8),   w38 => Pw(70)(38*8-1 downto 37*8),   w39 => Pw(70)(39*8-1 downto 38*8),   w40 => Pw(70)(40*8-1 downto 39*8),  
w41 => Pw(70)(41*8-1 downto 40*8),   w42 => Pw(70)(42*8-1 downto 41*8),   w43 => Pw(70)(43*8-1 downto 42*8),   w44 => Pw(70)(44*8-1 downto 43*8),   w45 => Pw(70)(45*8-1 downto 44*8),   w46 => Pw(70)(46*8-1 downto 45*8),   w47 => Pw(70)(47*8-1 downto 46*8),   w48 => Pw(70)(48*8-1 downto 47*8),  
w49 => Pw(70)(49*8-1 downto 48*8),   w50 => Pw(70)(50*8-1 downto 49*8),   w51 => Pw(70)(51*8-1 downto 50*8),   w52 => Pw(70)(52*8-1 downto 51*8),   w53 => Pw(70)(53*8-1 downto 52*8),   w54 => Pw(70)(54*8-1 downto 53*8),   w55 => Pw(70)(55*8-1 downto 54*8),   w56 => Pw(70)(56*8-1 downto 55*8),  
w57 => Pw(70)(57*8-1 downto 56*8),   w58 => Pw(70)(58*8-1 downto 57*8),   w59 => Pw(70)(59*8-1 downto 58*8),   w60 => Pw(70)(60*8-1 downto 59*8),   w61 => Pw(70)(61*8-1 downto 60*8),   w62 => Pw(70)(62*8-1 downto 61*8),   w63 => Pw(70)(63*8-1 downto 62*8),   w64 => Pw(70)(64*8-1 downto 63*8), 
w65 => Pw(70)( 65*8-1 downto  64*8), w66 => Pw(70)( 66*8-1 downto  65*8), w67 => Pw(70)( 67*8-1 downto  66*8), w68 => Pw(70)( 68*8-1 downto  67*8), w69 => Pw(70)( 69*8-1 downto  68*8), w70 => Pw(70)( 70*8-1 downto  69*8), w71 => Pw(70)( 71*8-1 downto  70*8), w72 => Pw(70)( 72*8-1 downto  71*8), 
w73 => Pw(70)( 73*8-1 downto  72*8), w74 => Pw(70)( 74*8-1 downto  73*8), w75 => Pw(70)( 75*8-1 downto  74*8), w76 => Pw(70)( 76*8-1 downto  75*8), w77 => Pw(70)( 77*8-1 downto  76*8), w78 => Pw(70)( 78*8-1 downto  77*8), w79 => Pw(70)( 79*8-1 downto  78*8), w80 => Pw(70)( 80*8-1 downto  79*8), 
w81 => Pw(70)( 81*8-1 downto  80*8), w82 => Pw(70)( 82*8-1 downto  81*8), w83 => Pw(70)( 83*8-1 downto  82*8), w84 => Pw(70)( 84*8-1 downto  83*8), w85 => Pw(70)( 85*8-1 downto  84*8), w86 => Pw(70)( 86*8-1 downto  85*8), w87 => Pw(70)( 87*8-1 downto  86*8), w88 => Pw(70)( 88*8-1 downto  87*8), 
w89 => Pw(70)( 89*8-1 downto  88*8), w90 => Pw(70)( 90*8-1 downto  89*8), w91 => Pw(70)( 91*8-1 downto  90*8), w92 => Pw(70)( 92*8-1 downto  91*8), w93 => Pw(70)( 93*8-1 downto  92*8), w94 => Pw(70)( 94*8-1 downto  93*8), w95 => Pw(70)( 95*8-1 downto  94*8), w96 => Pw(70)( 96*8-1 downto  95*8), 
w97 => Pw(70)( 97*8-1 downto  96*8), w98 => Pw(70)( 98*8-1 downto  97*8), w99 => Pw(70)( 99*8-1 downto  98*8), w100=> Pw(70)(100*8-1 downto  99*8), w101=> Pw(70)(101*8-1 downto 100*8), w102=> Pw(70)(102*8-1 downto 101*8), w103=> Pw(70)(103*8-1 downto 102*8), w104=> Pw(70)(104*8-1 downto 103*8), 
w105=> Pw(70)(105*8-1 downto 104*8), w106=> Pw(70)(106*8-1 downto 105*8), w107=> Pw(70)(107*8-1 downto 106*8), w108=> Pw(70)(108*8-1 downto 107*8), w109=> Pw(70)(109*8-1 downto 108*8), w110=> Pw(70)(110*8-1 downto 109*8), w111=> Pw(70)(111*8-1 downto 110*8), w112=> Pw(70)(112*8-1 downto 111*8), 
w113=> Pw(70)(113*8-1 downto 112*8), w114=> Pw(70)(114*8-1 downto 113*8), w115=> Pw(70)(115*8-1 downto 114*8), w116=> Pw(70)(116*8-1 downto 115*8), w117=> Pw(70)(117*8-1 downto 116*8), w118=> Pw(70)(118*8-1 downto 117*8), w119=> Pw(70)(119*8-1 downto 118*8), w120=> Pw(70)(120*8-1 downto 119*8), 
w121=> Pw(70)(121*8-1 downto 120*8), w122=> Pw(70)(122*8-1 downto 121*8), w123=> Pw(70)(123*8-1 downto 122*8), w124=> Pw(70)(124*8-1 downto 123*8), w125=> Pw(70)(125*8-1 downto 124*8), w126=> Pw(70)(126*8-1 downto 125*8), w127=> Pw(70)(127*8-1 downto 126*8), w128=> Pw(70)(128*8-1 downto 127*8), 
           d_out   => pca_d70_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_71_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(71)(     7 downto    0),   w02 => Pw(71)( 2*8-1 downto    8),   w03 => Pw(71)( 3*8-1 downto  2*8),   w04 => Pw(71)( 4*8-1 downto  3*8),   w05 => Pw(71)( 5*8-1 downto  4*8),   w06 => Pw(71)( 6*8-1 downto  5*8),   w07 => Pw(71)( 7*8-1 downto  6*8),   w08 => Pw(71)( 8*8-1 downto  7*8),  
w09 => Pw(71)( 9*8-1 downto  8*8),   w10 => Pw(71)(10*8-1 downto  9*8),   w11 => Pw(71)(11*8-1 downto 10*8),   w12 => Pw(71)(12*8-1 downto 11*8),   w13 => Pw(71)(13*8-1 downto 12*8),   w14 => Pw(71)(14*8-1 downto 13*8),   w15 => Pw(71)(15*8-1 downto 14*8),   w16 => Pw(71)(16*8-1 downto 15*8),  
w17 => Pw(71)(17*8-1 downto 16*8),   w18 => Pw(71)(18*8-1 downto 17*8),   w19 => Pw(71)(19*8-1 downto 18*8),   w20 => Pw(71)(20*8-1 downto 19*8),   w21 => Pw(71)(21*8-1 downto 20*8),   w22 => Pw(71)(22*8-1 downto 21*8),   w23 => Pw(71)(23*8-1 downto 22*8),   w24 => Pw(71)(24*8-1 downto 23*8),  
w25 => Pw(71)(25*8-1 downto 24*8),   w26 => Pw(71)(26*8-1 downto 25*8),   w27 => Pw(71)(27*8-1 downto 26*8),   w28 => Pw(71)(28*8-1 downto 27*8),   w29 => Pw(71)(29*8-1 downto 28*8),   w30 => Pw(71)(30*8-1 downto 29*8),   w31 => Pw(71)(31*8-1 downto 30*8),   w32 => Pw(71)(32*8-1 downto 31*8),  
w33 => Pw(71)(33*8-1 downto 32*8),   w34 => Pw(71)(34*8-1 downto 33*8),   w35 => Pw(71)(35*8-1 downto 34*8),   w36 => Pw(71)(36*8-1 downto 35*8),   w37 => Pw(71)(37*8-1 downto 36*8),   w38 => Pw(71)(38*8-1 downto 37*8),   w39 => Pw(71)(39*8-1 downto 38*8),   w40 => Pw(71)(40*8-1 downto 39*8),  
w41 => Pw(71)(41*8-1 downto 40*8),   w42 => Pw(71)(42*8-1 downto 41*8),   w43 => Pw(71)(43*8-1 downto 42*8),   w44 => Pw(71)(44*8-1 downto 43*8),   w45 => Pw(71)(45*8-1 downto 44*8),   w46 => Pw(71)(46*8-1 downto 45*8),   w47 => Pw(71)(47*8-1 downto 46*8),   w48 => Pw(71)(48*8-1 downto 47*8),  
w49 => Pw(71)(49*8-1 downto 48*8),   w50 => Pw(71)(50*8-1 downto 49*8),   w51 => Pw(71)(51*8-1 downto 50*8),   w52 => Pw(71)(52*8-1 downto 51*8),   w53 => Pw(71)(53*8-1 downto 52*8),   w54 => Pw(71)(54*8-1 downto 53*8),   w55 => Pw(71)(55*8-1 downto 54*8),   w56 => Pw(71)(56*8-1 downto 55*8),  
w57 => Pw(71)(57*8-1 downto 56*8),   w58 => Pw(71)(58*8-1 downto 57*8),   w59 => Pw(71)(59*8-1 downto 58*8),   w60 => Pw(71)(60*8-1 downto 59*8),   w61 => Pw(71)(61*8-1 downto 60*8),   w62 => Pw(71)(62*8-1 downto 61*8),   w63 => Pw(71)(63*8-1 downto 62*8),   w64 => Pw(71)(64*8-1 downto 63*8), 
w65 => Pw(71)( 65*8-1 downto  64*8), w66 => Pw(71)( 66*8-1 downto  65*8), w67 => Pw(71)( 67*8-1 downto  66*8), w68 => Pw(71)( 68*8-1 downto  67*8), w69 => Pw(71)( 69*8-1 downto  68*8), w70 => Pw(71)( 70*8-1 downto  69*8), w71 => Pw(71)( 71*8-1 downto  70*8), w72 => Pw(71)( 72*8-1 downto  71*8), 
w73 => Pw(71)( 73*8-1 downto  72*8), w74 => Pw(71)( 74*8-1 downto  73*8), w75 => Pw(71)( 75*8-1 downto  74*8), w76 => Pw(71)( 76*8-1 downto  75*8), w77 => Pw(71)( 77*8-1 downto  76*8), w78 => Pw(71)( 78*8-1 downto  77*8), w79 => Pw(71)( 79*8-1 downto  78*8), w80 => Pw(71)( 80*8-1 downto  79*8), 
w81 => Pw(71)( 81*8-1 downto  80*8), w82 => Pw(71)( 82*8-1 downto  81*8), w83 => Pw(71)( 83*8-1 downto  82*8), w84 => Pw(71)( 84*8-1 downto  83*8), w85 => Pw(71)( 85*8-1 downto  84*8), w86 => Pw(71)( 86*8-1 downto  85*8), w87 => Pw(71)( 87*8-1 downto  86*8), w88 => Pw(71)( 88*8-1 downto  87*8), 
w89 => Pw(71)( 89*8-1 downto  88*8), w90 => Pw(71)( 90*8-1 downto  89*8), w91 => Pw(71)( 91*8-1 downto  90*8), w92 => Pw(71)( 92*8-1 downto  91*8), w93 => Pw(71)( 93*8-1 downto  92*8), w94 => Pw(71)( 94*8-1 downto  93*8), w95 => Pw(71)( 95*8-1 downto  94*8), w96 => Pw(71)( 96*8-1 downto  95*8), 
w97 => Pw(71)( 97*8-1 downto  96*8), w98 => Pw(71)( 98*8-1 downto  97*8), w99 => Pw(71)( 99*8-1 downto  98*8), w100=> Pw(71)(100*8-1 downto  99*8), w101=> Pw(71)(101*8-1 downto 100*8), w102=> Pw(71)(102*8-1 downto 101*8), w103=> Pw(71)(103*8-1 downto 102*8), w104=> Pw(71)(104*8-1 downto 103*8), 
w105=> Pw(71)(105*8-1 downto 104*8), w106=> Pw(71)(106*8-1 downto 105*8), w107=> Pw(71)(107*8-1 downto 106*8), w108=> Pw(71)(108*8-1 downto 107*8), w109=> Pw(71)(109*8-1 downto 108*8), w110=> Pw(71)(110*8-1 downto 109*8), w111=> Pw(71)(111*8-1 downto 110*8), w112=> Pw(71)(112*8-1 downto 111*8), 
w113=> Pw(71)(113*8-1 downto 112*8), w114=> Pw(71)(114*8-1 downto 113*8), w115=> Pw(71)(115*8-1 downto 114*8), w116=> Pw(71)(116*8-1 downto 115*8), w117=> Pw(71)(117*8-1 downto 116*8), w118=> Pw(71)(118*8-1 downto 117*8), w119=> Pw(71)(119*8-1 downto 118*8), w120=> Pw(71)(120*8-1 downto 119*8), 
w121=> Pw(71)(121*8-1 downto 120*8), w122=> Pw(71)(122*8-1 downto 121*8), w123=> Pw(71)(123*8-1 downto 122*8), w124=> Pw(71)(124*8-1 downto 123*8), w125=> Pw(71)(125*8-1 downto 124*8), w126=> Pw(71)(126*8-1 downto 125*8), w127=> Pw(71)(127*8-1 downto 126*8), w128=> Pw(71)(128*8-1 downto 127*8), 
           d_out   => pca_d71_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_72_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(72)(     7 downto    0),   w02 => Pw(72)( 2*8-1 downto    8),   w03 => Pw(72)( 3*8-1 downto  2*8),   w04 => Pw(72)( 4*8-1 downto  3*8),   w05 => Pw(72)( 5*8-1 downto  4*8),   w06 => Pw(72)( 6*8-1 downto  5*8),   w07 => Pw(72)( 7*8-1 downto  6*8),   w08 => Pw(72)( 8*8-1 downto  7*8),  
w09 => Pw(72)( 9*8-1 downto  8*8),   w10 => Pw(72)(10*8-1 downto  9*8),   w11 => Pw(72)(11*8-1 downto 10*8),   w12 => Pw(72)(12*8-1 downto 11*8),   w13 => Pw(72)(13*8-1 downto 12*8),   w14 => Pw(72)(14*8-1 downto 13*8),   w15 => Pw(72)(15*8-1 downto 14*8),   w16 => Pw(72)(16*8-1 downto 15*8),  
w17 => Pw(72)(17*8-1 downto 16*8),   w18 => Pw(72)(18*8-1 downto 17*8),   w19 => Pw(72)(19*8-1 downto 18*8),   w20 => Pw(72)(20*8-1 downto 19*8),   w21 => Pw(72)(21*8-1 downto 20*8),   w22 => Pw(72)(22*8-1 downto 21*8),   w23 => Pw(72)(23*8-1 downto 22*8),   w24 => Pw(72)(24*8-1 downto 23*8),  
w25 => Pw(72)(25*8-1 downto 24*8),   w26 => Pw(72)(26*8-1 downto 25*8),   w27 => Pw(72)(27*8-1 downto 26*8),   w28 => Pw(72)(28*8-1 downto 27*8),   w29 => Pw(72)(29*8-1 downto 28*8),   w30 => Pw(72)(30*8-1 downto 29*8),   w31 => Pw(72)(31*8-1 downto 30*8),   w32 => Pw(72)(32*8-1 downto 31*8),  
w33 => Pw(72)(33*8-1 downto 32*8),   w34 => Pw(72)(34*8-1 downto 33*8),   w35 => Pw(72)(35*8-1 downto 34*8),   w36 => Pw(72)(36*8-1 downto 35*8),   w37 => Pw(72)(37*8-1 downto 36*8),   w38 => Pw(72)(38*8-1 downto 37*8),   w39 => Pw(72)(39*8-1 downto 38*8),   w40 => Pw(72)(40*8-1 downto 39*8),  
w41 => Pw(72)(41*8-1 downto 40*8),   w42 => Pw(72)(42*8-1 downto 41*8),   w43 => Pw(72)(43*8-1 downto 42*8),   w44 => Pw(72)(44*8-1 downto 43*8),   w45 => Pw(72)(45*8-1 downto 44*8),   w46 => Pw(72)(46*8-1 downto 45*8),   w47 => Pw(72)(47*8-1 downto 46*8),   w48 => Pw(72)(48*8-1 downto 47*8),  
w49 => Pw(72)(49*8-1 downto 48*8),   w50 => Pw(72)(50*8-1 downto 49*8),   w51 => Pw(72)(51*8-1 downto 50*8),   w52 => Pw(72)(52*8-1 downto 51*8),   w53 => Pw(72)(53*8-1 downto 52*8),   w54 => Pw(72)(54*8-1 downto 53*8),   w55 => Pw(72)(55*8-1 downto 54*8),   w56 => Pw(72)(56*8-1 downto 55*8),  
w57 => Pw(72)(57*8-1 downto 56*8),   w58 => Pw(72)(58*8-1 downto 57*8),   w59 => Pw(72)(59*8-1 downto 58*8),   w60 => Pw(72)(60*8-1 downto 59*8),   w61 => Pw(72)(61*8-1 downto 60*8),   w62 => Pw(72)(62*8-1 downto 61*8),   w63 => Pw(72)(63*8-1 downto 62*8),   w64 => Pw(72)(64*8-1 downto 63*8), 
w65 => Pw(72)( 65*8-1 downto  64*8), w66 => Pw(72)( 66*8-1 downto  65*8), w67 => Pw(72)( 67*8-1 downto  66*8), w68 => Pw(72)( 68*8-1 downto  67*8), w69 => Pw(72)( 69*8-1 downto  68*8), w70 => Pw(72)( 70*8-1 downto  69*8), w71 => Pw(72)( 71*8-1 downto  70*8), w72 => Pw(72)( 72*8-1 downto  71*8), 
w73 => Pw(72)( 73*8-1 downto  72*8), w74 => Pw(72)( 74*8-1 downto  73*8), w75 => Pw(72)( 75*8-1 downto  74*8), w76 => Pw(72)( 76*8-1 downto  75*8), w77 => Pw(72)( 77*8-1 downto  76*8), w78 => Pw(72)( 78*8-1 downto  77*8), w79 => Pw(72)( 79*8-1 downto  78*8), w80 => Pw(72)( 80*8-1 downto  79*8), 
w81 => Pw(72)( 81*8-1 downto  80*8), w82 => Pw(72)( 82*8-1 downto  81*8), w83 => Pw(72)( 83*8-1 downto  82*8), w84 => Pw(72)( 84*8-1 downto  83*8), w85 => Pw(72)( 85*8-1 downto  84*8), w86 => Pw(72)( 86*8-1 downto  85*8), w87 => Pw(72)( 87*8-1 downto  86*8), w88 => Pw(72)( 88*8-1 downto  87*8), 
w89 => Pw(72)( 89*8-1 downto  88*8), w90 => Pw(72)( 90*8-1 downto  89*8), w91 => Pw(72)( 91*8-1 downto  90*8), w92 => Pw(72)( 92*8-1 downto  91*8), w93 => Pw(72)( 93*8-1 downto  92*8), w94 => Pw(72)( 94*8-1 downto  93*8), w95 => Pw(72)( 95*8-1 downto  94*8), w96 => Pw(72)( 96*8-1 downto  95*8), 
w97 => Pw(72)( 97*8-1 downto  96*8), w98 => Pw(72)( 98*8-1 downto  97*8), w99 => Pw(72)( 99*8-1 downto  98*8), w100=> Pw(72)(100*8-1 downto  99*8), w101=> Pw(72)(101*8-1 downto 100*8), w102=> Pw(72)(102*8-1 downto 101*8), w103=> Pw(72)(103*8-1 downto 102*8), w104=> Pw(72)(104*8-1 downto 103*8), 
w105=> Pw(72)(105*8-1 downto 104*8), w106=> Pw(72)(106*8-1 downto 105*8), w107=> Pw(72)(107*8-1 downto 106*8), w108=> Pw(72)(108*8-1 downto 107*8), w109=> Pw(72)(109*8-1 downto 108*8), w110=> Pw(72)(110*8-1 downto 109*8), w111=> Pw(72)(111*8-1 downto 110*8), w112=> Pw(72)(112*8-1 downto 111*8), 
w113=> Pw(72)(113*8-1 downto 112*8), w114=> Pw(72)(114*8-1 downto 113*8), w115=> Pw(72)(115*8-1 downto 114*8), w116=> Pw(72)(116*8-1 downto 115*8), w117=> Pw(72)(117*8-1 downto 116*8), w118=> Pw(72)(118*8-1 downto 117*8), w119=> Pw(72)(119*8-1 downto 118*8), w120=> Pw(72)(120*8-1 downto 119*8), 
w121=> Pw(72)(121*8-1 downto 120*8), w122=> Pw(72)(122*8-1 downto 121*8), w123=> Pw(72)(123*8-1 downto 122*8), w124=> Pw(72)(124*8-1 downto 123*8), w125=> Pw(72)(125*8-1 downto 124*8), w126=> Pw(72)(126*8-1 downto 125*8), w127=> Pw(72)(127*8-1 downto 126*8), w128=> Pw(72)(128*8-1 downto 127*8), 
           d_out   => pca_d72_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_73_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(73)(     7 downto    0),   w02 => Pw(73)( 2*8-1 downto    8),   w03 => Pw(73)( 3*8-1 downto  2*8),   w04 => Pw(73)( 4*8-1 downto  3*8),   w05 => Pw(73)( 5*8-1 downto  4*8),   w06 => Pw(73)( 6*8-1 downto  5*8),   w07 => Pw(73)( 7*8-1 downto  6*8),   w08 => Pw(73)( 8*8-1 downto  7*8),  
w09 => Pw(73)( 9*8-1 downto  8*8),   w10 => Pw(73)(10*8-1 downto  9*8),   w11 => Pw(73)(11*8-1 downto 10*8),   w12 => Pw(73)(12*8-1 downto 11*8),   w13 => Pw(73)(13*8-1 downto 12*8),   w14 => Pw(73)(14*8-1 downto 13*8),   w15 => Pw(73)(15*8-1 downto 14*8),   w16 => Pw(73)(16*8-1 downto 15*8),  
w17 => Pw(73)(17*8-1 downto 16*8),   w18 => Pw(73)(18*8-1 downto 17*8),   w19 => Pw(73)(19*8-1 downto 18*8),   w20 => Pw(73)(20*8-1 downto 19*8),   w21 => Pw(73)(21*8-1 downto 20*8),   w22 => Pw(73)(22*8-1 downto 21*8),   w23 => Pw(73)(23*8-1 downto 22*8),   w24 => Pw(73)(24*8-1 downto 23*8),  
w25 => Pw(73)(25*8-1 downto 24*8),   w26 => Pw(73)(26*8-1 downto 25*8),   w27 => Pw(73)(27*8-1 downto 26*8),   w28 => Pw(73)(28*8-1 downto 27*8),   w29 => Pw(73)(29*8-1 downto 28*8),   w30 => Pw(73)(30*8-1 downto 29*8),   w31 => Pw(73)(31*8-1 downto 30*8),   w32 => Pw(73)(32*8-1 downto 31*8),  
w33 => Pw(73)(33*8-1 downto 32*8),   w34 => Pw(73)(34*8-1 downto 33*8),   w35 => Pw(73)(35*8-1 downto 34*8),   w36 => Pw(73)(36*8-1 downto 35*8),   w37 => Pw(73)(37*8-1 downto 36*8),   w38 => Pw(73)(38*8-1 downto 37*8),   w39 => Pw(73)(39*8-1 downto 38*8),   w40 => Pw(73)(40*8-1 downto 39*8),  
w41 => Pw(73)(41*8-1 downto 40*8),   w42 => Pw(73)(42*8-1 downto 41*8),   w43 => Pw(73)(43*8-1 downto 42*8),   w44 => Pw(73)(44*8-1 downto 43*8),   w45 => Pw(73)(45*8-1 downto 44*8),   w46 => Pw(73)(46*8-1 downto 45*8),   w47 => Pw(73)(47*8-1 downto 46*8),   w48 => Pw(73)(48*8-1 downto 47*8),  
w49 => Pw(73)(49*8-1 downto 48*8),   w50 => Pw(73)(50*8-1 downto 49*8),   w51 => Pw(73)(51*8-1 downto 50*8),   w52 => Pw(73)(52*8-1 downto 51*8),   w53 => Pw(73)(53*8-1 downto 52*8),   w54 => Pw(73)(54*8-1 downto 53*8),   w55 => Pw(73)(55*8-1 downto 54*8),   w56 => Pw(73)(56*8-1 downto 55*8),  
w57 => Pw(73)(57*8-1 downto 56*8),   w58 => Pw(73)(58*8-1 downto 57*8),   w59 => Pw(73)(59*8-1 downto 58*8),   w60 => Pw(73)(60*8-1 downto 59*8),   w61 => Pw(73)(61*8-1 downto 60*8),   w62 => Pw(73)(62*8-1 downto 61*8),   w63 => Pw(73)(63*8-1 downto 62*8),   w64 => Pw(73)(64*8-1 downto 63*8), 
w65 => Pw(73)( 65*8-1 downto  64*8), w66 => Pw(73)( 66*8-1 downto  65*8), w67 => Pw(73)( 67*8-1 downto  66*8), w68 => Pw(73)( 68*8-1 downto  67*8), w69 => Pw(73)( 69*8-1 downto  68*8), w70 => Pw(73)( 70*8-1 downto  69*8), w71 => Pw(73)( 71*8-1 downto  70*8), w72 => Pw(73)( 72*8-1 downto  71*8), 
w73 => Pw(73)( 73*8-1 downto  72*8), w74 => Pw(73)( 74*8-1 downto  73*8), w75 => Pw(73)( 75*8-1 downto  74*8), w76 => Pw(73)( 76*8-1 downto  75*8), w77 => Pw(73)( 77*8-1 downto  76*8), w78 => Pw(73)( 78*8-1 downto  77*8), w79 => Pw(73)( 79*8-1 downto  78*8), w80 => Pw(73)( 80*8-1 downto  79*8), 
w81 => Pw(73)( 81*8-1 downto  80*8), w82 => Pw(73)( 82*8-1 downto  81*8), w83 => Pw(73)( 83*8-1 downto  82*8), w84 => Pw(73)( 84*8-1 downto  83*8), w85 => Pw(73)( 85*8-1 downto  84*8), w86 => Pw(73)( 86*8-1 downto  85*8), w87 => Pw(73)( 87*8-1 downto  86*8), w88 => Pw(73)( 88*8-1 downto  87*8), 
w89 => Pw(73)( 89*8-1 downto  88*8), w90 => Pw(73)( 90*8-1 downto  89*8), w91 => Pw(73)( 91*8-1 downto  90*8), w92 => Pw(73)( 92*8-1 downto  91*8), w93 => Pw(73)( 93*8-1 downto  92*8), w94 => Pw(73)( 94*8-1 downto  93*8), w95 => Pw(73)( 95*8-1 downto  94*8), w96 => Pw(73)( 96*8-1 downto  95*8), 
w97 => Pw(73)( 97*8-1 downto  96*8), w98 => Pw(73)( 98*8-1 downto  97*8), w99 => Pw(73)( 99*8-1 downto  98*8), w100=> Pw(73)(100*8-1 downto  99*8), w101=> Pw(73)(101*8-1 downto 100*8), w102=> Pw(73)(102*8-1 downto 101*8), w103=> Pw(73)(103*8-1 downto 102*8), w104=> Pw(73)(104*8-1 downto 103*8), 
w105=> Pw(73)(105*8-1 downto 104*8), w106=> Pw(73)(106*8-1 downto 105*8), w107=> Pw(73)(107*8-1 downto 106*8), w108=> Pw(73)(108*8-1 downto 107*8), w109=> Pw(73)(109*8-1 downto 108*8), w110=> Pw(73)(110*8-1 downto 109*8), w111=> Pw(73)(111*8-1 downto 110*8), w112=> Pw(73)(112*8-1 downto 111*8), 
w113=> Pw(73)(113*8-1 downto 112*8), w114=> Pw(73)(114*8-1 downto 113*8), w115=> Pw(73)(115*8-1 downto 114*8), w116=> Pw(73)(116*8-1 downto 115*8), w117=> Pw(73)(117*8-1 downto 116*8), w118=> Pw(73)(118*8-1 downto 117*8), w119=> Pw(73)(119*8-1 downto 118*8), w120=> Pw(73)(120*8-1 downto 119*8), 
w121=> Pw(73)(121*8-1 downto 120*8), w122=> Pw(73)(122*8-1 downto 121*8), w123=> Pw(73)(123*8-1 downto 122*8), w124=> Pw(73)(124*8-1 downto 123*8), w125=> Pw(73)(125*8-1 downto 124*8), w126=> Pw(73)(126*8-1 downto 125*8), w127=> Pw(73)(127*8-1 downto 126*8), w128=> Pw(73)(128*8-1 downto 127*8), 
           d_out   => pca_d73_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_74_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(74)(     7 downto    0),   w02 => Pw(74)( 2*8-1 downto    8),   w03 => Pw(74)( 3*8-1 downto  2*8),   w04 => Pw(74)( 4*8-1 downto  3*8),   w05 => Pw(74)( 5*8-1 downto  4*8),   w06 => Pw(74)( 6*8-1 downto  5*8),   w07 => Pw(74)( 7*8-1 downto  6*8),   w08 => Pw(74)( 8*8-1 downto  7*8),  
w09 => Pw(74)( 9*8-1 downto  8*8),   w10 => Pw(74)(10*8-1 downto  9*8),   w11 => Pw(74)(11*8-1 downto 10*8),   w12 => Pw(74)(12*8-1 downto 11*8),   w13 => Pw(74)(13*8-1 downto 12*8),   w14 => Pw(74)(14*8-1 downto 13*8),   w15 => Pw(74)(15*8-1 downto 14*8),   w16 => Pw(74)(16*8-1 downto 15*8),  
w17 => Pw(74)(17*8-1 downto 16*8),   w18 => Pw(74)(18*8-1 downto 17*8),   w19 => Pw(74)(19*8-1 downto 18*8),   w20 => Pw(74)(20*8-1 downto 19*8),   w21 => Pw(74)(21*8-1 downto 20*8),   w22 => Pw(74)(22*8-1 downto 21*8),   w23 => Pw(74)(23*8-1 downto 22*8),   w24 => Pw(74)(24*8-1 downto 23*8),  
w25 => Pw(74)(25*8-1 downto 24*8),   w26 => Pw(74)(26*8-1 downto 25*8),   w27 => Pw(74)(27*8-1 downto 26*8),   w28 => Pw(74)(28*8-1 downto 27*8),   w29 => Pw(74)(29*8-1 downto 28*8),   w30 => Pw(74)(30*8-1 downto 29*8),   w31 => Pw(74)(31*8-1 downto 30*8),   w32 => Pw(74)(32*8-1 downto 31*8),  
w33 => Pw(74)(33*8-1 downto 32*8),   w34 => Pw(74)(34*8-1 downto 33*8),   w35 => Pw(74)(35*8-1 downto 34*8),   w36 => Pw(74)(36*8-1 downto 35*8),   w37 => Pw(74)(37*8-1 downto 36*8),   w38 => Pw(74)(38*8-1 downto 37*8),   w39 => Pw(74)(39*8-1 downto 38*8),   w40 => Pw(74)(40*8-1 downto 39*8),  
w41 => Pw(74)(41*8-1 downto 40*8),   w42 => Pw(74)(42*8-1 downto 41*8),   w43 => Pw(74)(43*8-1 downto 42*8),   w44 => Pw(74)(44*8-1 downto 43*8),   w45 => Pw(74)(45*8-1 downto 44*8),   w46 => Pw(74)(46*8-1 downto 45*8),   w47 => Pw(74)(47*8-1 downto 46*8),   w48 => Pw(74)(48*8-1 downto 47*8),  
w49 => Pw(74)(49*8-1 downto 48*8),   w50 => Pw(74)(50*8-1 downto 49*8),   w51 => Pw(74)(51*8-1 downto 50*8),   w52 => Pw(74)(52*8-1 downto 51*8),   w53 => Pw(74)(53*8-1 downto 52*8),   w54 => Pw(74)(54*8-1 downto 53*8),   w55 => Pw(74)(55*8-1 downto 54*8),   w56 => Pw(74)(56*8-1 downto 55*8),  
w57 => Pw(74)(57*8-1 downto 56*8),   w58 => Pw(74)(58*8-1 downto 57*8),   w59 => Pw(74)(59*8-1 downto 58*8),   w60 => Pw(74)(60*8-1 downto 59*8),   w61 => Pw(74)(61*8-1 downto 60*8),   w62 => Pw(74)(62*8-1 downto 61*8),   w63 => Pw(74)(63*8-1 downto 62*8),   w64 => Pw(74)(64*8-1 downto 63*8), 
w65 => Pw(74)( 65*8-1 downto  64*8), w66 => Pw(74)( 66*8-1 downto  65*8), w67 => Pw(74)( 67*8-1 downto  66*8), w68 => Pw(74)( 68*8-1 downto  67*8), w69 => Pw(74)( 69*8-1 downto  68*8), w70 => Pw(74)( 70*8-1 downto  69*8), w71 => Pw(74)( 71*8-1 downto  70*8), w72 => Pw(74)( 72*8-1 downto  71*8), 
w73 => Pw(74)( 73*8-1 downto  72*8), w74 => Pw(74)( 74*8-1 downto  73*8), w75 => Pw(74)( 75*8-1 downto  74*8), w76 => Pw(74)( 76*8-1 downto  75*8), w77 => Pw(74)( 77*8-1 downto  76*8), w78 => Pw(74)( 78*8-1 downto  77*8), w79 => Pw(74)( 79*8-1 downto  78*8), w80 => Pw(74)( 80*8-1 downto  79*8), 
w81 => Pw(74)( 81*8-1 downto  80*8), w82 => Pw(74)( 82*8-1 downto  81*8), w83 => Pw(74)( 83*8-1 downto  82*8), w84 => Pw(74)( 84*8-1 downto  83*8), w85 => Pw(74)( 85*8-1 downto  84*8), w86 => Pw(74)( 86*8-1 downto  85*8), w87 => Pw(74)( 87*8-1 downto  86*8), w88 => Pw(74)( 88*8-1 downto  87*8), 
w89 => Pw(74)( 89*8-1 downto  88*8), w90 => Pw(74)( 90*8-1 downto  89*8), w91 => Pw(74)( 91*8-1 downto  90*8), w92 => Pw(74)( 92*8-1 downto  91*8), w93 => Pw(74)( 93*8-1 downto  92*8), w94 => Pw(74)( 94*8-1 downto  93*8), w95 => Pw(74)( 95*8-1 downto  94*8), w96 => Pw(74)( 96*8-1 downto  95*8), 
w97 => Pw(74)( 97*8-1 downto  96*8), w98 => Pw(74)( 98*8-1 downto  97*8), w99 => Pw(74)( 99*8-1 downto  98*8), w100=> Pw(74)(100*8-1 downto  99*8), w101=> Pw(74)(101*8-1 downto 100*8), w102=> Pw(74)(102*8-1 downto 101*8), w103=> Pw(74)(103*8-1 downto 102*8), w104=> Pw(74)(104*8-1 downto 103*8), 
w105=> Pw(74)(105*8-1 downto 104*8), w106=> Pw(74)(106*8-1 downto 105*8), w107=> Pw(74)(107*8-1 downto 106*8), w108=> Pw(74)(108*8-1 downto 107*8), w109=> Pw(74)(109*8-1 downto 108*8), w110=> Pw(74)(110*8-1 downto 109*8), w111=> Pw(74)(111*8-1 downto 110*8), w112=> Pw(74)(112*8-1 downto 111*8), 
w113=> Pw(74)(113*8-1 downto 112*8), w114=> Pw(74)(114*8-1 downto 113*8), w115=> Pw(74)(115*8-1 downto 114*8), w116=> Pw(74)(116*8-1 downto 115*8), w117=> Pw(74)(117*8-1 downto 116*8), w118=> Pw(74)(118*8-1 downto 117*8), w119=> Pw(74)(119*8-1 downto 118*8), w120=> Pw(74)(120*8-1 downto 119*8), 
w121=> Pw(74)(121*8-1 downto 120*8), w122=> Pw(74)(122*8-1 downto 121*8), w123=> Pw(74)(123*8-1 downto 122*8), w124=> Pw(74)(124*8-1 downto 123*8), w125=> Pw(74)(125*8-1 downto 124*8), w126=> Pw(74)(126*8-1 downto 125*8), w127=> Pw(74)(127*8-1 downto 126*8), w128=> Pw(74)(128*8-1 downto 127*8), 
           d_out   => pca_d74_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_75_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(75)(     7 downto    0),   w02 => Pw(75)( 2*8-1 downto    8),   w03 => Pw(75)( 3*8-1 downto  2*8),   w04 => Pw(75)( 4*8-1 downto  3*8),   w05 => Pw(75)( 5*8-1 downto  4*8),   w06 => Pw(75)( 6*8-1 downto  5*8),   w07 => Pw(75)( 7*8-1 downto  6*8),   w08 => Pw(75)( 8*8-1 downto  7*8),  
w09 => Pw(75)( 9*8-1 downto  8*8),   w10 => Pw(75)(10*8-1 downto  9*8),   w11 => Pw(75)(11*8-1 downto 10*8),   w12 => Pw(75)(12*8-1 downto 11*8),   w13 => Pw(75)(13*8-1 downto 12*8),   w14 => Pw(75)(14*8-1 downto 13*8),   w15 => Pw(75)(15*8-1 downto 14*8),   w16 => Pw(75)(16*8-1 downto 15*8),  
w17 => Pw(75)(17*8-1 downto 16*8),   w18 => Pw(75)(18*8-1 downto 17*8),   w19 => Pw(75)(19*8-1 downto 18*8),   w20 => Pw(75)(20*8-1 downto 19*8),   w21 => Pw(75)(21*8-1 downto 20*8),   w22 => Pw(75)(22*8-1 downto 21*8),   w23 => Pw(75)(23*8-1 downto 22*8),   w24 => Pw(75)(24*8-1 downto 23*8),  
w25 => Pw(75)(25*8-1 downto 24*8),   w26 => Pw(75)(26*8-1 downto 25*8),   w27 => Pw(75)(27*8-1 downto 26*8),   w28 => Pw(75)(28*8-1 downto 27*8),   w29 => Pw(75)(29*8-1 downto 28*8),   w30 => Pw(75)(30*8-1 downto 29*8),   w31 => Pw(75)(31*8-1 downto 30*8),   w32 => Pw(75)(32*8-1 downto 31*8),  
w33 => Pw(75)(33*8-1 downto 32*8),   w34 => Pw(75)(34*8-1 downto 33*8),   w35 => Pw(75)(35*8-1 downto 34*8),   w36 => Pw(75)(36*8-1 downto 35*8),   w37 => Pw(75)(37*8-1 downto 36*8),   w38 => Pw(75)(38*8-1 downto 37*8),   w39 => Pw(75)(39*8-1 downto 38*8),   w40 => Pw(75)(40*8-1 downto 39*8),  
w41 => Pw(75)(41*8-1 downto 40*8),   w42 => Pw(75)(42*8-1 downto 41*8),   w43 => Pw(75)(43*8-1 downto 42*8),   w44 => Pw(75)(44*8-1 downto 43*8),   w45 => Pw(75)(45*8-1 downto 44*8),   w46 => Pw(75)(46*8-1 downto 45*8),   w47 => Pw(75)(47*8-1 downto 46*8),   w48 => Pw(75)(48*8-1 downto 47*8),  
w49 => Pw(75)(49*8-1 downto 48*8),   w50 => Pw(75)(50*8-1 downto 49*8),   w51 => Pw(75)(51*8-1 downto 50*8),   w52 => Pw(75)(52*8-1 downto 51*8),   w53 => Pw(75)(53*8-1 downto 52*8),   w54 => Pw(75)(54*8-1 downto 53*8),   w55 => Pw(75)(55*8-1 downto 54*8),   w56 => Pw(75)(56*8-1 downto 55*8),  
w57 => Pw(75)(57*8-1 downto 56*8),   w58 => Pw(75)(58*8-1 downto 57*8),   w59 => Pw(75)(59*8-1 downto 58*8),   w60 => Pw(75)(60*8-1 downto 59*8),   w61 => Pw(75)(61*8-1 downto 60*8),   w62 => Pw(75)(62*8-1 downto 61*8),   w63 => Pw(75)(63*8-1 downto 62*8),   w64 => Pw(75)(64*8-1 downto 63*8), 
w65 => Pw(75)( 65*8-1 downto  64*8), w66 => Pw(75)( 66*8-1 downto  65*8), w67 => Pw(75)( 67*8-1 downto  66*8), w68 => Pw(75)( 68*8-1 downto  67*8), w69 => Pw(75)( 69*8-1 downto  68*8), w70 => Pw(75)( 70*8-1 downto  69*8), w71 => Pw(75)( 71*8-1 downto  70*8), w72 => Pw(75)( 72*8-1 downto  71*8), 
w73 => Pw(75)( 73*8-1 downto  72*8), w74 => Pw(75)( 74*8-1 downto  73*8), w75 => Pw(75)( 75*8-1 downto  74*8), w76 => Pw(75)( 76*8-1 downto  75*8), w77 => Pw(75)( 77*8-1 downto  76*8), w78 => Pw(75)( 78*8-1 downto  77*8), w79 => Pw(75)( 79*8-1 downto  78*8), w80 => Pw(75)( 80*8-1 downto  79*8), 
w81 => Pw(75)( 81*8-1 downto  80*8), w82 => Pw(75)( 82*8-1 downto  81*8), w83 => Pw(75)( 83*8-1 downto  82*8), w84 => Pw(75)( 84*8-1 downto  83*8), w85 => Pw(75)( 85*8-1 downto  84*8), w86 => Pw(75)( 86*8-1 downto  85*8), w87 => Pw(75)( 87*8-1 downto  86*8), w88 => Pw(75)( 88*8-1 downto  87*8), 
w89 => Pw(75)( 89*8-1 downto  88*8), w90 => Pw(75)( 90*8-1 downto  89*8), w91 => Pw(75)( 91*8-1 downto  90*8), w92 => Pw(75)( 92*8-1 downto  91*8), w93 => Pw(75)( 93*8-1 downto  92*8), w94 => Pw(75)( 94*8-1 downto  93*8), w95 => Pw(75)( 95*8-1 downto  94*8), w96 => Pw(75)( 96*8-1 downto  95*8), 
w97 => Pw(75)( 97*8-1 downto  96*8), w98 => Pw(75)( 98*8-1 downto  97*8), w99 => Pw(75)( 99*8-1 downto  98*8), w100=> Pw(75)(100*8-1 downto  99*8), w101=> Pw(75)(101*8-1 downto 100*8), w102=> Pw(75)(102*8-1 downto 101*8), w103=> Pw(75)(103*8-1 downto 102*8), w104=> Pw(75)(104*8-1 downto 103*8), 
w105=> Pw(75)(105*8-1 downto 104*8), w106=> Pw(75)(106*8-1 downto 105*8), w107=> Pw(75)(107*8-1 downto 106*8), w108=> Pw(75)(108*8-1 downto 107*8), w109=> Pw(75)(109*8-1 downto 108*8), w110=> Pw(75)(110*8-1 downto 109*8), w111=> Pw(75)(111*8-1 downto 110*8), w112=> Pw(75)(112*8-1 downto 111*8), 
w113=> Pw(75)(113*8-1 downto 112*8), w114=> Pw(75)(114*8-1 downto 113*8), w115=> Pw(75)(115*8-1 downto 114*8), w116=> Pw(75)(116*8-1 downto 115*8), w117=> Pw(75)(117*8-1 downto 116*8), w118=> Pw(75)(118*8-1 downto 117*8), w119=> Pw(75)(119*8-1 downto 118*8), w120=> Pw(75)(120*8-1 downto 119*8), 
w121=> Pw(75)(121*8-1 downto 120*8), w122=> Pw(75)(122*8-1 downto 121*8), w123=> Pw(75)(123*8-1 downto 122*8), w124=> Pw(75)(124*8-1 downto 123*8), w125=> Pw(75)(125*8-1 downto 124*8), w126=> Pw(75)(126*8-1 downto 125*8), w127=> Pw(75)(127*8-1 downto 126*8), w128=> Pw(75)(128*8-1 downto 127*8), 
           d_out   => pca_d75_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_76_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(76)(     7 downto    0),   w02 => Pw(76)( 2*8-1 downto    8),   w03 => Pw(76)( 3*8-1 downto  2*8),   w04 => Pw(76)( 4*8-1 downto  3*8),   w05 => Pw(76)( 5*8-1 downto  4*8),   w06 => Pw(76)( 6*8-1 downto  5*8),   w07 => Pw(76)( 7*8-1 downto  6*8),   w08 => Pw(76)( 8*8-1 downto  7*8),  
w09 => Pw(76)( 9*8-1 downto  8*8),   w10 => Pw(76)(10*8-1 downto  9*8),   w11 => Pw(76)(11*8-1 downto 10*8),   w12 => Pw(76)(12*8-1 downto 11*8),   w13 => Pw(76)(13*8-1 downto 12*8),   w14 => Pw(76)(14*8-1 downto 13*8),   w15 => Pw(76)(15*8-1 downto 14*8),   w16 => Pw(76)(16*8-1 downto 15*8),  
w17 => Pw(76)(17*8-1 downto 16*8),   w18 => Pw(76)(18*8-1 downto 17*8),   w19 => Pw(76)(19*8-1 downto 18*8),   w20 => Pw(76)(20*8-1 downto 19*8),   w21 => Pw(76)(21*8-1 downto 20*8),   w22 => Pw(76)(22*8-1 downto 21*8),   w23 => Pw(76)(23*8-1 downto 22*8),   w24 => Pw(76)(24*8-1 downto 23*8),  
w25 => Pw(76)(25*8-1 downto 24*8),   w26 => Pw(76)(26*8-1 downto 25*8),   w27 => Pw(76)(27*8-1 downto 26*8),   w28 => Pw(76)(28*8-1 downto 27*8),   w29 => Pw(76)(29*8-1 downto 28*8),   w30 => Pw(76)(30*8-1 downto 29*8),   w31 => Pw(76)(31*8-1 downto 30*8),   w32 => Pw(76)(32*8-1 downto 31*8),  
w33 => Pw(76)(33*8-1 downto 32*8),   w34 => Pw(76)(34*8-1 downto 33*8),   w35 => Pw(76)(35*8-1 downto 34*8),   w36 => Pw(76)(36*8-1 downto 35*8),   w37 => Pw(76)(37*8-1 downto 36*8),   w38 => Pw(76)(38*8-1 downto 37*8),   w39 => Pw(76)(39*8-1 downto 38*8),   w40 => Pw(76)(40*8-1 downto 39*8),  
w41 => Pw(76)(41*8-1 downto 40*8),   w42 => Pw(76)(42*8-1 downto 41*8),   w43 => Pw(76)(43*8-1 downto 42*8),   w44 => Pw(76)(44*8-1 downto 43*8),   w45 => Pw(76)(45*8-1 downto 44*8),   w46 => Pw(76)(46*8-1 downto 45*8),   w47 => Pw(76)(47*8-1 downto 46*8),   w48 => Pw(76)(48*8-1 downto 47*8),  
w49 => Pw(76)(49*8-1 downto 48*8),   w50 => Pw(76)(50*8-1 downto 49*8),   w51 => Pw(76)(51*8-1 downto 50*8),   w52 => Pw(76)(52*8-1 downto 51*8),   w53 => Pw(76)(53*8-1 downto 52*8),   w54 => Pw(76)(54*8-1 downto 53*8),   w55 => Pw(76)(55*8-1 downto 54*8),   w56 => Pw(76)(56*8-1 downto 55*8),  
w57 => Pw(76)(57*8-1 downto 56*8),   w58 => Pw(76)(58*8-1 downto 57*8),   w59 => Pw(76)(59*8-1 downto 58*8),   w60 => Pw(76)(60*8-1 downto 59*8),   w61 => Pw(76)(61*8-1 downto 60*8),   w62 => Pw(76)(62*8-1 downto 61*8),   w63 => Pw(76)(63*8-1 downto 62*8),   w64 => Pw(76)(64*8-1 downto 63*8), 
w65 => Pw(76)( 65*8-1 downto  64*8), w66 => Pw(76)( 66*8-1 downto  65*8), w67 => Pw(76)( 67*8-1 downto  66*8), w68 => Pw(76)( 68*8-1 downto  67*8), w69 => Pw(76)( 69*8-1 downto  68*8), w70 => Pw(76)( 70*8-1 downto  69*8), w71 => Pw(76)( 71*8-1 downto  70*8), w72 => Pw(76)( 72*8-1 downto  71*8), 
w73 => Pw(76)( 73*8-1 downto  72*8), w74 => Pw(76)( 74*8-1 downto  73*8), w75 => Pw(76)( 75*8-1 downto  74*8), w76 => Pw(76)( 76*8-1 downto  75*8), w77 => Pw(76)( 77*8-1 downto  76*8), w78 => Pw(76)( 78*8-1 downto  77*8), w79 => Pw(76)( 79*8-1 downto  78*8), w80 => Pw(76)( 80*8-1 downto  79*8), 
w81 => Pw(76)( 81*8-1 downto  80*8), w82 => Pw(76)( 82*8-1 downto  81*8), w83 => Pw(76)( 83*8-1 downto  82*8), w84 => Pw(76)( 84*8-1 downto  83*8), w85 => Pw(76)( 85*8-1 downto  84*8), w86 => Pw(76)( 86*8-1 downto  85*8), w87 => Pw(76)( 87*8-1 downto  86*8), w88 => Pw(76)( 88*8-1 downto  87*8), 
w89 => Pw(76)( 89*8-1 downto  88*8), w90 => Pw(76)( 90*8-1 downto  89*8), w91 => Pw(76)( 91*8-1 downto  90*8), w92 => Pw(76)( 92*8-1 downto  91*8), w93 => Pw(76)( 93*8-1 downto  92*8), w94 => Pw(76)( 94*8-1 downto  93*8), w95 => Pw(76)( 95*8-1 downto  94*8), w96 => Pw(76)( 96*8-1 downto  95*8), 
w97 => Pw(76)( 97*8-1 downto  96*8), w98 => Pw(76)( 98*8-1 downto  97*8), w99 => Pw(76)( 99*8-1 downto  98*8), w100=> Pw(76)(100*8-1 downto  99*8), w101=> Pw(76)(101*8-1 downto 100*8), w102=> Pw(76)(102*8-1 downto 101*8), w103=> Pw(76)(103*8-1 downto 102*8), w104=> Pw(76)(104*8-1 downto 103*8), 
w105=> Pw(76)(105*8-1 downto 104*8), w106=> Pw(76)(106*8-1 downto 105*8), w107=> Pw(76)(107*8-1 downto 106*8), w108=> Pw(76)(108*8-1 downto 107*8), w109=> Pw(76)(109*8-1 downto 108*8), w110=> Pw(76)(110*8-1 downto 109*8), w111=> Pw(76)(111*8-1 downto 110*8), w112=> Pw(76)(112*8-1 downto 111*8), 
w113=> Pw(76)(113*8-1 downto 112*8), w114=> Pw(76)(114*8-1 downto 113*8), w115=> Pw(76)(115*8-1 downto 114*8), w116=> Pw(76)(116*8-1 downto 115*8), w117=> Pw(76)(117*8-1 downto 116*8), w118=> Pw(76)(118*8-1 downto 117*8), w119=> Pw(76)(119*8-1 downto 118*8), w120=> Pw(76)(120*8-1 downto 119*8), 
w121=> Pw(76)(121*8-1 downto 120*8), w122=> Pw(76)(122*8-1 downto 121*8), w123=> Pw(76)(123*8-1 downto 122*8), w124=> Pw(76)(124*8-1 downto 123*8), w125=> Pw(76)(125*8-1 downto 124*8), w126=> Pw(76)(126*8-1 downto 125*8), w127=> Pw(76)(127*8-1 downto 126*8), w128=> Pw(76)(128*8-1 downto 127*8), 
           d_out   => pca_d76_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_77_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(77)(     7 downto    0),   w02 => Pw(77)( 2*8-1 downto    8),   w03 => Pw(77)( 3*8-1 downto  2*8),   w04 => Pw(77)( 4*8-1 downto  3*8),   w05 => Pw(77)( 5*8-1 downto  4*8),   w06 => Pw(77)( 6*8-1 downto  5*8),   w07 => Pw(77)( 7*8-1 downto  6*8),   w08 => Pw(77)( 8*8-1 downto  7*8),  
w09 => Pw(77)( 9*8-1 downto  8*8),   w10 => Pw(77)(10*8-1 downto  9*8),   w11 => Pw(77)(11*8-1 downto 10*8),   w12 => Pw(77)(12*8-1 downto 11*8),   w13 => Pw(77)(13*8-1 downto 12*8),   w14 => Pw(77)(14*8-1 downto 13*8),   w15 => Pw(77)(15*8-1 downto 14*8),   w16 => Pw(77)(16*8-1 downto 15*8),  
w17 => Pw(77)(17*8-1 downto 16*8),   w18 => Pw(77)(18*8-1 downto 17*8),   w19 => Pw(77)(19*8-1 downto 18*8),   w20 => Pw(77)(20*8-1 downto 19*8),   w21 => Pw(77)(21*8-1 downto 20*8),   w22 => Pw(77)(22*8-1 downto 21*8),   w23 => Pw(77)(23*8-1 downto 22*8),   w24 => Pw(77)(24*8-1 downto 23*8),  
w25 => Pw(77)(25*8-1 downto 24*8),   w26 => Pw(77)(26*8-1 downto 25*8),   w27 => Pw(77)(27*8-1 downto 26*8),   w28 => Pw(77)(28*8-1 downto 27*8),   w29 => Pw(77)(29*8-1 downto 28*8),   w30 => Pw(77)(30*8-1 downto 29*8),   w31 => Pw(77)(31*8-1 downto 30*8),   w32 => Pw(77)(32*8-1 downto 31*8),  
w33 => Pw(77)(33*8-1 downto 32*8),   w34 => Pw(77)(34*8-1 downto 33*8),   w35 => Pw(77)(35*8-1 downto 34*8),   w36 => Pw(77)(36*8-1 downto 35*8),   w37 => Pw(77)(37*8-1 downto 36*8),   w38 => Pw(77)(38*8-1 downto 37*8),   w39 => Pw(77)(39*8-1 downto 38*8),   w40 => Pw(77)(40*8-1 downto 39*8),  
w41 => Pw(77)(41*8-1 downto 40*8),   w42 => Pw(77)(42*8-1 downto 41*8),   w43 => Pw(77)(43*8-1 downto 42*8),   w44 => Pw(77)(44*8-1 downto 43*8),   w45 => Pw(77)(45*8-1 downto 44*8),   w46 => Pw(77)(46*8-1 downto 45*8),   w47 => Pw(77)(47*8-1 downto 46*8),   w48 => Pw(77)(48*8-1 downto 47*8),  
w49 => Pw(77)(49*8-1 downto 48*8),   w50 => Pw(77)(50*8-1 downto 49*8),   w51 => Pw(77)(51*8-1 downto 50*8),   w52 => Pw(77)(52*8-1 downto 51*8),   w53 => Pw(77)(53*8-1 downto 52*8),   w54 => Pw(77)(54*8-1 downto 53*8),   w55 => Pw(77)(55*8-1 downto 54*8),   w56 => Pw(77)(56*8-1 downto 55*8),  
w57 => Pw(77)(57*8-1 downto 56*8),   w58 => Pw(77)(58*8-1 downto 57*8),   w59 => Pw(77)(59*8-1 downto 58*8),   w60 => Pw(77)(60*8-1 downto 59*8),   w61 => Pw(77)(61*8-1 downto 60*8),   w62 => Pw(77)(62*8-1 downto 61*8),   w63 => Pw(77)(63*8-1 downto 62*8),   w64 => Pw(77)(64*8-1 downto 63*8), 
w65 => Pw(77)( 65*8-1 downto  64*8), w66 => Pw(77)( 66*8-1 downto  65*8), w67 => Pw(77)( 67*8-1 downto  66*8), w68 => Pw(77)( 68*8-1 downto  67*8), w69 => Pw(77)( 69*8-1 downto  68*8), w70 => Pw(77)( 70*8-1 downto  69*8), w71 => Pw(77)( 71*8-1 downto  70*8), w72 => Pw(77)( 72*8-1 downto  71*8), 
w73 => Pw(77)( 73*8-1 downto  72*8), w74 => Pw(77)( 74*8-1 downto  73*8), w75 => Pw(77)( 75*8-1 downto  74*8), w76 => Pw(77)( 76*8-1 downto  75*8), w77 => Pw(77)( 77*8-1 downto  76*8), w78 => Pw(77)( 78*8-1 downto  77*8), w79 => Pw(77)( 79*8-1 downto  78*8), w80 => Pw(77)( 80*8-1 downto  79*8), 
w81 => Pw(77)( 81*8-1 downto  80*8), w82 => Pw(77)( 82*8-1 downto  81*8), w83 => Pw(77)( 83*8-1 downto  82*8), w84 => Pw(77)( 84*8-1 downto  83*8), w85 => Pw(77)( 85*8-1 downto  84*8), w86 => Pw(77)( 86*8-1 downto  85*8), w87 => Pw(77)( 87*8-1 downto  86*8), w88 => Pw(77)( 88*8-1 downto  87*8), 
w89 => Pw(77)( 89*8-1 downto  88*8), w90 => Pw(77)( 90*8-1 downto  89*8), w91 => Pw(77)( 91*8-1 downto  90*8), w92 => Pw(77)( 92*8-1 downto  91*8), w93 => Pw(77)( 93*8-1 downto  92*8), w94 => Pw(77)( 94*8-1 downto  93*8), w95 => Pw(77)( 95*8-1 downto  94*8), w96 => Pw(77)( 96*8-1 downto  95*8), 
w97 => Pw(77)( 97*8-1 downto  96*8), w98 => Pw(77)( 98*8-1 downto  97*8), w99 => Pw(77)( 99*8-1 downto  98*8), w100=> Pw(77)(100*8-1 downto  99*8), w101=> Pw(77)(101*8-1 downto 100*8), w102=> Pw(77)(102*8-1 downto 101*8), w103=> Pw(77)(103*8-1 downto 102*8), w104=> Pw(77)(104*8-1 downto 103*8), 
w105=> Pw(77)(105*8-1 downto 104*8), w106=> Pw(77)(106*8-1 downto 105*8), w107=> Pw(77)(107*8-1 downto 106*8), w108=> Pw(77)(108*8-1 downto 107*8), w109=> Pw(77)(109*8-1 downto 108*8), w110=> Pw(77)(110*8-1 downto 109*8), w111=> Pw(77)(111*8-1 downto 110*8), w112=> Pw(77)(112*8-1 downto 111*8), 
w113=> Pw(77)(113*8-1 downto 112*8), w114=> Pw(77)(114*8-1 downto 113*8), w115=> Pw(77)(115*8-1 downto 114*8), w116=> Pw(77)(116*8-1 downto 115*8), w117=> Pw(77)(117*8-1 downto 116*8), w118=> Pw(77)(118*8-1 downto 117*8), w119=> Pw(77)(119*8-1 downto 118*8), w120=> Pw(77)(120*8-1 downto 119*8), 
w121=> Pw(77)(121*8-1 downto 120*8), w122=> Pw(77)(122*8-1 downto 121*8), w123=> Pw(77)(123*8-1 downto 122*8), w124=> Pw(77)(124*8-1 downto 123*8), w125=> Pw(77)(125*8-1 downto 124*8), w126=> Pw(77)(126*8-1 downto 125*8), w127=> Pw(77)(127*8-1 downto 126*8), w128=> Pw(77)(128*8-1 downto 127*8), 
           d_out   => pca_d77_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_78_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(78)(     7 downto    0),   w02 => Pw(78)( 2*8-1 downto    8),   w03 => Pw(78)( 3*8-1 downto  2*8),   w04 => Pw(78)( 4*8-1 downto  3*8),   w05 => Pw(78)( 5*8-1 downto  4*8),   w06 => Pw(78)( 6*8-1 downto  5*8),   w07 => Pw(78)( 7*8-1 downto  6*8),   w08 => Pw(78)( 8*8-1 downto  7*8),  
w09 => Pw(78)( 9*8-1 downto  8*8),   w10 => Pw(78)(10*8-1 downto  9*8),   w11 => Pw(78)(11*8-1 downto 10*8),   w12 => Pw(78)(12*8-1 downto 11*8),   w13 => Pw(78)(13*8-1 downto 12*8),   w14 => Pw(78)(14*8-1 downto 13*8),   w15 => Pw(78)(15*8-1 downto 14*8),   w16 => Pw(78)(16*8-1 downto 15*8),  
w17 => Pw(78)(17*8-1 downto 16*8),   w18 => Pw(78)(18*8-1 downto 17*8),   w19 => Pw(78)(19*8-1 downto 18*8),   w20 => Pw(78)(20*8-1 downto 19*8),   w21 => Pw(78)(21*8-1 downto 20*8),   w22 => Pw(78)(22*8-1 downto 21*8),   w23 => Pw(78)(23*8-1 downto 22*8),   w24 => Pw(78)(24*8-1 downto 23*8),  
w25 => Pw(78)(25*8-1 downto 24*8),   w26 => Pw(78)(26*8-1 downto 25*8),   w27 => Pw(78)(27*8-1 downto 26*8),   w28 => Pw(78)(28*8-1 downto 27*8),   w29 => Pw(78)(29*8-1 downto 28*8),   w30 => Pw(78)(30*8-1 downto 29*8),   w31 => Pw(78)(31*8-1 downto 30*8),   w32 => Pw(78)(32*8-1 downto 31*8),  
w33 => Pw(78)(33*8-1 downto 32*8),   w34 => Pw(78)(34*8-1 downto 33*8),   w35 => Pw(78)(35*8-1 downto 34*8),   w36 => Pw(78)(36*8-1 downto 35*8),   w37 => Pw(78)(37*8-1 downto 36*8),   w38 => Pw(78)(38*8-1 downto 37*8),   w39 => Pw(78)(39*8-1 downto 38*8),   w40 => Pw(78)(40*8-1 downto 39*8),  
w41 => Pw(78)(41*8-1 downto 40*8),   w42 => Pw(78)(42*8-1 downto 41*8),   w43 => Pw(78)(43*8-1 downto 42*8),   w44 => Pw(78)(44*8-1 downto 43*8),   w45 => Pw(78)(45*8-1 downto 44*8),   w46 => Pw(78)(46*8-1 downto 45*8),   w47 => Pw(78)(47*8-1 downto 46*8),   w48 => Pw(78)(48*8-1 downto 47*8),  
w49 => Pw(78)(49*8-1 downto 48*8),   w50 => Pw(78)(50*8-1 downto 49*8),   w51 => Pw(78)(51*8-1 downto 50*8),   w52 => Pw(78)(52*8-1 downto 51*8),   w53 => Pw(78)(53*8-1 downto 52*8),   w54 => Pw(78)(54*8-1 downto 53*8),   w55 => Pw(78)(55*8-1 downto 54*8),   w56 => Pw(78)(56*8-1 downto 55*8),  
w57 => Pw(78)(57*8-1 downto 56*8),   w58 => Pw(78)(58*8-1 downto 57*8),   w59 => Pw(78)(59*8-1 downto 58*8),   w60 => Pw(78)(60*8-1 downto 59*8),   w61 => Pw(78)(61*8-1 downto 60*8),   w62 => Pw(78)(62*8-1 downto 61*8),   w63 => Pw(78)(63*8-1 downto 62*8),   w64 => Pw(78)(64*8-1 downto 63*8), 
w65 => Pw(78)( 65*8-1 downto  64*8), w66 => Pw(78)( 66*8-1 downto  65*8), w67 => Pw(78)( 67*8-1 downto  66*8), w68 => Pw(78)( 68*8-1 downto  67*8), w69 => Pw(78)( 69*8-1 downto  68*8), w70 => Pw(78)( 70*8-1 downto  69*8), w71 => Pw(78)( 71*8-1 downto  70*8), w72 => Pw(78)( 72*8-1 downto  71*8), 
w73 => Pw(78)( 73*8-1 downto  72*8), w74 => Pw(78)( 74*8-1 downto  73*8), w75 => Pw(78)( 75*8-1 downto  74*8), w76 => Pw(78)( 76*8-1 downto  75*8), w77 => Pw(78)( 77*8-1 downto  76*8), w78 => Pw(78)( 78*8-1 downto  77*8), w79 => Pw(78)( 79*8-1 downto  78*8), w80 => Pw(78)( 80*8-1 downto  79*8), 
w81 => Pw(78)( 81*8-1 downto  80*8), w82 => Pw(78)( 82*8-1 downto  81*8), w83 => Pw(78)( 83*8-1 downto  82*8), w84 => Pw(78)( 84*8-1 downto  83*8), w85 => Pw(78)( 85*8-1 downto  84*8), w86 => Pw(78)( 86*8-1 downto  85*8), w87 => Pw(78)( 87*8-1 downto  86*8), w88 => Pw(78)( 88*8-1 downto  87*8), 
w89 => Pw(78)( 89*8-1 downto  88*8), w90 => Pw(78)( 90*8-1 downto  89*8), w91 => Pw(78)( 91*8-1 downto  90*8), w92 => Pw(78)( 92*8-1 downto  91*8), w93 => Pw(78)( 93*8-1 downto  92*8), w94 => Pw(78)( 94*8-1 downto  93*8), w95 => Pw(78)( 95*8-1 downto  94*8), w96 => Pw(78)( 96*8-1 downto  95*8), 
w97 => Pw(78)( 97*8-1 downto  96*8), w98 => Pw(78)( 98*8-1 downto  97*8), w99 => Pw(78)( 99*8-1 downto  98*8), w100=> Pw(78)(100*8-1 downto  99*8), w101=> Pw(78)(101*8-1 downto 100*8), w102=> Pw(78)(102*8-1 downto 101*8), w103=> Pw(78)(103*8-1 downto 102*8), w104=> Pw(78)(104*8-1 downto 103*8), 
w105=> Pw(78)(105*8-1 downto 104*8), w106=> Pw(78)(106*8-1 downto 105*8), w107=> Pw(78)(107*8-1 downto 106*8), w108=> Pw(78)(108*8-1 downto 107*8), w109=> Pw(78)(109*8-1 downto 108*8), w110=> Pw(78)(110*8-1 downto 109*8), w111=> Pw(78)(111*8-1 downto 110*8), w112=> Pw(78)(112*8-1 downto 111*8), 
w113=> Pw(78)(113*8-1 downto 112*8), w114=> Pw(78)(114*8-1 downto 113*8), w115=> Pw(78)(115*8-1 downto 114*8), w116=> Pw(78)(116*8-1 downto 115*8), w117=> Pw(78)(117*8-1 downto 116*8), w118=> Pw(78)(118*8-1 downto 117*8), w119=> Pw(78)(119*8-1 downto 118*8), w120=> Pw(78)(120*8-1 downto 119*8), 
w121=> Pw(78)(121*8-1 downto 120*8), w122=> Pw(78)(122*8-1 downto 121*8), w123=> Pw(78)(123*8-1 downto 122*8), w124=> Pw(78)(124*8-1 downto 123*8), w125=> Pw(78)(125*8-1 downto 124*8), w126=> Pw(78)(126*8-1 downto 125*8), w127=> Pw(78)(127*8-1 downto 126*8), w128=> Pw(78)(128*8-1 downto 127*8), 
           d_out   => pca_d78_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_79_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(79)(     7 downto    0),   w02 => Pw(79)( 2*8-1 downto    8),   w03 => Pw(79)( 3*8-1 downto  2*8),   w04 => Pw(79)( 4*8-1 downto  3*8),   w05 => Pw(79)( 5*8-1 downto  4*8),   w06 => Pw(79)( 6*8-1 downto  5*8),   w07 => Pw(79)( 7*8-1 downto  6*8),   w08 => Pw(79)( 8*8-1 downto  7*8),  
w09 => Pw(79)( 9*8-1 downto  8*8),   w10 => Pw(79)(10*8-1 downto  9*8),   w11 => Pw(79)(11*8-1 downto 10*8),   w12 => Pw(79)(12*8-1 downto 11*8),   w13 => Pw(79)(13*8-1 downto 12*8),   w14 => Pw(79)(14*8-1 downto 13*8),   w15 => Pw(79)(15*8-1 downto 14*8),   w16 => Pw(79)(16*8-1 downto 15*8),  
w17 => Pw(79)(17*8-1 downto 16*8),   w18 => Pw(79)(18*8-1 downto 17*8),   w19 => Pw(79)(19*8-1 downto 18*8),   w20 => Pw(79)(20*8-1 downto 19*8),   w21 => Pw(79)(21*8-1 downto 20*8),   w22 => Pw(79)(22*8-1 downto 21*8),   w23 => Pw(79)(23*8-1 downto 22*8),   w24 => Pw(79)(24*8-1 downto 23*8),  
w25 => Pw(79)(25*8-1 downto 24*8),   w26 => Pw(79)(26*8-1 downto 25*8),   w27 => Pw(79)(27*8-1 downto 26*8),   w28 => Pw(79)(28*8-1 downto 27*8),   w29 => Pw(79)(29*8-1 downto 28*8),   w30 => Pw(79)(30*8-1 downto 29*8),   w31 => Pw(79)(31*8-1 downto 30*8),   w32 => Pw(79)(32*8-1 downto 31*8),  
w33 => Pw(79)(33*8-1 downto 32*8),   w34 => Pw(79)(34*8-1 downto 33*8),   w35 => Pw(79)(35*8-1 downto 34*8),   w36 => Pw(79)(36*8-1 downto 35*8),   w37 => Pw(79)(37*8-1 downto 36*8),   w38 => Pw(79)(38*8-1 downto 37*8),   w39 => Pw(79)(39*8-1 downto 38*8),   w40 => Pw(79)(40*8-1 downto 39*8),  
w41 => Pw(79)(41*8-1 downto 40*8),   w42 => Pw(79)(42*8-1 downto 41*8),   w43 => Pw(79)(43*8-1 downto 42*8),   w44 => Pw(79)(44*8-1 downto 43*8),   w45 => Pw(79)(45*8-1 downto 44*8),   w46 => Pw(79)(46*8-1 downto 45*8),   w47 => Pw(79)(47*8-1 downto 46*8),   w48 => Pw(79)(48*8-1 downto 47*8),  
w49 => Pw(79)(49*8-1 downto 48*8),   w50 => Pw(79)(50*8-1 downto 49*8),   w51 => Pw(79)(51*8-1 downto 50*8),   w52 => Pw(79)(52*8-1 downto 51*8),   w53 => Pw(79)(53*8-1 downto 52*8),   w54 => Pw(79)(54*8-1 downto 53*8),   w55 => Pw(79)(55*8-1 downto 54*8),   w56 => Pw(79)(56*8-1 downto 55*8),  
w57 => Pw(79)(57*8-1 downto 56*8),   w58 => Pw(79)(58*8-1 downto 57*8),   w59 => Pw(79)(59*8-1 downto 58*8),   w60 => Pw(79)(60*8-1 downto 59*8),   w61 => Pw(79)(61*8-1 downto 60*8),   w62 => Pw(79)(62*8-1 downto 61*8),   w63 => Pw(79)(63*8-1 downto 62*8),   w64 => Pw(79)(64*8-1 downto 63*8), 
w65 => Pw(79)( 65*8-1 downto  64*8), w66 => Pw(79)( 66*8-1 downto  65*8), w67 => Pw(79)( 67*8-1 downto  66*8), w68 => Pw(79)( 68*8-1 downto  67*8), w69 => Pw(79)( 69*8-1 downto  68*8), w70 => Pw(79)( 70*8-1 downto  69*8), w71 => Pw(79)( 71*8-1 downto  70*8), w72 => Pw(79)( 72*8-1 downto  71*8), 
w73 => Pw(79)( 73*8-1 downto  72*8), w74 => Pw(79)( 74*8-1 downto  73*8), w75 => Pw(79)( 75*8-1 downto  74*8), w76 => Pw(79)( 76*8-1 downto  75*8), w77 => Pw(79)( 77*8-1 downto  76*8), w78 => Pw(79)( 78*8-1 downto  77*8), w79 => Pw(79)( 79*8-1 downto  78*8), w80 => Pw(79)( 80*8-1 downto  79*8), 
w81 => Pw(79)( 81*8-1 downto  80*8), w82 => Pw(79)( 82*8-1 downto  81*8), w83 => Pw(79)( 83*8-1 downto  82*8), w84 => Pw(79)( 84*8-1 downto  83*8), w85 => Pw(79)( 85*8-1 downto  84*8), w86 => Pw(79)( 86*8-1 downto  85*8), w87 => Pw(79)( 87*8-1 downto  86*8), w88 => Pw(79)( 88*8-1 downto  87*8), 
w89 => Pw(79)( 89*8-1 downto  88*8), w90 => Pw(79)( 90*8-1 downto  89*8), w91 => Pw(79)( 91*8-1 downto  90*8), w92 => Pw(79)( 92*8-1 downto  91*8), w93 => Pw(79)( 93*8-1 downto  92*8), w94 => Pw(79)( 94*8-1 downto  93*8), w95 => Pw(79)( 95*8-1 downto  94*8), w96 => Pw(79)( 96*8-1 downto  95*8), 
w97 => Pw(79)( 97*8-1 downto  96*8), w98 => Pw(79)( 98*8-1 downto  97*8), w99 => Pw(79)( 99*8-1 downto  98*8), w100=> Pw(79)(100*8-1 downto  99*8), w101=> Pw(79)(101*8-1 downto 100*8), w102=> Pw(79)(102*8-1 downto 101*8), w103=> Pw(79)(103*8-1 downto 102*8), w104=> Pw(79)(104*8-1 downto 103*8), 
w105=> Pw(79)(105*8-1 downto 104*8), w106=> Pw(79)(106*8-1 downto 105*8), w107=> Pw(79)(107*8-1 downto 106*8), w108=> Pw(79)(108*8-1 downto 107*8), w109=> Pw(79)(109*8-1 downto 108*8), w110=> Pw(79)(110*8-1 downto 109*8), w111=> Pw(79)(111*8-1 downto 110*8), w112=> Pw(79)(112*8-1 downto 111*8), 
w113=> Pw(79)(113*8-1 downto 112*8), w114=> Pw(79)(114*8-1 downto 113*8), w115=> Pw(79)(115*8-1 downto 114*8), w116=> Pw(79)(116*8-1 downto 115*8), w117=> Pw(79)(117*8-1 downto 116*8), w118=> Pw(79)(118*8-1 downto 117*8), w119=> Pw(79)(119*8-1 downto 118*8), w120=> Pw(79)(120*8-1 downto 119*8), 
w121=> Pw(79)(121*8-1 downto 120*8), w122=> Pw(79)(122*8-1 downto 121*8), w123=> Pw(79)(123*8-1 downto 122*8), w124=> Pw(79)(124*8-1 downto 123*8), w125=> Pw(79)(125*8-1 downto 124*8), w126=> Pw(79)(126*8-1 downto 125*8), w127=> Pw(79)(127*8-1 downto 126*8), w128=> Pw(79)(128*8-1 downto 127*8), 
           d_out   => pca_d79_out   ,
           en_out  => open  ,
           sof_out => open );

  PCA128_80_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(80)(     7 downto    0),   w02 => Pw(80)( 2*8-1 downto    8),   w03 => Pw(80)( 3*8-1 downto  2*8),   w04 => Pw(80)( 4*8-1 downto  3*8),   w05 => Pw(80)( 5*8-1 downto  4*8),   w06 => Pw(80)( 6*8-1 downto  5*8),   w07 => Pw(80)( 7*8-1 downto  6*8),   w08 => Pw(80)( 8*8-1 downto  7*8),  
w09 => Pw(80)( 9*8-1 downto  8*8),   w10 => Pw(80)(10*8-1 downto  9*8),   w11 => Pw(80)(11*8-1 downto 10*8),   w12 => Pw(80)(12*8-1 downto 11*8),   w13 => Pw(80)(13*8-1 downto 12*8),   w14 => Pw(80)(14*8-1 downto 13*8),   w15 => Pw(80)(15*8-1 downto 14*8),   w16 => Pw(80)(16*8-1 downto 15*8),  
w17 => Pw(80)(17*8-1 downto 16*8),   w18 => Pw(80)(18*8-1 downto 17*8),   w19 => Pw(80)(19*8-1 downto 18*8),   w20 => Pw(80)(20*8-1 downto 19*8),   w21 => Pw(80)(21*8-1 downto 20*8),   w22 => Pw(80)(22*8-1 downto 21*8),   w23 => Pw(80)(23*8-1 downto 22*8),   w24 => Pw(80)(24*8-1 downto 23*8),  
w25 => Pw(80)(25*8-1 downto 24*8),   w26 => Pw(80)(26*8-1 downto 25*8),   w27 => Pw(80)(27*8-1 downto 26*8),   w28 => Pw(80)(28*8-1 downto 27*8),   w29 => Pw(80)(29*8-1 downto 28*8),   w30 => Pw(80)(30*8-1 downto 29*8),   w31 => Pw(80)(31*8-1 downto 30*8),   w32 => Pw(80)(32*8-1 downto 31*8),  
w33 => Pw(80)(33*8-1 downto 32*8),   w34 => Pw(80)(34*8-1 downto 33*8),   w35 => Pw(80)(35*8-1 downto 34*8),   w36 => Pw(80)(36*8-1 downto 35*8),   w37 => Pw(80)(37*8-1 downto 36*8),   w38 => Pw(80)(38*8-1 downto 37*8),   w39 => Pw(80)(39*8-1 downto 38*8),   w40 => Pw(80)(40*8-1 downto 39*8),  
w41 => Pw(80)(41*8-1 downto 40*8),   w42 => Pw(80)(42*8-1 downto 41*8),   w43 => Pw(80)(43*8-1 downto 42*8),   w44 => Pw(80)(44*8-1 downto 43*8),   w45 => Pw(80)(45*8-1 downto 44*8),   w46 => Pw(80)(46*8-1 downto 45*8),   w47 => Pw(80)(47*8-1 downto 46*8),   w48 => Pw(80)(48*8-1 downto 47*8),  
w49 => Pw(80)(49*8-1 downto 48*8),   w50 => Pw(80)(50*8-1 downto 49*8),   w51 => Pw(80)(51*8-1 downto 50*8),   w52 => Pw(80)(52*8-1 downto 51*8),   w53 => Pw(80)(53*8-1 downto 52*8),   w54 => Pw(80)(54*8-1 downto 53*8),   w55 => Pw(80)(55*8-1 downto 54*8),   w56 => Pw(80)(56*8-1 downto 55*8),  
w57 => Pw(80)(57*8-1 downto 56*8),   w58 => Pw(80)(58*8-1 downto 57*8),   w59 => Pw(80)(59*8-1 downto 58*8),   w60 => Pw(80)(60*8-1 downto 59*8),   w61 => Pw(80)(61*8-1 downto 60*8),   w62 => Pw(80)(62*8-1 downto 61*8),   w63 => Pw(80)(63*8-1 downto 62*8),   w64 => Pw(80)(64*8-1 downto 63*8), 
w65 => Pw(80)( 65*8-1 downto  64*8), w66 => Pw(80)( 66*8-1 downto  65*8), w67 => Pw(80)( 67*8-1 downto  66*8), w68 => Pw(80)( 68*8-1 downto  67*8), w69 => Pw(80)( 69*8-1 downto  68*8), w70 => Pw(80)( 70*8-1 downto  69*8), w71 => Pw(80)( 71*8-1 downto  70*8), w72 => Pw(80)( 72*8-1 downto  71*8), 
w73 => Pw(80)( 73*8-1 downto  72*8), w74 => Pw(80)( 74*8-1 downto  73*8), w75 => Pw(80)( 75*8-1 downto  74*8), w76 => Pw(80)( 76*8-1 downto  75*8), w77 => Pw(80)( 77*8-1 downto  76*8), w78 => Pw(80)( 78*8-1 downto  77*8), w79 => Pw(80)( 79*8-1 downto  78*8), w80 => Pw(80)( 80*8-1 downto  79*8), 
w81 => Pw(80)( 81*8-1 downto  80*8), w82 => Pw(80)( 82*8-1 downto  81*8), w83 => Pw(80)( 83*8-1 downto  82*8), w84 => Pw(80)( 84*8-1 downto  83*8), w85 => Pw(80)( 85*8-1 downto  84*8), w86 => Pw(80)( 86*8-1 downto  85*8), w87 => Pw(80)( 87*8-1 downto  86*8), w88 => Pw(80)( 88*8-1 downto  87*8), 
w89 => Pw(80)( 89*8-1 downto  88*8), w90 => Pw(80)( 90*8-1 downto  89*8), w91 => Pw(80)( 91*8-1 downto  90*8), w92 => Pw(80)( 92*8-1 downto  91*8), w93 => Pw(80)( 93*8-1 downto  92*8), w94 => Pw(80)( 94*8-1 downto  93*8), w95 => Pw(80)( 95*8-1 downto  94*8), w96 => Pw(80)( 96*8-1 downto  95*8), 
w97 => Pw(80)( 97*8-1 downto  96*8), w98 => Pw(80)( 98*8-1 downto  97*8), w99 => Pw(80)( 99*8-1 downto  98*8), w100=> Pw(80)(100*8-1 downto  99*8), w101=> Pw(80)(101*8-1 downto 100*8), w102=> Pw(80)(102*8-1 downto 101*8), w103=> Pw(80)(103*8-1 downto 102*8), w104=> Pw(80)(104*8-1 downto 103*8), 
w105=> Pw(80)(105*8-1 downto 104*8), w106=> Pw(80)(106*8-1 downto 105*8), w107=> Pw(80)(107*8-1 downto 106*8), w108=> Pw(80)(108*8-1 downto 107*8), w109=> Pw(80)(109*8-1 downto 108*8), w110=> Pw(80)(110*8-1 downto 109*8), w111=> Pw(80)(111*8-1 downto 110*8), w112=> Pw(80)(112*8-1 downto 111*8), 
w113=> Pw(80)(113*8-1 downto 112*8), w114=> Pw(80)(114*8-1 downto 113*8), w115=> Pw(80)(115*8-1 downto 114*8), w116=> Pw(80)(116*8-1 downto 115*8), w117=> Pw(80)(117*8-1 downto 116*8), w118=> Pw(80)(118*8-1 downto 117*8), w119=> Pw(80)(119*8-1 downto 118*8), w120=> Pw(80)(120*8-1 downto 119*8), 
w121=> Pw(80)(121*8-1 downto 120*8), w122=> Pw(80)(122*8-1 downto 121*8), w123=> Pw(80)(123*8-1 downto 122*8), w124=> Pw(80)(124*8-1 downto 123*8), w125=> Pw(80)(125*8-1 downto 124*8), w126=> Pw(80)(126*8-1 downto 125*8), w127=> Pw(80)(127*8-1 downto 126*8), w128=> Pw(80)(128*8-1 downto 127*8), 
           d_out   => pca_d80_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_81_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(81)(     7 downto    0),   w02 => Pw(81)( 2*8-1 downto    8),   w03 => Pw(81)( 3*8-1 downto  2*8),   w04 => Pw(81)( 4*8-1 downto  3*8),   w05 => Pw(81)( 5*8-1 downto  4*8),   w06 => Pw(81)( 6*8-1 downto  5*8),   w07 => Pw(81)( 7*8-1 downto  6*8),   w08 => Pw(81)( 8*8-1 downto  7*8),  
w09 => Pw(81)( 9*8-1 downto  8*8),   w10 => Pw(81)(10*8-1 downto  9*8),   w11 => Pw(81)(11*8-1 downto 10*8),   w12 => Pw(81)(12*8-1 downto 11*8),   w13 => Pw(81)(13*8-1 downto 12*8),   w14 => Pw(81)(14*8-1 downto 13*8),   w15 => Pw(81)(15*8-1 downto 14*8),   w16 => Pw(81)(16*8-1 downto 15*8),  
w17 => Pw(81)(17*8-1 downto 16*8),   w18 => Pw(81)(18*8-1 downto 17*8),   w19 => Pw(81)(19*8-1 downto 18*8),   w20 => Pw(81)(20*8-1 downto 19*8),   w21 => Pw(81)(21*8-1 downto 20*8),   w22 => Pw(81)(22*8-1 downto 21*8),   w23 => Pw(81)(23*8-1 downto 22*8),   w24 => Pw(81)(24*8-1 downto 23*8),  
w25 => Pw(81)(25*8-1 downto 24*8),   w26 => Pw(81)(26*8-1 downto 25*8),   w27 => Pw(81)(27*8-1 downto 26*8),   w28 => Pw(81)(28*8-1 downto 27*8),   w29 => Pw(81)(29*8-1 downto 28*8),   w30 => Pw(81)(30*8-1 downto 29*8),   w31 => Pw(81)(31*8-1 downto 30*8),   w32 => Pw(81)(32*8-1 downto 31*8),  
w33 => Pw(81)(33*8-1 downto 32*8),   w34 => Pw(81)(34*8-1 downto 33*8),   w35 => Pw(81)(35*8-1 downto 34*8),   w36 => Pw(81)(36*8-1 downto 35*8),   w37 => Pw(81)(37*8-1 downto 36*8),   w38 => Pw(81)(38*8-1 downto 37*8),   w39 => Pw(81)(39*8-1 downto 38*8),   w40 => Pw(81)(40*8-1 downto 39*8),  
w41 => Pw(81)(41*8-1 downto 40*8),   w42 => Pw(81)(42*8-1 downto 41*8),   w43 => Pw(81)(43*8-1 downto 42*8),   w44 => Pw(81)(44*8-1 downto 43*8),   w45 => Pw(81)(45*8-1 downto 44*8),   w46 => Pw(81)(46*8-1 downto 45*8),   w47 => Pw(81)(47*8-1 downto 46*8),   w48 => Pw(81)(48*8-1 downto 47*8),  
w49 => Pw(81)(49*8-1 downto 48*8),   w50 => Pw(81)(50*8-1 downto 49*8),   w51 => Pw(81)(51*8-1 downto 50*8),   w52 => Pw(81)(52*8-1 downto 51*8),   w53 => Pw(81)(53*8-1 downto 52*8),   w54 => Pw(81)(54*8-1 downto 53*8),   w55 => Pw(81)(55*8-1 downto 54*8),   w56 => Pw(81)(56*8-1 downto 55*8),  
w57 => Pw(81)(57*8-1 downto 56*8),   w58 => Pw(81)(58*8-1 downto 57*8),   w59 => Pw(81)(59*8-1 downto 58*8),   w60 => Pw(81)(60*8-1 downto 59*8),   w61 => Pw(81)(61*8-1 downto 60*8),   w62 => Pw(81)(62*8-1 downto 61*8),   w63 => Pw(81)(63*8-1 downto 62*8),   w64 => Pw(81)(64*8-1 downto 63*8), 
w65 => Pw(81)( 65*8-1 downto  64*8), w66 => Pw(81)( 66*8-1 downto  65*8), w67 => Pw(81)( 67*8-1 downto  66*8), w68 => Pw(81)( 68*8-1 downto  67*8), w69 => Pw(81)( 69*8-1 downto  68*8), w70 => Pw(81)( 70*8-1 downto  69*8), w71 => Pw(81)( 71*8-1 downto  70*8), w72 => Pw(81)( 72*8-1 downto  71*8), 
w73 => Pw(81)( 73*8-1 downto  72*8), w74 => Pw(81)( 74*8-1 downto  73*8), w75 => Pw(81)( 75*8-1 downto  74*8), w76 => Pw(81)( 76*8-1 downto  75*8), w77 => Pw(81)( 77*8-1 downto  76*8), w78 => Pw(81)( 78*8-1 downto  77*8), w79 => Pw(81)( 79*8-1 downto  78*8), w80 => Pw(81)( 80*8-1 downto  79*8), 
w81 => Pw(81)( 81*8-1 downto  80*8), w82 => Pw(81)( 82*8-1 downto  81*8), w83 => Pw(81)( 83*8-1 downto  82*8), w84 => Pw(81)( 84*8-1 downto  83*8), w85 => Pw(81)( 85*8-1 downto  84*8), w86 => Pw(81)( 86*8-1 downto  85*8), w87 => Pw(81)( 87*8-1 downto  86*8), w88 => Pw(81)( 88*8-1 downto  87*8), 
w89 => Pw(81)( 89*8-1 downto  88*8), w90 => Pw(81)( 90*8-1 downto  89*8), w91 => Pw(81)( 91*8-1 downto  90*8), w92 => Pw(81)( 92*8-1 downto  91*8), w93 => Pw(81)( 93*8-1 downto  92*8), w94 => Pw(81)( 94*8-1 downto  93*8), w95 => Pw(81)( 95*8-1 downto  94*8), w96 => Pw(81)( 96*8-1 downto  95*8), 
w97 => Pw(81)( 97*8-1 downto  96*8), w98 => Pw(81)( 98*8-1 downto  97*8), w99 => Pw(81)( 99*8-1 downto  98*8), w100=> Pw(81)(100*8-1 downto  99*8), w101=> Pw(81)(101*8-1 downto 100*8), w102=> Pw(81)(102*8-1 downto 101*8), w103=> Pw(81)(103*8-1 downto 102*8), w104=> Pw(81)(104*8-1 downto 103*8), 
w105=> Pw(81)(105*8-1 downto 104*8), w106=> Pw(81)(106*8-1 downto 105*8), w107=> Pw(81)(107*8-1 downto 106*8), w108=> Pw(81)(108*8-1 downto 107*8), w109=> Pw(81)(109*8-1 downto 108*8), w110=> Pw(81)(110*8-1 downto 109*8), w111=> Pw(81)(111*8-1 downto 110*8), w112=> Pw(81)(112*8-1 downto 111*8), 
w113=> Pw(81)(113*8-1 downto 112*8), w114=> Pw(81)(114*8-1 downto 113*8), w115=> Pw(81)(115*8-1 downto 114*8), w116=> Pw(81)(116*8-1 downto 115*8), w117=> Pw(81)(117*8-1 downto 116*8), w118=> Pw(81)(118*8-1 downto 117*8), w119=> Pw(81)(119*8-1 downto 118*8), w120=> Pw(81)(120*8-1 downto 119*8), 
w121=> Pw(81)(121*8-1 downto 120*8), w122=> Pw(81)(122*8-1 downto 121*8), w123=> Pw(81)(123*8-1 downto 122*8), w124=> Pw(81)(124*8-1 downto 123*8), w125=> Pw(81)(125*8-1 downto 124*8), w126=> Pw(81)(126*8-1 downto 125*8), w127=> Pw(81)(127*8-1 downto 126*8), w128=> Pw(81)(128*8-1 downto 127*8), 
           d_out   => pca_d81_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_82_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(82)(     7 downto    0),   w02 => Pw(82)( 2*8-1 downto    8),   w03 => Pw(82)( 3*8-1 downto  2*8),   w04 => Pw(82)( 4*8-1 downto  3*8),   w05 => Pw(82)( 5*8-1 downto  4*8),   w06 => Pw(82)( 6*8-1 downto  5*8),   w07 => Pw(82)( 7*8-1 downto  6*8),   w08 => Pw(82)( 8*8-1 downto  7*8),  
w09 => Pw(82)( 9*8-1 downto  8*8),   w10 => Pw(82)(10*8-1 downto  9*8),   w11 => Pw(82)(11*8-1 downto 10*8),   w12 => Pw(82)(12*8-1 downto 11*8),   w13 => Pw(82)(13*8-1 downto 12*8),   w14 => Pw(82)(14*8-1 downto 13*8),   w15 => Pw(82)(15*8-1 downto 14*8),   w16 => Pw(82)(16*8-1 downto 15*8),  
w17 => Pw(82)(17*8-1 downto 16*8),   w18 => Pw(82)(18*8-1 downto 17*8),   w19 => Pw(82)(19*8-1 downto 18*8),   w20 => Pw(82)(20*8-1 downto 19*8),   w21 => Pw(82)(21*8-1 downto 20*8),   w22 => Pw(82)(22*8-1 downto 21*8),   w23 => Pw(82)(23*8-1 downto 22*8),   w24 => Pw(82)(24*8-1 downto 23*8),  
w25 => Pw(82)(25*8-1 downto 24*8),   w26 => Pw(82)(26*8-1 downto 25*8),   w27 => Pw(82)(27*8-1 downto 26*8),   w28 => Pw(82)(28*8-1 downto 27*8),   w29 => Pw(82)(29*8-1 downto 28*8),   w30 => Pw(82)(30*8-1 downto 29*8),   w31 => Pw(82)(31*8-1 downto 30*8),   w32 => Pw(82)(32*8-1 downto 31*8),  
w33 => Pw(82)(33*8-1 downto 32*8),   w34 => Pw(82)(34*8-1 downto 33*8),   w35 => Pw(82)(35*8-1 downto 34*8),   w36 => Pw(82)(36*8-1 downto 35*8),   w37 => Pw(82)(37*8-1 downto 36*8),   w38 => Pw(82)(38*8-1 downto 37*8),   w39 => Pw(82)(39*8-1 downto 38*8),   w40 => Pw(82)(40*8-1 downto 39*8),  
w41 => Pw(82)(41*8-1 downto 40*8),   w42 => Pw(82)(42*8-1 downto 41*8),   w43 => Pw(82)(43*8-1 downto 42*8),   w44 => Pw(82)(44*8-1 downto 43*8),   w45 => Pw(82)(45*8-1 downto 44*8),   w46 => Pw(82)(46*8-1 downto 45*8),   w47 => Pw(82)(47*8-1 downto 46*8),   w48 => Pw(82)(48*8-1 downto 47*8),  
w49 => Pw(82)(49*8-1 downto 48*8),   w50 => Pw(82)(50*8-1 downto 49*8),   w51 => Pw(82)(51*8-1 downto 50*8),   w52 => Pw(82)(52*8-1 downto 51*8),   w53 => Pw(82)(53*8-1 downto 52*8),   w54 => Pw(82)(54*8-1 downto 53*8),   w55 => Pw(82)(55*8-1 downto 54*8),   w56 => Pw(82)(56*8-1 downto 55*8),  
w57 => Pw(82)(57*8-1 downto 56*8),   w58 => Pw(82)(58*8-1 downto 57*8),   w59 => Pw(82)(59*8-1 downto 58*8),   w60 => Pw(82)(60*8-1 downto 59*8),   w61 => Pw(82)(61*8-1 downto 60*8),   w62 => Pw(82)(62*8-1 downto 61*8),   w63 => Pw(82)(63*8-1 downto 62*8),   w64 => Pw(82)(64*8-1 downto 63*8), 
w65 => Pw(82)( 65*8-1 downto  64*8), w66 => Pw(82)( 66*8-1 downto  65*8), w67 => Pw(82)( 67*8-1 downto  66*8), w68 => Pw(82)( 68*8-1 downto  67*8), w69 => Pw(82)( 69*8-1 downto  68*8), w70 => Pw(82)( 70*8-1 downto  69*8), w71 => Pw(82)( 71*8-1 downto  70*8), w72 => Pw(82)( 72*8-1 downto  71*8), 
w73 => Pw(82)( 73*8-1 downto  72*8), w74 => Pw(82)( 74*8-1 downto  73*8), w75 => Pw(82)( 75*8-1 downto  74*8), w76 => Pw(82)( 76*8-1 downto  75*8), w77 => Pw(82)( 77*8-1 downto  76*8), w78 => Pw(82)( 78*8-1 downto  77*8), w79 => Pw(82)( 79*8-1 downto  78*8), w80 => Pw(82)( 80*8-1 downto  79*8), 
w81 => Pw(82)( 81*8-1 downto  80*8), w82 => Pw(82)( 82*8-1 downto  81*8), w83 => Pw(82)( 83*8-1 downto  82*8), w84 => Pw(82)( 84*8-1 downto  83*8), w85 => Pw(82)( 85*8-1 downto  84*8), w86 => Pw(82)( 86*8-1 downto  85*8), w87 => Pw(82)( 87*8-1 downto  86*8), w88 => Pw(82)( 88*8-1 downto  87*8), 
w89 => Pw(82)( 89*8-1 downto  88*8), w90 => Pw(82)( 90*8-1 downto  89*8), w91 => Pw(82)( 91*8-1 downto  90*8), w92 => Pw(82)( 92*8-1 downto  91*8), w93 => Pw(82)( 93*8-1 downto  92*8), w94 => Pw(82)( 94*8-1 downto  93*8), w95 => Pw(82)( 95*8-1 downto  94*8), w96 => Pw(82)( 96*8-1 downto  95*8), 
w97 => Pw(82)( 97*8-1 downto  96*8), w98 => Pw(82)( 98*8-1 downto  97*8), w99 => Pw(82)( 99*8-1 downto  98*8), w100=> Pw(82)(100*8-1 downto  99*8), w101=> Pw(82)(101*8-1 downto 100*8), w102=> Pw(82)(102*8-1 downto 101*8), w103=> Pw(82)(103*8-1 downto 102*8), w104=> Pw(82)(104*8-1 downto 103*8), 
w105=> Pw(82)(105*8-1 downto 104*8), w106=> Pw(82)(106*8-1 downto 105*8), w107=> Pw(82)(107*8-1 downto 106*8), w108=> Pw(82)(108*8-1 downto 107*8), w109=> Pw(82)(109*8-1 downto 108*8), w110=> Pw(82)(110*8-1 downto 109*8), w111=> Pw(82)(111*8-1 downto 110*8), w112=> Pw(82)(112*8-1 downto 111*8), 
w113=> Pw(82)(113*8-1 downto 112*8), w114=> Pw(82)(114*8-1 downto 113*8), w115=> Pw(82)(115*8-1 downto 114*8), w116=> Pw(82)(116*8-1 downto 115*8), w117=> Pw(82)(117*8-1 downto 116*8), w118=> Pw(82)(118*8-1 downto 117*8), w119=> Pw(82)(119*8-1 downto 118*8), w120=> Pw(82)(120*8-1 downto 119*8), 
w121=> Pw(82)(121*8-1 downto 120*8), w122=> Pw(82)(122*8-1 downto 121*8), w123=> Pw(82)(123*8-1 downto 122*8), w124=> Pw(82)(124*8-1 downto 123*8), w125=> Pw(82)(125*8-1 downto 124*8), w126=> Pw(82)(126*8-1 downto 125*8), w127=> Pw(82)(127*8-1 downto 126*8), w128=> Pw(82)(128*8-1 downto 127*8), 
           d_out   => pca_d82_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_83_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(83)(     7 downto    0),   w02 => Pw(83)( 2*8-1 downto    8),   w03 => Pw(83)( 3*8-1 downto  2*8),   w04 => Pw(83)( 4*8-1 downto  3*8),   w05 => Pw(83)( 5*8-1 downto  4*8),   w06 => Pw(83)( 6*8-1 downto  5*8),   w07 => Pw(83)( 7*8-1 downto  6*8),   w08 => Pw(83)( 8*8-1 downto  7*8),  
w09 => Pw(83)( 9*8-1 downto  8*8),   w10 => Pw(83)(10*8-1 downto  9*8),   w11 => Pw(83)(11*8-1 downto 10*8),   w12 => Pw(83)(12*8-1 downto 11*8),   w13 => Pw(83)(13*8-1 downto 12*8),   w14 => Pw(83)(14*8-1 downto 13*8),   w15 => Pw(83)(15*8-1 downto 14*8),   w16 => Pw(83)(16*8-1 downto 15*8),  
w17 => Pw(83)(17*8-1 downto 16*8),   w18 => Pw(83)(18*8-1 downto 17*8),   w19 => Pw(83)(19*8-1 downto 18*8),   w20 => Pw(83)(20*8-1 downto 19*8),   w21 => Pw(83)(21*8-1 downto 20*8),   w22 => Pw(83)(22*8-1 downto 21*8),   w23 => Pw(83)(23*8-1 downto 22*8),   w24 => Pw(83)(24*8-1 downto 23*8),  
w25 => Pw(83)(25*8-1 downto 24*8),   w26 => Pw(83)(26*8-1 downto 25*8),   w27 => Pw(83)(27*8-1 downto 26*8),   w28 => Pw(83)(28*8-1 downto 27*8),   w29 => Pw(83)(29*8-1 downto 28*8),   w30 => Pw(83)(30*8-1 downto 29*8),   w31 => Pw(83)(31*8-1 downto 30*8),   w32 => Pw(83)(32*8-1 downto 31*8),  
w33 => Pw(83)(33*8-1 downto 32*8),   w34 => Pw(83)(34*8-1 downto 33*8),   w35 => Pw(83)(35*8-1 downto 34*8),   w36 => Pw(83)(36*8-1 downto 35*8),   w37 => Pw(83)(37*8-1 downto 36*8),   w38 => Pw(83)(38*8-1 downto 37*8),   w39 => Pw(83)(39*8-1 downto 38*8),   w40 => Pw(83)(40*8-1 downto 39*8),  
w41 => Pw(83)(41*8-1 downto 40*8),   w42 => Pw(83)(42*8-1 downto 41*8),   w43 => Pw(83)(43*8-1 downto 42*8),   w44 => Pw(83)(44*8-1 downto 43*8),   w45 => Pw(83)(45*8-1 downto 44*8),   w46 => Pw(83)(46*8-1 downto 45*8),   w47 => Pw(83)(47*8-1 downto 46*8),   w48 => Pw(83)(48*8-1 downto 47*8),  
w49 => Pw(83)(49*8-1 downto 48*8),   w50 => Pw(83)(50*8-1 downto 49*8),   w51 => Pw(83)(51*8-1 downto 50*8),   w52 => Pw(83)(52*8-1 downto 51*8),   w53 => Pw(83)(53*8-1 downto 52*8),   w54 => Pw(83)(54*8-1 downto 53*8),   w55 => Pw(83)(55*8-1 downto 54*8),   w56 => Pw(83)(56*8-1 downto 55*8),  
w57 => Pw(83)(57*8-1 downto 56*8),   w58 => Pw(83)(58*8-1 downto 57*8),   w59 => Pw(83)(59*8-1 downto 58*8),   w60 => Pw(83)(60*8-1 downto 59*8),   w61 => Pw(83)(61*8-1 downto 60*8),   w62 => Pw(83)(62*8-1 downto 61*8),   w63 => Pw(83)(63*8-1 downto 62*8),   w64 => Pw(83)(64*8-1 downto 63*8), 
w65 => Pw(83)( 65*8-1 downto  64*8), w66 => Pw(83)( 66*8-1 downto  65*8), w67 => Pw(83)( 67*8-1 downto  66*8), w68 => Pw(83)( 68*8-1 downto  67*8), w69 => Pw(83)( 69*8-1 downto  68*8), w70 => Pw(83)( 70*8-1 downto  69*8), w71 => Pw(83)( 71*8-1 downto  70*8), w72 => Pw(83)( 72*8-1 downto  71*8), 
w73 => Pw(83)( 73*8-1 downto  72*8), w74 => Pw(83)( 74*8-1 downto  73*8), w75 => Pw(83)( 75*8-1 downto  74*8), w76 => Pw(83)( 76*8-1 downto  75*8), w77 => Pw(83)( 77*8-1 downto  76*8), w78 => Pw(83)( 78*8-1 downto  77*8), w79 => Pw(83)( 79*8-1 downto  78*8), w80 => Pw(83)( 80*8-1 downto  79*8), 
w81 => Pw(83)( 81*8-1 downto  80*8), w82 => Pw(83)( 82*8-1 downto  81*8), w83 => Pw(83)( 83*8-1 downto  82*8), w84 => Pw(83)( 84*8-1 downto  83*8), w85 => Pw(83)( 85*8-1 downto  84*8), w86 => Pw(83)( 86*8-1 downto  85*8), w87 => Pw(83)( 87*8-1 downto  86*8), w88 => Pw(83)( 88*8-1 downto  87*8), 
w89 => Pw(83)( 89*8-1 downto  88*8), w90 => Pw(83)( 90*8-1 downto  89*8), w91 => Pw(83)( 91*8-1 downto  90*8), w92 => Pw(83)( 92*8-1 downto  91*8), w93 => Pw(83)( 93*8-1 downto  92*8), w94 => Pw(83)( 94*8-1 downto  93*8), w95 => Pw(83)( 95*8-1 downto  94*8), w96 => Pw(83)( 96*8-1 downto  95*8), 
w97 => Pw(83)( 97*8-1 downto  96*8), w98 => Pw(83)( 98*8-1 downto  97*8), w99 => Pw(83)( 99*8-1 downto  98*8), w100=> Pw(83)(100*8-1 downto  99*8), w101=> Pw(83)(101*8-1 downto 100*8), w102=> Pw(83)(102*8-1 downto 101*8), w103=> Pw(83)(103*8-1 downto 102*8), w104=> Pw(83)(104*8-1 downto 103*8), 
w105=> Pw(83)(105*8-1 downto 104*8), w106=> Pw(83)(106*8-1 downto 105*8), w107=> Pw(83)(107*8-1 downto 106*8), w108=> Pw(83)(108*8-1 downto 107*8), w109=> Pw(83)(109*8-1 downto 108*8), w110=> Pw(83)(110*8-1 downto 109*8), w111=> Pw(83)(111*8-1 downto 110*8), w112=> Pw(83)(112*8-1 downto 111*8), 
w113=> Pw(83)(113*8-1 downto 112*8), w114=> Pw(83)(114*8-1 downto 113*8), w115=> Pw(83)(115*8-1 downto 114*8), w116=> Pw(83)(116*8-1 downto 115*8), w117=> Pw(83)(117*8-1 downto 116*8), w118=> Pw(83)(118*8-1 downto 117*8), w119=> Pw(83)(119*8-1 downto 118*8), w120=> Pw(83)(120*8-1 downto 119*8), 
w121=> Pw(83)(121*8-1 downto 120*8), w122=> Pw(83)(122*8-1 downto 121*8), w123=> Pw(83)(123*8-1 downto 122*8), w124=> Pw(83)(124*8-1 downto 123*8), w125=> Pw(83)(125*8-1 downto 124*8), w126=> Pw(83)(126*8-1 downto 125*8), w127=> Pw(83)(127*8-1 downto 126*8), w128=> Pw(83)(128*8-1 downto 127*8), 
           d_out   => pca_d83_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_84_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(84)(     7 downto    0),   w02 => Pw(84)( 2*8-1 downto    8),   w03 => Pw(84)( 3*8-1 downto  2*8),   w04 => Pw(84)( 4*8-1 downto  3*8),   w05 => Pw(84)( 5*8-1 downto  4*8),   w06 => Pw(84)( 6*8-1 downto  5*8),   w07 => Pw(84)( 7*8-1 downto  6*8),   w08 => Pw(84)( 8*8-1 downto  7*8),  
w09 => Pw(84)( 9*8-1 downto  8*8),   w10 => Pw(84)(10*8-1 downto  9*8),   w11 => Pw(84)(11*8-1 downto 10*8),   w12 => Pw(84)(12*8-1 downto 11*8),   w13 => Pw(84)(13*8-1 downto 12*8),   w14 => Pw(84)(14*8-1 downto 13*8),   w15 => Pw(84)(15*8-1 downto 14*8),   w16 => Pw(84)(16*8-1 downto 15*8),  
w17 => Pw(84)(17*8-1 downto 16*8),   w18 => Pw(84)(18*8-1 downto 17*8),   w19 => Pw(84)(19*8-1 downto 18*8),   w20 => Pw(84)(20*8-1 downto 19*8),   w21 => Pw(84)(21*8-1 downto 20*8),   w22 => Pw(84)(22*8-1 downto 21*8),   w23 => Pw(84)(23*8-1 downto 22*8),   w24 => Pw(84)(24*8-1 downto 23*8),  
w25 => Pw(84)(25*8-1 downto 24*8),   w26 => Pw(84)(26*8-1 downto 25*8),   w27 => Pw(84)(27*8-1 downto 26*8),   w28 => Pw(84)(28*8-1 downto 27*8),   w29 => Pw(84)(29*8-1 downto 28*8),   w30 => Pw(84)(30*8-1 downto 29*8),   w31 => Pw(84)(31*8-1 downto 30*8),   w32 => Pw(84)(32*8-1 downto 31*8),  
w33 => Pw(84)(33*8-1 downto 32*8),   w34 => Pw(84)(34*8-1 downto 33*8),   w35 => Pw(84)(35*8-1 downto 34*8),   w36 => Pw(84)(36*8-1 downto 35*8),   w37 => Pw(84)(37*8-1 downto 36*8),   w38 => Pw(84)(38*8-1 downto 37*8),   w39 => Pw(84)(39*8-1 downto 38*8),   w40 => Pw(84)(40*8-1 downto 39*8),  
w41 => Pw(84)(41*8-1 downto 40*8),   w42 => Pw(84)(42*8-1 downto 41*8),   w43 => Pw(84)(43*8-1 downto 42*8),   w44 => Pw(84)(44*8-1 downto 43*8),   w45 => Pw(84)(45*8-1 downto 44*8),   w46 => Pw(84)(46*8-1 downto 45*8),   w47 => Pw(84)(47*8-1 downto 46*8),   w48 => Pw(84)(48*8-1 downto 47*8),  
w49 => Pw(84)(49*8-1 downto 48*8),   w50 => Pw(84)(50*8-1 downto 49*8),   w51 => Pw(84)(51*8-1 downto 50*8),   w52 => Pw(84)(52*8-1 downto 51*8),   w53 => Pw(84)(53*8-1 downto 52*8),   w54 => Pw(84)(54*8-1 downto 53*8),   w55 => Pw(84)(55*8-1 downto 54*8),   w56 => Pw(84)(56*8-1 downto 55*8),  
w57 => Pw(84)(57*8-1 downto 56*8),   w58 => Pw(84)(58*8-1 downto 57*8),   w59 => Pw(84)(59*8-1 downto 58*8),   w60 => Pw(84)(60*8-1 downto 59*8),   w61 => Pw(84)(61*8-1 downto 60*8),   w62 => Pw(84)(62*8-1 downto 61*8),   w63 => Pw(84)(63*8-1 downto 62*8),   w64 => Pw(84)(64*8-1 downto 63*8), 
w65 => Pw(84)( 65*8-1 downto  64*8), w66 => Pw(84)( 66*8-1 downto  65*8), w67 => Pw(84)( 67*8-1 downto  66*8), w68 => Pw(84)( 68*8-1 downto  67*8), w69 => Pw(84)( 69*8-1 downto  68*8), w70 => Pw(84)( 70*8-1 downto  69*8), w71 => Pw(84)( 71*8-1 downto  70*8), w72 => Pw(84)( 72*8-1 downto  71*8), 
w73 => Pw(84)( 73*8-1 downto  72*8), w74 => Pw(84)( 74*8-1 downto  73*8), w75 => Pw(84)( 75*8-1 downto  74*8), w76 => Pw(84)( 76*8-1 downto  75*8), w77 => Pw(84)( 77*8-1 downto  76*8), w78 => Pw(84)( 78*8-1 downto  77*8), w79 => Pw(84)( 79*8-1 downto  78*8), w80 => Pw(84)( 80*8-1 downto  79*8), 
w81 => Pw(84)( 81*8-1 downto  80*8), w82 => Pw(84)( 82*8-1 downto  81*8), w83 => Pw(84)( 83*8-1 downto  82*8), w84 => Pw(84)( 84*8-1 downto  83*8), w85 => Pw(84)( 85*8-1 downto  84*8), w86 => Pw(84)( 86*8-1 downto  85*8), w87 => Pw(84)( 87*8-1 downto  86*8), w88 => Pw(84)( 88*8-1 downto  87*8), 
w89 => Pw(84)( 89*8-1 downto  88*8), w90 => Pw(84)( 90*8-1 downto  89*8), w91 => Pw(84)( 91*8-1 downto  90*8), w92 => Pw(84)( 92*8-1 downto  91*8), w93 => Pw(84)( 93*8-1 downto  92*8), w94 => Pw(84)( 94*8-1 downto  93*8), w95 => Pw(84)( 95*8-1 downto  94*8), w96 => Pw(84)( 96*8-1 downto  95*8), 
w97 => Pw(84)( 97*8-1 downto  96*8), w98 => Pw(84)( 98*8-1 downto  97*8), w99 => Pw(84)( 99*8-1 downto  98*8), w100=> Pw(84)(100*8-1 downto  99*8), w101=> Pw(84)(101*8-1 downto 100*8), w102=> Pw(84)(102*8-1 downto 101*8), w103=> Pw(84)(103*8-1 downto 102*8), w104=> Pw(84)(104*8-1 downto 103*8), 
w105=> Pw(84)(105*8-1 downto 104*8), w106=> Pw(84)(106*8-1 downto 105*8), w107=> Pw(84)(107*8-1 downto 106*8), w108=> Pw(84)(108*8-1 downto 107*8), w109=> Pw(84)(109*8-1 downto 108*8), w110=> Pw(84)(110*8-1 downto 109*8), w111=> Pw(84)(111*8-1 downto 110*8), w112=> Pw(84)(112*8-1 downto 111*8), 
w113=> Pw(84)(113*8-1 downto 112*8), w114=> Pw(84)(114*8-1 downto 113*8), w115=> Pw(84)(115*8-1 downto 114*8), w116=> Pw(84)(116*8-1 downto 115*8), w117=> Pw(84)(117*8-1 downto 116*8), w118=> Pw(84)(118*8-1 downto 117*8), w119=> Pw(84)(119*8-1 downto 118*8), w120=> Pw(84)(120*8-1 downto 119*8), 
w121=> Pw(84)(121*8-1 downto 120*8), w122=> Pw(84)(122*8-1 downto 121*8), w123=> Pw(84)(123*8-1 downto 122*8), w124=> Pw(84)(124*8-1 downto 123*8), w125=> Pw(84)(125*8-1 downto 124*8), w126=> Pw(84)(126*8-1 downto 125*8), w127=> Pw(84)(127*8-1 downto 126*8), w128=> Pw(84)(128*8-1 downto 127*8), 
           d_out   => pca_d84_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_85_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(85)(     7 downto    0),   w02 => Pw(85)( 2*8-1 downto    8),   w03 => Pw(85)( 3*8-1 downto  2*8),   w04 => Pw(85)( 4*8-1 downto  3*8),   w05 => Pw(85)( 5*8-1 downto  4*8),   w06 => Pw(85)( 6*8-1 downto  5*8),   w07 => Pw(85)( 7*8-1 downto  6*8),   w08 => Pw(85)( 8*8-1 downto  7*8),  
w09 => Pw(85)( 9*8-1 downto  8*8),   w10 => Pw(85)(10*8-1 downto  9*8),   w11 => Pw(85)(11*8-1 downto 10*8),   w12 => Pw(85)(12*8-1 downto 11*8),   w13 => Pw(85)(13*8-1 downto 12*8),   w14 => Pw(85)(14*8-1 downto 13*8),   w15 => Pw(85)(15*8-1 downto 14*8),   w16 => Pw(85)(16*8-1 downto 15*8),  
w17 => Pw(85)(17*8-1 downto 16*8),   w18 => Pw(85)(18*8-1 downto 17*8),   w19 => Pw(85)(19*8-1 downto 18*8),   w20 => Pw(85)(20*8-1 downto 19*8),   w21 => Pw(85)(21*8-1 downto 20*8),   w22 => Pw(85)(22*8-1 downto 21*8),   w23 => Pw(85)(23*8-1 downto 22*8),   w24 => Pw(85)(24*8-1 downto 23*8),  
w25 => Pw(85)(25*8-1 downto 24*8),   w26 => Pw(85)(26*8-1 downto 25*8),   w27 => Pw(85)(27*8-1 downto 26*8),   w28 => Pw(85)(28*8-1 downto 27*8),   w29 => Pw(85)(29*8-1 downto 28*8),   w30 => Pw(85)(30*8-1 downto 29*8),   w31 => Pw(85)(31*8-1 downto 30*8),   w32 => Pw(85)(32*8-1 downto 31*8),  
w33 => Pw(85)(33*8-1 downto 32*8),   w34 => Pw(85)(34*8-1 downto 33*8),   w35 => Pw(85)(35*8-1 downto 34*8),   w36 => Pw(85)(36*8-1 downto 35*8),   w37 => Pw(85)(37*8-1 downto 36*8),   w38 => Pw(85)(38*8-1 downto 37*8),   w39 => Pw(85)(39*8-1 downto 38*8),   w40 => Pw(85)(40*8-1 downto 39*8),  
w41 => Pw(85)(41*8-1 downto 40*8),   w42 => Pw(85)(42*8-1 downto 41*8),   w43 => Pw(85)(43*8-1 downto 42*8),   w44 => Pw(85)(44*8-1 downto 43*8),   w45 => Pw(85)(45*8-1 downto 44*8),   w46 => Pw(85)(46*8-1 downto 45*8),   w47 => Pw(85)(47*8-1 downto 46*8),   w48 => Pw(85)(48*8-1 downto 47*8),  
w49 => Pw(85)(49*8-1 downto 48*8),   w50 => Pw(85)(50*8-1 downto 49*8),   w51 => Pw(85)(51*8-1 downto 50*8),   w52 => Pw(85)(52*8-1 downto 51*8),   w53 => Pw(85)(53*8-1 downto 52*8),   w54 => Pw(85)(54*8-1 downto 53*8),   w55 => Pw(85)(55*8-1 downto 54*8),   w56 => Pw(85)(56*8-1 downto 55*8),  
w57 => Pw(85)(57*8-1 downto 56*8),   w58 => Pw(85)(58*8-1 downto 57*8),   w59 => Pw(85)(59*8-1 downto 58*8),   w60 => Pw(85)(60*8-1 downto 59*8),   w61 => Pw(85)(61*8-1 downto 60*8),   w62 => Pw(85)(62*8-1 downto 61*8),   w63 => Pw(85)(63*8-1 downto 62*8),   w64 => Pw(85)(64*8-1 downto 63*8), 
w65 => Pw(85)( 65*8-1 downto  64*8), w66 => Pw(85)( 66*8-1 downto  65*8), w67 => Pw(85)( 67*8-1 downto  66*8), w68 => Pw(85)( 68*8-1 downto  67*8), w69 => Pw(85)( 69*8-1 downto  68*8), w70 => Pw(85)( 70*8-1 downto  69*8), w71 => Pw(85)( 71*8-1 downto  70*8), w72 => Pw(85)( 72*8-1 downto  71*8), 
w73 => Pw(85)( 73*8-1 downto  72*8), w74 => Pw(85)( 74*8-1 downto  73*8), w75 => Pw(85)( 75*8-1 downto  74*8), w76 => Pw(85)( 76*8-1 downto  75*8), w77 => Pw(85)( 77*8-1 downto  76*8), w78 => Pw(85)( 78*8-1 downto  77*8), w79 => Pw(85)( 79*8-1 downto  78*8), w80 => Pw(85)( 80*8-1 downto  79*8), 
w81 => Pw(85)( 81*8-1 downto  80*8), w82 => Pw(85)( 82*8-1 downto  81*8), w83 => Pw(85)( 83*8-1 downto  82*8), w84 => Pw(85)( 84*8-1 downto  83*8), w85 => Pw(85)( 85*8-1 downto  84*8), w86 => Pw(85)( 86*8-1 downto  85*8), w87 => Pw(85)( 87*8-1 downto  86*8), w88 => Pw(85)( 88*8-1 downto  87*8), 
w89 => Pw(85)( 89*8-1 downto  88*8), w90 => Pw(85)( 90*8-1 downto  89*8), w91 => Pw(85)( 91*8-1 downto  90*8), w92 => Pw(85)( 92*8-1 downto  91*8), w93 => Pw(85)( 93*8-1 downto  92*8), w94 => Pw(85)( 94*8-1 downto  93*8), w95 => Pw(85)( 95*8-1 downto  94*8), w96 => Pw(85)( 96*8-1 downto  95*8), 
w97 => Pw(85)( 97*8-1 downto  96*8), w98 => Pw(85)( 98*8-1 downto  97*8), w99 => Pw(85)( 99*8-1 downto  98*8), w100=> Pw(85)(100*8-1 downto  99*8), w101=> Pw(85)(101*8-1 downto 100*8), w102=> Pw(85)(102*8-1 downto 101*8), w103=> Pw(85)(103*8-1 downto 102*8), w104=> Pw(85)(104*8-1 downto 103*8), 
w105=> Pw(85)(105*8-1 downto 104*8), w106=> Pw(85)(106*8-1 downto 105*8), w107=> Pw(85)(107*8-1 downto 106*8), w108=> Pw(85)(108*8-1 downto 107*8), w109=> Pw(85)(109*8-1 downto 108*8), w110=> Pw(85)(110*8-1 downto 109*8), w111=> Pw(85)(111*8-1 downto 110*8), w112=> Pw(85)(112*8-1 downto 111*8), 
w113=> Pw(85)(113*8-1 downto 112*8), w114=> Pw(85)(114*8-1 downto 113*8), w115=> Pw(85)(115*8-1 downto 114*8), w116=> Pw(85)(116*8-1 downto 115*8), w117=> Pw(85)(117*8-1 downto 116*8), w118=> Pw(85)(118*8-1 downto 117*8), w119=> Pw(85)(119*8-1 downto 118*8), w120=> Pw(85)(120*8-1 downto 119*8), 
w121=> Pw(85)(121*8-1 downto 120*8), w122=> Pw(85)(122*8-1 downto 121*8), w123=> Pw(85)(123*8-1 downto 122*8), w124=> Pw(85)(124*8-1 downto 123*8), w125=> Pw(85)(125*8-1 downto 124*8), w126=> Pw(85)(126*8-1 downto 125*8), w127=> Pw(85)(127*8-1 downto 126*8), w128=> Pw(85)(128*8-1 downto 127*8), 
           d_out   => pca_d85_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_86_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(86)(     7 downto    0),   w02 => Pw(86)( 2*8-1 downto    8),   w03 => Pw(86)( 3*8-1 downto  2*8),   w04 => Pw(86)( 4*8-1 downto  3*8),   w05 => Pw(86)( 5*8-1 downto  4*8),   w06 => Pw(86)( 6*8-1 downto  5*8),   w07 => Pw(86)( 7*8-1 downto  6*8),   w08 => Pw(86)( 8*8-1 downto  7*8),  
w09 => Pw(86)( 9*8-1 downto  8*8),   w10 => Pw(86)(10*8-1 downto  9*8),   w11 => Pw(86)(11*8-1 downto 10*8),   w12 => Pw(86)(12*8-1 downto 11*8),   w13 => Pw(86)(13*8-1 downto 12*8),   w14 => Pw(86)(14*8-1 downto 13*8),   w15 => Pw(86)(15*8-1 downto 14*8),   w16 => Pw(86)(16*8-1 downto 15*8),  
w17 => Pw(86)(17*8-1 downto 16*8),   w18 => Pw(86)(18*8-1 downto 17*8),   w19 => Pw(86)(19*8-1 downto 18*8),   w20 => Pw(86)(20*8-1 downto 19*8),   w21 => Pw(86)(21*8-1 downto 20*8),   w22 => Pw(86)(22*8-1 downto 21*8),   w23 => Pw(86)(23*8-1 downto 22*8),   w24 => Pw(86)(24*8-1 downto 23*8),  
w25 => Pw(86)(25*8-1 downto 24*8),   w26 => Pw(86)(26*8-1 downto 25*8),   w27 => Pw(86)(27*8-1 downto 26*8),   w28 => Pw(86)(28*8-1 downto 27*8),   w29 => Pw(86)(29*8-1 downto 28*8),   w30 => Pw(86)(30*8-1 downto 29*8),   w31 => Pw(86)(31*8-1 downto 30*8),   w32 => Pw(86)(32*8-1 downto 31*8),  
w33 => Pw(86)(33*8-1 downto 32*8),   w34 => Pw(86)(34*8-1 downto 33*8),   w35 => Pw(86)(35*8-1 downto 34*8),   w36 => Pw(86)(36*8-1 downto 35*8),   w37 => Pw(86)(37*8-1 downto 36*8),   w38 => Pw(86)(38*8-1 downto 37*8),   w39 => Pw(86)(39*8-1 downto 38*8),   w40 => Pw(86)(40*8-1 downto 39*8),  
w41 => Pw(86)(41*8-1 downto 40*8),   w42 => Pw(86)(42*8-1 downto 41*8),   w43 => Pw(86)(43*8-1 downto 42*8),   w44 => Pw(86)(44*8-1 downto 43*8),   w45 => Pw(86)(45*8-1 downto 44*8),   w46 => Pw(86)(46*8-1 downto 45*8),   w47 => Pw(86)(47*8-1 downto 46*8),   w48 => Pw(86)(48*8-1 downto 47*8),  
w49 => Pw(86)(49*8-1 downto 48*8),   w50 => Pw(86)(50*8-1 downto 49*8),   w51 => Pw(86)(51*8-1 downto 50*8),   w52 => Pw(86)(52*8-1 downto 51*8),   w53 => Pw(86)(53*8-1 downto 52*8),   w54 => Pw(86)(54*8-1 downto 53*8),   w55 => Pw(86)(55*8-1 downto 54*8),   w56 => Pw(86)(56*8-1 downto 55*8),  
w57 => Pw(86)(57*8-1 downto 56*8),   w58 => Pw(86)(58*8-1 downto 57*8),   w59 => Pw(86)(59*8-1 downto 58*8),   w60 => Pw(86)(60*8-1 downto 59*8),   w61 => Pw(86)(61*8-1 downto 60*8),   w62 => Pw(86)(62*8-1 downto 61*8),   w63 => Pw(86)(63*8-1 downto 62*8),   w64 => Pw(86)(64*8-1 downto 63*8), 
w65 => Pw(86)( 65*8-1 downto  64*8), w66 => Pw(86)( 66*8-1 downto  65*8), w67 => Pw(86)( 67*8-1 downto  66*8), w68 => Pw(86)( 68*8-1 downto  67*8), w69 => Pw(86)( 69*8-1 downto  68*8), w70 => Pw(86)( 70*8-1 downto  69*8), w71 => Pw(86)( 71*8-1 downto  70*8), w72 => Pw(86)( 72*8-1 downto  71*8), 
w73 => Pw(86)( 73*8-1 downto  72*8), w74 => Pw(86)( 74*8-1 downto  73*8), w75 => Pw(86)( 75*8-1 downto  74*8), w76 => Pw(86)( 76*8-1 downto  75*8), w77 => Pw(86)( 77*8-1 downto  76*8), w78 => Pw(86)( 78*8-1 downto  77*8), w79 => Pw(86)( 79*8-1 downto  78*8), w80 => Pw(86)( 80*8-1 downto  79*8), 
w81 => Pw(86)( 81*8-1 downto  80*8), w82 => Pw(86)( 82*8-1 downto  81*8), w83 => Pw(86)( 83*8-1 downto  82*8), w84 => Pw(86)( 84*8-1 downto  83*8), w85 => Pw(86)( 85*8-1 downto  84*8), w86 => Pw(86)( 86*8-1 downto  85*8), w87 => Pw(86)( 87*8-1 downto  86*8), w88 => Pw(86)( 88*8-1 downto  87*8), 
w89 => Pw(86)( 89*8-1 downto  88*8), w90 => Pw(86)( 90*8-1 downto  89*8), w91 => Pw(86)( 91*8-1 downto  90*8), w92 => Pw(86)( 92*8-1 downto  91*8), w93 => Pw(86)( 93*8-1 downto  92*8), w94 => Pw(86)( 94*8-1 downto  93*8), w95 => Pw(86)( 95*8-1 downto  94*8), w96 => Pw(86)( 96*8-1 downto  95*8), 
w97 => Pw(86)( 97*8-1 downto  96*8), w98 => Pw(86)( 98*8-1 downto  97*8), w99 => Pw(86)( 99*8-1 downto  98*8), w100=> Pw(86)(100*8-1 downto  99*8), w101=> Pw(86)(101*8-1 downto 100*8), w102=> Pw(86)(102*8-1 downto 101*8), w103=> Pw(86)(103*8-1 downto 102*8), w104=> Pw(86)(104*8-1 downto 103*8), 
w105=> Pw(86)(105*8-1 downto 104*8), w106=> Pw(86)(106*8-1 downto 105*8), w107=> Pw(86)(107*8-1 downto 106*8), w108=> Pw(86)(108*8-1 downto 107*8), w109=> Pw(86)(109*8-1 downto 108*8), w110=> Pw(86)(110*8-1 downto 109*8), w111=> Pw(86)(111*8-1 downto 110*8), w112=> Pw(86)(112*8-1 downto 111*8), 
w113=> Pw(86)(113*8-1 downto 112*8), w114=> Pw(86)(114*8-1 downto 113*8), w115=> Pw(86)(115*8-1 downto 114*8), w116=> Pw(86)(116*8-1 downto 115*8), w117=> Pw(86)(117*8-1 downto 116*8), w118=> Pw(86)(118*8-1 downto 117*8), w119=> Pw(86)(119*8-1 downto 118*8), w120=> Pw(86)(120*8-1 downto 119*8), 
w121=> Pw(86)(121*8-1 downto 120*8), w122=> Pw(86)(122*8-1 downto 121*8), w123=> Pw(86)(123*8-1 downto 122*8), w124=> Pw(86)(124*8-1 downto 123*8), w125=> Pw(86)(125*8-1 downto 124*8), w126=> Pw(86)(126*8-1 downto 125*8), w127=> Pw(86)(127*8-1 downto 126*8), w128=> Pw(86)(128*8-1 downto 127*8), 
           d_out   => pca_d86_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_87_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(87)(     7 downto    0),   w02 => Pw(87)( 2*8-1 downto    8),   w03 => Pw(87)( 3*8-1 downto  2*8),   w04 => Pw(87)( 4*8-1 downto  3*8),   w05 => Pw(87)( 5*8-1 downto  4*8),   w06 => Pw(87)( 6*8-1 downto  5*8),   w07 => Pw(87)( 7*8-1 downto  6*8),   w08 => Pw(87)( 8*8-1 downto  7*8),  
w09 => Pw(87)( 9*8-1 downto  8*8),   w10 => Pw(87)(10*8-1 downto  9*8),   w11 => Pw(87)(11*8-1 downto 10*8),   w12 => Pw(87)(12*8-1 downto 11*8),   w13 => Pw(87)(13*8-1 downto 12*8),   w14 => Pw(87)(14*8-1 downto 13*8),   w15 => Pw(87)(15*8-1 downto 14*8),   w16 => Pw(87)(16*8-1 downto 15*8),  
w17 => Pw(87)(17*8-1 downto 16*8),   w18 => Pw(87)(18*8-1 downto 17*8),   w19 => Pw(87)(19*8-1 downto 18*8),   w20 => Pw(87)(20*8-1 downto 19*8),   w21 => Pw(87)(21*8-1 downto 20*8),   w22 => Pw(87)(22*8-1 downto 21*8),   w23 => Pw(87)(23*8-1 downto 22*8),   w24 => Pw(87)(24*8-1 downto 23*8),  
w25 => Pw(87)(25*8-1 downto 24*8),   w26 => Pw(87)(26*8-1 downto 25*8),   w27 => Pw(87)(27*8-1 downto 26*8),   w28 => Pw(87)(28*8-1 downto 27*8),   w29 => Pw(87)(29*8-1 downto 28*8),   w30 => Pw(87)(30*8-1 downto 29*8),   w31 => Pw(87)(31*8-1 downto 30*8),   w32 => Pw(87)(32*8-1 downto 31*8),  
w33 => Pw(87)(33*8-1 downto 32*8),   w34 => Pw(87)(34*8-1 downto 33*8),   w35 => Pw(87)(35*8-1 downto 34*8),   w36 => Pw(87)(36*8-1 downto 35*8),   w37 => Pw(87)(37*8-1 downto 36*8),   w38 => Pw(87)(38*8-1 downto 37*8),   w39 => Pw(87)(39*8-1 downto 38*8),   w40 => Pw(87)(40*8-1 downto 39*8),  
w41 => Pw(87)(41*8-1 downto 40*8),   w42 => Pw(87)(42*8-1 downto 41*8),   w43 => Pw(87)(43*8-1 downto 42*8),   w44 => Pw(87)(44*8-1 downto 43*8),   w45 => Pw(87)(45*8-1 downto 44*8),   w46 => Pw(87)(46*8-1 downto 45*8),   w47 => Pw(87)(47*8-1 downto 46*8),   w48 => Pw(87)(48*8-1 downto 47*8),  
w49 => Pw(87)(49*8-1 downto 48*8),   w50 => Pw(87)(50*8-1 downto 49*8),   w51 => Pw(87)(51*8-1 downto 50*8),   w52 => Pw(87)(52*8-1 downto 51*8),   w53 => Pw(87)(53*8-1 downto 52*8),   w54 => Pw(87)(54*8-1 downto 53*8),   w55 => Pw(87)(55*8-1 downto 54*8),   w56 => Pw(87)(56*8-1 downto 55*8),  
w57 => Pw(87)(57*8-1 downto 56*8),   w58 => Pw(87)(58*8-1 downto 57*8),   w59 => Pw(87)(59*8-1 downto 58*8),   w60 => Pw(87)(60*8-1 downto 59*8),   w61 => Pw(87)(61*8-1 downto 60*8),   w62 => Pw(87)(62*8-1 downto 61*8),   w63 => Pw(87)(63*8-1 downto 62*8),   w64 => Pw(87)(64*8-1 downto 63*8), 
w65 => Pw(87)( 65*8-1 downto  64*8), w66 => Pw(87)( 66*8-1 downto  65*8), w67 => Pw(87)( 67*8-1 downto  66*8), w68 => Pw(87)( 68*8-1 downto  67*8), w69 => Pw(87)( 69*8-1 downto  68*8), w70 => Pw(87)( 70*8-1 downto  69*8), w71 => Pw(87)( 71*8-1 downto  70*8), w72 => Pw(87)( 72*8-1 downto  71*8), 
w73 => Pw(87)( 73*8-1 downto  72*8), w74 => Pw(87)( 74*8-1 downto  73*8), w75 => Pw(87)( 75*8-1 downto  74*8), w76 => Pw(87)( 76*8-1 downto  75*8), w77 => Pw(87)( 77*8-1 downto  76*8), w78 => Pw(87)( 78*8-1 downto  77*8), w79 => Pw(87)( 79*8-1 downto  78*8), w80 => Pw(87)( 80*8-1 downto  79*8), 
w81 => Pw(87)( 81*8-1 downto  80*8), w82 => Pw(87)( 82*8-1 downto  81*8), w83 => Pw(87)( 83*8-1 downto  82*8), w84 => Pw(87)( 84*8-1 downto  83*8), w85 => Pw(87)( 85*8-1 downto  84*8), w86 => Pw(87)( 86*8-1 downto  85*8), w87 => Pw(87)( 87*8-1 downto  86*8), w88 => Pw(87)( 88*8-1 downto  87*8), 
w89 => Pw(87)( 89*8-1 downto  88*8), w90 => Pw(87)( 90*8-1 downto  89*8), w91 => Pw(87)( 91*8-1 downto  90*8), w92 => Pw(87)( 92*8-1 downto  91*8), w93 => Pw(87)( 93*8-1 downto  92*8), w94 => Pw(87)( 94*8-1 downto  93*8), w95 => Pw(87)( 95*8-1 downto  94*8), w96 => Pw(87)( 96*8-1 downto  95*8), 
w97 => Pw(87)( 97*8-1 downto  96*8), w98 => Pw(87)( 98*8-1 downto  97*8), w99 => Pw(87)( 99*8-1 downto  98*8), w100=> Pw(87)(100*8-1 downto  99*8), w101=> Pw(87)(101*8-1 downto 100*8), w102=> Pw(87)(102*8-1 downto 101*8), w103=> Pw(87)(103*8-1 downto 102*8), w104=> Pw(87)(104*8-1 downto 103*8), 
w105=> Pw(87)(105*8-1 downto 104*8), w106=> Pw(87)(106*8-1 downto 105*8), w107=> Pw(87)(107*8-1 downto 106*8), w108=> Pw(87)(108*8-1 downto 107*8), w109=> Pw(87)(109*8-1 downto 108*8), w110=> Pw(87)(110*8-1 downto 109*8), w111=> Pw(87)(111*8-1 downto 110*8), w112=> Pw(87)(112*8-1 downto 111*8), 
w113=> Pw(87)(113*8-1 downto 112*8), w114=> Pw(87)(114*8-1 downto 113*8), w115=> Pw(87)(115*8-1 downto 114*8), w116=> Pw(87)(116*8-1 downto 115*8), w117=> Pw(87)(117*8-1 downto 116*8), w118=> Pw(87)(118*8-1 downto 117*8), w119=> Pw(87)(119*8-1 downto 118*8), w120=> Pw(87)(120*8-1 downto 119*8), 
w121=> Pw(87)(121*8-1 downto 120*8), w122=> Pw(87)(122*8-1 downto 121*8), w123=> Pw(87)(123*8-1 downto 122*8), w124=> Pw(87)(124*8-1 downto 123*8), w125=> Pw(87)(125*8-1 downto 124*8), w126=> Pw(87)(126*8-1 downto 125*8), w127=> Pw(87)(127*8-1 downto 126*8), w128=> Pw(87)(128*8-1 downto 127*8), 
           d_out   => pca_d87_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_88_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(88)(     7 downto    0),   w02 => Pw(88)( 2*8-1 downto    8),   w03 => Pw(88)( 3*8-1 downto  2*8),   w04 => Pw(88)( 4*8-1 downto  3*8),   w05 => Pw(88)( 5*8-1 downto  4*8),   w06 => Pw(88)( 6*8-1 downto  5*8),   w07 => Pw(88)( 7*8-1 downto  6*8),   w08 => Pw(88)( 8*8-1 downto  7*8),  
w09 => Pw(88)( 9*8-1 downto  8*8),   w10 => Pw(88)(10*8-1 downto  9*8),   w11 => Pw(88)(11*8-1 downto 10*8),   w12 => Pw(88)(12*8-1 downto 11*8),   w13 => Pw(88)(13*8-1 downto 12*8),   w14 => Pw(88)(14*8-1 downto 13*8),   w15 => Pw(88)(15*8-1 downto 14*8),   w16 => Pw(88)(16*8-1 downto 15*8),  
w17 => Pw(88)(17*8-1 downto 16*8),   w18 => Pw(88)(18*8-1 downto 17*8),   w19 => Pw(88)(19*8-1 downto 18*8),   w20 => Pw(88)(20*8-1 downto 19*8),   w21 => Pw(88)(21*8-1 downto 20*8),   w22 => Pw(88)(22*8-1 downto 21*8),   w23 => Pw(88)(23*8-1 downto 22*8),   w24 => Pw(88)(24*8-1 downto 23*8),  
w25 => Pw(88)(25*8-1 downto 24*8),   w26 => Pw(88)(26*8-1 downto 25*8),   w27 => Pw(88)(27*8-1 downto 26*8),   w28 => Pw(88)(28*8-1 downto 27*8),   w29 => Pw(88)(29*8-1 downto 28*8),   w30 => Pw(88)(30*8-1 downto 29*8),   w31 => Pw(88)(31*8-1 downto 30*8),   w32 => Pw(88)(32*8-1 downto 31*8),  
w33 => Pw(88)(33*8-1 downto 32*8),   w34 => Pw(88)(34*8-1 downto 33*8),   w35 => Pw(88)(35*8-1 downto 34*8),   w36 => Pw(88)(36*8-1 downto 35*8),   w37 => Pw(88)(37*8-1 downto 36*8),   w38 => Pw(88)(38*8-1 downto 37*8),   w39 => Pw(88)(39*8-1 downto 38*8),   w40 => Pw(88)(40*8-1 downto 39*8),  
w41 => Pw(88)(41*8-1 downto 40*8),   w42 => Pw(88)(42*8-1 downto 41*8),   w43 => Pw(88)(43*8-1 downto 42*8),   w44 => Pw(88)(44*8-1 downto 43*8),   w45 => Pw(88)(45*8-1 downto 44*8),   w46 => Pw(88)(46*8-1 downto 45*8),   w47 => Pw(88)(47*8-1 downto 46*8),   w48 => Pw(88)(48*8-1 downto 47*8),  
w49 => Pw(88)(49*8-1 downto 48*8),   w50 => Pw(88)(50*8-1 downto 49*8),   w51 => Pw(88)(51*8-1 downto 50*8),   w52 => Pw(88)(52*8-1 downto 51*8),   w53 => Pw(88)(53*8-1 downto 52*8),   w54 => Pw(88)(54*8-1 downto 53*8),   w55 => Pw(88)(55*8-1 downto 54*8),   w56 => Pw(88)(56*8-1 downto 55*8),  
w57 => Pw(88)(57*8-1 downto 56*8),   w58 => Pw(88)(58*8-1 downto 57*8),   w59 => Pw(88)(59*8-1 downto 58*8),   w60 => Pw(88)(60*8-1 downto 59*8),   w61 => Pw(88)(61*8-1 downto 60*8),   w62 => Pw(88)(62*8-1 downto 61*8),   w63 => Pw(88)(63*8-1 downto 62*8),   w64 => Pw(88)(64*8-1 downto 63*8), 
w65 => Pw(88)( 65*8-1 downto  64*8), w66 => Pw(88)( 66*8-1 downto  65*8), w67 => Pw(88)( 67*8-1 downto  66*8), w68 => Pw(88)( 68*8-1 downto  67*8), w69 => Pw(88)( 69*8-1 downto  68*8), w70 => Pw(88)( 70*8-1 downto  69*8), w71 => Pw(88)( 71*8-1 downto  70*8), w72 => Pw(88)( 72*8-1 downto  71*8), 
w73 => Pw(88)( 73*8-1 downto  72*8), w74 => Pw(88)( 74*8-1 downto  73*8), w75 => Pw(88)( 75*8-1 downto  74*8), w76 => Pw(88)( 76*8-1 downto  75*8), w77 => Pw(88)( 77*8-1 downto  76*8), w78 => Pw(88)( 78*8-1 downto  77*8), w79 => Pw(88)( 79*8-1 downto  78*8), w80 => Pw(88)( 80*8-1 downto  79*8), 
w81 => Pw(88)( 81*8-1 downto  80*8), w82 => Pw(88)( 82*8-1 downto  81*8), w83 => Pw(88)( 83*8-1 downto  82*8), w84 => Pw(88)( 84*8-1 downto  83*8), w85 => Pw(88)( 85*8-1 downto  84*8), w86 => Pw(88)( 86*8-1 downto  85*8), w87 => Pw(88)( 87*8-1 downto  86*8), w88 => Pw(88)( 88*8-1 downto  87*8), 
w89 => Pw(88)( 89*8-1 downto  88*8), w90 => Pw(88)( 90*8-1 downto  89*8), w91 => Pw(88)( 91*8-1 downto  90*8), w92 => Pw(88)( 92*8-1 downto  91*8), w93 => Pw(88)( 93*8-1 downto  92*8), w94 => Pw(88)( 94*8-1 downto  93*8), w95 => Pw(88)( 95*8-1 downto  94*8), w96 => Pw(88)( 96*8-1 downto  95*8), 
w97 => Pw(88)( 97*8-1 downto  96*8), w98 => Pw(88)( 98*8-1 downto  97*8), w99 => Pw(88)( 99*8-1 downto  98*8), w100=> Pw(88)(100*8-1 downto  99*8), w101=> Pw(88)(101*8-1 downto 100*8), w102=> Pw(88)(102*8-1 downto 101*8), w103=> Pw(88)(103*8-1 downto 102*8), w104=> Pw(88)(104*8-1 downto 103*8), 
w105=> Pw(88)(105*8-1 downto 104*8), w106=> Pw(88)(106*8-1 downto 105*8), w107=> Pw(88)(107*8-1 downto 106*8), w108=> Pw(88)(108*8-1 downto 107*8), w109=> Pw(88)(109*8-1 downto 108*8), w110=> Pw(88)(110*8-1 downto 109*8), w111=> Pw(88)(111*8-1 downto 110*8), w112=> Pw(88)(112*8-1 downto 111*8), 
w113=> Pw(88)(113*8-1 downto 112*8), w114=> Pw(88)(114*8-1 downto 113*8), w115=> Pw(88)(115*8-1 downto 114*8), w116=> Pw(88)(116*8-1 downto 115*8), w117=> Pw(88)(117*8-1 downto 116*8), w118=> Pw(88)(118*8-1 downto 117*8), w119=> Pw(88)(119*8-1 downto 118*8), w120=> Pw(88)(120*8-1 downto 119*8), 
w121=> Pw(88)(121*8-1 downto 120*8), w122=> Pw(88)(122*8-1 downto 121*8), w123=> Pw(88)(123*8-1 downto 122*8), w124=> Pw(88)(124*8-1 downto 123*8), w125=> Pw(88)(125*8-1 downto 124*8), w126=> Pw(88)(126*8-1 downto 125*8), w127=> Pw(88)(127*8-1 downto 126*8), w128=> Pw(88)(128*8-1 downto 127*8), 
           d_out   => pca_d88_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_89_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(89)(     7 downto    0),   w02 => Pw(89)( 2*8-1 downto    8),   w03 => Pw(89)( 3*8-1 downto  2*8),   w04 => Pw(89)( 4*8-1 downto  3*8),   w05 => Pw(89)( 5*8-1 downto  4*8),   w06 => Pw(89)( 6*8-1 downto  5*8),   w07 => Pw(89)( 7*8-1 downto  6*8),   w08 => Pw(89)( 8*8-1 downto  7*8),  
w09 => Pw(89)( 9*8-1 downto  8*8),   w10 => Pw(89)(10*8-1 downto  9*8),   w11 => Pw(89)(11*8-1 downto 10*8),   w12 => Pw(89)(12*8-1 downto 11*8),   w13 => Pw(89)(13*8-1 downto 12*8),   w14 => Pw(89)(14*8-1 downto 13*8),   w15 => Pw(89)(15*8-1 downto 14*8),   w16 => Pw(89)(16*8-1 downto 15*8),  
w17 => Pw(89)(17*8-1 downto 16*8),   w18 => Pw(89)(18*8-1 downto 17*8),   w19 => Pw(89)(19*8-1 downto 18*8),   w20 => Pw(89)(20*8-1 downto 19*8),   w21 => Pw(89)(21*8-1 downto 20*8),   w22 => Pw(89)(22*8-1 downto 21*8),   w23 => Pw(89)(23*8-1 downto 22*8),   w24 => Pw(89)(24*8-1 downto 23*8),  
w25 => Pw(89)(25*8-1 downto 24*8),   w26 => Pw(89)(26*8-1 downto 25*8),   w27 => Pw(89)(27*8-1 downto 26*8),   w28 => Pw(89)(28*8-1 downto 27*8),   w29 => Pw(89)(29*8-1 downto 28*8),   w30 => Pw(89)(30*8-1 downto 29*8),   w31 => Pw(89)(31*8-1 downto 30*8),   w32 => Pw(89)(32*8-1 downto 31*8),  
w33 => Pw(89)(33*8-1 downto 32*8),   w34 => Pw(89)(34*8-1 downto 33*8),   w35 => Pw(89)(35*8-1 downto 34*8),   w36 => Pw(89)(36*8-1 downto 35*8),   w37 => Pw(89)(37*8-1 downto 36*8),   w38 => Pw(89)(38*8-1 downto 37*8),   w39 => Pw(89)(39*8-1 downto 38*8),   w40 => Pw(89)(40*8-1 downto 39*8),  
w41 => Pw(89)(41*8-1 downto 40*8),   w42 => Pw(89)(42*8-1 downto 41*8),   w43 => Pw(89)(43*8-1 downto 42*8),   w44 => Pw(89)(44*8-1 downto 43*8),   w45 => Pw(89)(45*8-1 downto 44*8),   w46 => Pw(89)(46*8-1 downto 45*8),   w47 => Pw(89)(47*8-1 downto 46*8),   w48 => Pw(89)(48*8-1 downto 47*8),  
w49 => Pw(89)(49*8-1 downto 48*8),   w50 => Pw(89)(50*8-1 downto 49*8),   w51 => Pw(89)(51*8-1 downto 50*8),   w52 => Pw(89)(52*8-1 downto 51*8),   w53 => Pw(89)(53*8-1 downto 52*8),   w54 => Pw(89)(54*8-1 downto 53*8),   w55 => Pw(89)(55*8-1 downto 54*8),   w56 => Pw(89)(56*8-1 downto 55*8),  
w57 => Pw(89)(57*8-1 downto 56*8),   w58 => Pw(89)(58*8-1 downto 57*8),   w59 => Pw(89)(59*8-1 downto 58*8),   w60 => Pw(89)(60*8-1 downto 59*8),   w61 => Pw(89)(61*8-1 downto 60*8),   w62 => Pw(89)(62*8-1 downto 61*8),   w63 => Pw(89)(63*8-1 downto 62*8),   w64 => Pw(89)(64*8-1 downto 63*8), 
w65 => Pw(89)( 65*8-1 downto  64*8), w66 => Pw(89)( 66*8-1 downto  65*8), w67 => Pw(89)( 67*8-1 downto  66*8), w68 => Pw(89)( 68*8-1 downto  67*8), w69 => Pw(89)( 69*8-1 downto  68*8), w70 => Pw(89)( 70*8-1 downto  69*8), w71 => Pw(89)( 71*8-1 downto  70*8), w72 => Pw(89)( 72*8-1 downto  71*8), 
w73 => Pw(89)( 73*8-1 downto  72*8), w74 => Pw(89)( 74*8-1 downto  73*8), w75 => Pw(89)( 75*8-1 downto  74*8), w76 => Pw(89)( 76*8-1 downto  75*8), w77 => Pw(89)( 77*8-1 downto  76*8), w78 => Pw(89)( 78*8-1 downto  77*8), w79 => Pw(89)( 79*8-1 downto  78*8), w80 => Pw(89)( 80*8-1 downto  79*8), 
w81 => Pw(89)( 81*8-1 downto  80*8), w82 => Pw(89)( 82*8-1 downto  81*8), w83 => Pw(89)( 83*8-1 downto  82*8), w84 => Pw(89)( 84*8-1 downto  83*8), w85 => Pw(89)( 85*8-1 downto  84*8), w86 => Pw(89)( 86*8-1 downto  85*8), w87 => Pw(89)( 87*8-1 downto  86*8), w88 => Pw(89)( 88*8-1 downto  87*8), 
w89 => Pw(89)( 89*8-1 downto  88*8), w90 => Pw(89)( 90*8-1 downto  89*8), w91 => Pw(89)( 91*8-1 downto  90*8), w92 => Pw(89)( 92*8-1 downto  91*8), w93 => Pw(89)( 93*8-1 downto  92*8), w94 => Pw(89)( 94*8-1 downto  93*8), w95 => Pw(89)( 95*8-1 downto  94*8), w96 => Pw(89)( 96*8-1 downto  95*8), 
w97 => Pw(89)( 97*8-1 downto  96*8), w98 => Pw(89)( 98*8-1 downto  97*8), w99 => Pw(89)( 99*8-1 downto  98*8), w100=> Pw(89)(100*8-1 downto  99*8), w101=> Pw(89)(101*8-1 downto 100*8), w102=> Pw(89)(102*8-1 downto 101*8), w103=> Pw(89)(103*8-1 downto 102*8), w104=> Pw(89)(104*8-1 downto 103*8), 
w105=> Pw(89)(105*8-1 downto 104*8), w106=> Pw(89)(106*8-1 downto 105*8), w107=> Pw(89)(107*8-1 downto 106*8), w108=> Pw(89)(108*8-1 downto 107*8), w109=> Pw(89)(109*8-1 downto 108*8), w110=> Pw(89)(110*8-1 downto 109*8), w111=> Pw(89)(111*8-1 downto 110*8), w112=> Pw(89)(112*8-1 downto 111*8), 
w113=> Pw(89)(113*8-1 downto 112*8), w114=> Pw(89)(114*8-1 downto 113*8), w115=> Pw(89)(115*8-1 downto 114*8), w116=> Pw(89)(116*8-1 downto 115*8), w117=> Pw(89)(117*8-1 downto 116*8), w118=> Pw(89)(118*8-1 downto 117*8), w119=> Pw(89)(119*8-1 downto 118*8), w120=> Pw(89)(120*8-1 downto 119*8), 
w121=> Pw(89)(121*8-1 downto 120*8), w122=> Pw(89)(122*8-1 downto 121*8), w123=> Pw(89)(123*8-1 downto 122*8), w124=> Pw(89)(124*8-1 downto 123*8), w125=> Pw(89)(125*8-1 downto 124*8), w126=> Pw(89)(126*8-1 downto 125*8), w127=> Pw(89)(127*8-1 downto 126*8), w128=> Pw(89)(128*8-1 downto 127*8), 
           d_out   => pca_d89_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_90_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(90)(     7 downto    0),   w02 => Pw(90)( 2*8-1 downto    8),   w03 => Pw(90)( 3*8-1 downto  2*8),   w04 => Pw(90)( 4*8-1 downto  3*8),   w05 => Pw(90)( 5*8-1 downto  4*8),   w06 => Pw(90)( 6*8-1 downto  5*8),   w07 => Pw(90)( 7*8-1 downto  6*8),   w08 => Pw(90)( 8*8-1 downto  7*8),  
w09 => Pw(90)( 9*8-1 downto  8*8),   w10 => Pw(90)(10*8-1 downto  9*8),   w11 => Pw(90)(11*8-1 downto 10*8),   w12 => Pw(90)(12*8-1 downto 11*8),   w13 => Pw(90)(13*8-1 downto 12*8),   w14 => Pw(90)(14*8-1 downto 13*8),   w15 => Pw(90)(15*8-1 downto 14*8),   w16 => Pw(90)(16*8-1 downto 15*8),  
w17 => Pw(90)(17*8-1 downto 16*8),   w18 => Pw(90)(18*8-1 downto 17*8),   w19 => Pw(90)(19*8-1 downto 18*8),   w20 => Pw(90)(20*8-1 downto 19*8),   w21 => Pw(90)(21*8-1 downto 20*8),   w22 => Pw(90)(22*8-1 downto 21*8),   w23 => Pw(90)(23*8-1 downto 22*8),   w24 => Pw(90)(24*8-1 downto 23*8),  
w25 => Pw(90)(25*8-1 downto 24*8),   w26 => Pw(90)(26*8-1 downto 25*8),   w27 => Pw(90)(27*8-1 downto 26*8),   w28 => Pw(90)(28*8-1 downto 27*8),   w29 => Pw(90)(29*8-1 downto 28*8),   w30 => Pw(90)(30*8-1 downto 29*8),   w31 => Pw(90)(31*8-1 downto 30*8),   w32 => Pw(90)(32*8-1 downto 31*8),  
w33 => Pw(90)(33*8-1 downto 32*8),   w34 => Pw(90)(34*8-1 downto 33*8),   w35 => Pw(90)(35*8-1 downto 34*8),   w36 => Pw(90)(36*8-1 downto 35*8),   w37 => Pw(90)(37*8-1 downto 36*8),   w38 => Pw(90)(38*8-1 downto 37*8),   w39 => Pw(90)(39*8-1 downto 38*8),   w40 => Pw(90)(40*8-1 downto 39*8),  
w41 => Pw(90)(41*8-1 downto 40*8),   w42 => Pw(90)(42*8-1 downto 41*8),   w43 => Pw(90)(43*8-1 downto 42*8),   w44 => Pw(90)(44*8-1 downto 43*8),   w45 => Pw(90)(45*8-1 downto 44*8),   w46 => Pw(90)(46*8-1 downto 45*8),   w47 => Pw(90)(47*8-1 downto 46*8),   w48 => Pw(90)(48*8-1 downto 47*8),  
w49 => Pw(90)(49*8-1 downto 48*8),   w50 => Pw(90)(50*8-1 downto 49*8),   w51 => Pw(90)(51*8-1 downto 50*8),   w52 => Pw(90)(52*8-1 downto 51*8),   w53 => Pw(90)(53*8-1 downto 52*8),   w54 => Pw(90)(54*8-1 downto 53*8),   w55 => Pw(90)(55*8-1 downto 54*8),   w56 => Pw(90)(56*8-1 downto 55*8),  
w57 => Pw(90)(57*8-1 downto 56*8),   w58 => Pw(90)(58*8-1 downto 57*8),   w59 => Pw(90)(59*8-1 downto 58*8),   w60 => Pw(90)(60*8-1 downto 59*8),   w61 => Pw(90)(61*8-1 downto 60*8),   w62 => Pw(90)(62*8-1 downto 61*8),   w63 => Pw(90)(63*8-1 downto 62*8),   w64 => Pw(90)(64*8-1 downto 63*8), 
w65 => Pw(90)( 65*8-1 downto  64*8), w66 => Pw(90)( 66*8-1 downto  65*8), w67 => Pw(90)( 67*8-1 downto  66*8), w68 => Pw(90)( 68*8-1 downto  67*8), w69 => Pw(90)( 69*8-1 downto  68*8), w70 => Pw(90)( 70*8-1 downto  69*8), w71 => Pw(90)( 71*8-1 downto  70*8), w72 => Pw(90)( 72*8-1 downto  71*8), 
w73 => Pw(90)( 73*8-1 downto  72*8), w74 => Pw(90)( 74*8-1 downto  73*8), w75 => Pw(90)( 75*8-1 downto  74*8), w76 => Pw(90)( 76*8-1 downto  75*8), w77 => Pw(90)( 77*8-1 downto  76*8), w78 => Pw(90)( 78*8-1 downto  77*8), w79 => Pw(90)( 79*8-1 downto  78*8), w80 => Pw(90)( 80*8-1 downto  79*8), 
w81 => Pw(90)( 81*8-1 downto  80*8), w82 => Pw(90)( 82*8-1 downto  81*8), w83 => Pw(90)( 83*8-1 downto  82*8), w84 => Pw(90)( 84*8-1 downto  83*8), w85 => Pw(90)( 85*8-1 downto  84*8), w86 => Pw(90)( 86*8-1 downto  85*8), w87 => Pw(90)( 87*8-1 downto  86*8), w88 => Pw(90)( 88*8-1 downto  87*8), 
w89 => Pw(90)( 89*8-1 downto  88*8), w90 => Pw(90)( 90*8-1 downto  89*8), w91 => Pw(90)( 91*8-1 downto  90*8), w92 => Pw(90)( 92*8-1 downto  91*8), w93 => Pw(90)( 93*8-1 downto  92*8), w94 => Pw(90)( 94*8-1 downto  93*8), w95 => Pw(90)( 95*8-1 downto  94*8), w96 => Pw(90)( 96*8-1 downto  95*8), 
w97 => Pw(90)( 97*8-1 downto  96*8), w98 => Pw(90)( 98*8-1 downto  97*8), w99 => Pw(90)( 99*8-1 downto  98*8), w100=> Pw(90)(100*8-1 downto  99*8), w101=> Pw(90)(101*8-1 downto 100*8), w102=> Pw(90)(102*8-1 downto 101*8), w103=> Pw(90)(103*8-1 downto 102*8), w104=> Pw(90)(104*8-1 downto 103*8), 
w105=> Pw(90)(105*8-1 downto 104*8), w106=> Pw(90)(106*8-1 downto 105*8), w107=> Pw(90)(107*8-1 downto 106*8), w108=> Pw(90)(108*8-1 downto 107*8), w109=> Pw(90)(109*8-1 downto 108*8), w110=> Pw(90)(110*8-1 downto 109*8), w111=> Pw(90)(111*8-1 downto 110*8), w112=> Pw(90)(112*8-1 downto 111*8), 
w113=> Pw(90)(113*8-1 downto 112*8), w114=> Pw(90)(114*8-1 downto 113*8), w115=> Pw(90)(115*8-1 downto 114*8), w116=> Pw(90)(116*8-1 downto 115*8), w117=> Pw(90)(117*8-1 downto 116*8), w118=> Pw(90)(118*8-1 downto 117*8), w119=> Pw(90)(119*8-1 downto 118*8), w120=> Pw(90)(120*8-1 downto 119*8), 
w121=> Pw(90)(121*8-1 downto 120*8), w122=> Pw(90)(122*8-1 downto 121*8), w123=> Pw(90)(123*8-1 downto 122*8), w124=> Pw(90)(124*8-1 downto 123*8), w125=> Pw(90)(125*8-1 downto 124*8), w126=> Pw(90)(126*8-1 downto 125*8), w127=> Pw(90)(127*8-1 downto 126*8), w128=> Pw(90)(128*8-1 downto 127*8), 
           d_out   => pca_d90_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_91_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(91)(     7 downto    0),   w02 => Pw(91)( 2*8-1 downto    8),   w03 => Pw(91)( 3*8-1 downto  2*8),   w04 => Pw(91)( 4*8-1 downto  3*8),   w05 => Pw(91)( 5*8-1 downto  4*8),   w06 => Pw(91)( 6*8-1 downto  5*8),   w07 => Pw(91)( 7*8-1 downto  6*8),   w08 => Pw(91)( 8*8-1 downto  7*8),  
w09 => Pw(91)( 9*8-1 downto  8*8),   w10 => Pw(91)(10*8-1 downto  9*8),   w11 => Pw(91)(11*8-1 downto 10*8),   w12 => Pw(91)(12*8-1 downto 11*8),   w13 => Pw(91)(13*8-1 downto 12*8),   w14 => Pw(91)(14*8-1 downto 13*8),   w15 => Pw(91)(15*8-1 downto 14*8),   w16 => Pw(91)(16*8-1 downto 15*8),  
w17 => Pw(91)(17*8-1 downto 16*8),   w18 => Pw(91)(18*8-1 downto 17*8),   w19 => Pw(91)(19*8-1 downto 18*8),   w20 => Pw(91)(20*8-1 downto 19*8),   w21 => Pw(91)(21*8-1 downto 20*8),   w22 => Pw(91)(22*8-1 downto 21*8),   w23 => Pw(91)(23*8-1 downto 22*8),   w24 => Pw(91)(24*8-1 downto 23*8),  
w25 => Pw(91)(25*8-1 downto 24*8),   w26 => Pw(91)(26*8-1 downto 25*8),   w27 => Pw(91)(27*8-1 downto 26*8),   w28 => Pw(91)(28*8-1 downto 27*8),   w29 => Pw(91)(29*8-1 downto 28*8),   w30 => Pw(91)(30*8-1 downto 29*8),   w31 => Pw(91)(31*8-1 downto 30*8),   w32 => Pw(91)(32*8-1 downto 31*8),  
w33 => Pw(91)(33*8-1 downto 32*8),   w34 => Pw(91)(34*8-1 downto 33*8),   w35 => Pw(91)(35*8-1 downto 34*8),   w36 => Pw(91)(36*8-1 downto 35*8),   w37 => Pw(91)(37*8-1 downto 36*8),   w38 => Pw(91)(38*8-1 downto 37*8),   w39 => Pw(91)(39*8-1 downto 38*8),   w40 => Pw(91)(40*8-1 downto 39*8),  
w41 => Pw(91)(41*8-1 downto 40*8),   w42 => Pw(91)(42*8-1 downto 41*8),   w43 => Pw(91)(43*8-1 downto 42*8),   w44 => Pw(91)(44*8-1 downto 43*8),   w45 => Pw(91)(45*8-1 downto 44*8),   w46 => Pw(91)(46*8-1 downto 45*8),   w47 => Pw(91)(47*8-1 downto 46*8),   w48 => Pw(91)(48*8-1 downto 47*8),  
w49 => Pw(91)(49*8-1 downto 48*8),   w50 => Pw(91)(50*8-1 downto 49*8),   w51 => Pw(91)(51*8-1 downto 50*8),   w52 => Pw(91)(52*8-1 downto 51*8),   w53 => Pw(91)(53*8-1 downto 52*8),   w54 => Pw(91)(54*8-1 downto 53*8),   w55 => Pw(91)(55*8-1 downto 54*8),   w56 => Pw(91)(56*8-1 downto 55*8),  
w57 => Pw(91)(57*8-1 downto 56*8),   w58 => Pw(91)(58*8-1 downto 57*8),   w59 => Pw(91)(59*8-1 downto 58*8),   w60 => Pw(91)(60*8-1 downto 59*8),   w61 => Pw(91)(61*8-1 downto 60*8),   w62 => Pw(91)(62*8-1 downto 61*8),   w63 => Pw(91)(63*8-1 downto 62*8),   w64 => Pw(91)(64*8-1 downto 63*8), 
w65 => Pw(91)( 65*8-1 downto  64*8), w66 => Pw(91)( 66*8-1 downto  65*8), w67 => Pw(91)( 67*8-1 downto  66*8), w68 => Pw(91)( 68*8-1 downto  67*8), w69 => Pw(91)( 69*8-1 downto  68*8), w70 => Pw(91)( 70*8-1 downto  69*8), w71 => Pw(91)( 71*8-1 downto  70*8), w72 => Pw(91)( 72*8-1 downto  71*8), 
w73 => Pw(91)( 73*8-1 downto  72*8), w74 => Pw(91)( 74*8-1 downto  73*8), w75 => Pw(91)( 75*8-1 downto  74*8), w76 => Pw(91)( 76*8-1 downto  75*8), w77 => Pw(91)( 77*8-1 downto  76*8), w78 => Pw(91)( 78*8-1 downto  77*8), w79 => Pw(91)( 79*8-1 downto  78*8), w80 => Pw(91)( 80*8-1 downto  79*8), 
w81 => Pw(91)( 81*8-1 downto  80*8), w82 => Pw(91)( 82*8-1 downto  81*8), w83 => Pw(91)( 83*8-1 downto  82*8), w84 => Pw(91)( 84*8-1 downto  83*8), w85 => Pw(91)( 85*8-1 downto  84*8), w86 => Pw(91)( 86*8-1 downto  85*8), w87 => Pw(91)( 87*8-1 downto  86*8), w88 => Pw(91)( 88*8-1 downto  87*8), 
w89 => Pw(91)( 89*8-1 downto  88*8), w90 => Pw(91)( 90*8-1 downto  89*8), w91 => Pw(91)( 91*8-1 downto  90*8), w92 => Pw(91)( 92*8-1 downto  91*8), w93 => Pw(91)( 93*8-1 downto  92*8), w94 => Pw(91)( 94*8-1 downto  93*8), w95 => Pw(91)( 95*8-1 downto  94*8), w96 => Pw(91)( 96*8-1 downto  95*8), 
w97 => Pw(91)( 97*8-1 downto  96*8), w98 => Pw(91)( 98*8-1 downto  97*8), w99 => Pw(91)( 99*8-1 downto  98*8), w100=> Pw(91)(100*8-1 downto  99*8), w101=> Pw(91)(101*8-1 downto 100*8), w102=> Pw(91)(102*8-1 downto 101*8), w103=> Pw(91)(103*8-1 downto 102*8), w104=> Pw(91)(104*8-1 downto 103*8), 
w105=> Pw(91)(105*8-1 downto 104*8), w106=> Pw(91)(106*8-1 downto 105*8), w107=> Pw(91)(107*8-1 downto 106*8), w108=> Pw(91)(108*8-1 downto 107*8), w109=> Pw(91)(109*8-1 downto 108*8), w110=> Pw(91)(110*8-1 downto 109*8), w111=> Pw(91)(111*8-1 downto 110*8), w112=> Pw(91)(112*8-1 downto 111*8), 
w113=> Pw(91)(113*8-1 downto 112*8), w114=> Pw(91)(114*8-1 downto 113*8), w115=> Pw(91)(115*8-1 downto 114*8), w116=> Pw(91)(116*8-1 downto 115*8), w117=> Pw(91)(117*8-1 downto 116*8), w118=> Pw(91)(118*8-1 downto 117*8), w119=> Pw(91)(119*8-1 downto 118*8), w120=> Pw(91)(120*8-1 downto 119*8), 
w121=> Pw(91)(121*8-1 downto 120*8), w122=> Pw(91)(122*8-1 downto 121*8), w123=> Pw(91)(123*8-1 downto 122*8), w124=> Pw(91)(124*8-1 downto 123*8), w125=> Pw(91)(125*8-1 downto 124*8), w126=> Pw(91)(126*8-1 downto 125*8), w127=> Pw(91)(127*8-1 downto 126*8), w128=> Pw(91)(128*8-1 downto 127*8), 
           d_out   => pca_d91_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_92_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(92)(     7 downto    0),   w02 => Pw(92)( 2*8-1 downto    8),   w03 => Pw(92)( 3*8-1 downto  2*8),   w04 => Pw(92)( 4*8-1 downto  3*8),   w05 => Pw(92)( 5*8-1 downto  4*8),   w06 => Pw(92)( 6*8-1 downto  5*8),   w07 => Pw(92)( 7*8-1 downto  6*8),   w08 => Pw(92)( 8*8-1 downto  7*8),  
w09 => Pw(92)( 9*8-1 downto  8*8),   w10 => Pw(92)(10*8-1 downto  9*8),   w11 => Pw(92)(11*8-1 downto 10*8),   w12 => Pw(92)(12*8-1 downto 11*8),   w13 => Pw(92)(13*8-1 downto 12*8),   w14 => Pw(92)(14*8-1 downto 13*8),   w15 => Pw(92)(15*8-1 downto 14*8),   w16 => Pw(92)(16*8-1 downto 15*8),  
w17 => Pw(92)(17*8-1 downto 16*8),   w18 => Pw(92)(18*8-1 downto 17*8),   w19 => Pw(92)(19*8-1 downto 18*8),   w20 => Pw(92)(20*8-1 downto 19*8),   w21 => Pw(92)(21*8-1 downto 20*8),   w22 => Pw(92)(22*8-1 downto 21*8),   w23 => Pw(92)(23*8-1 downto 22*8),   w24 => Pw(92)(24*8-1 downto 23*8),  
w25 => Pw(92)(25*8-1 downto 24*8),   w26 => Pw(92)(26*8-1 downto 25*8),   w27 => Pw(92)(27*8-1 downto 26*8),   w28 => Pw(92)(28*8-1 downto 27*8),   w29 => Pw(92)(29*8-1 downto 28*8),   w30 => Pw(92)(30*8-1 downto 29*8),   w31 => Pw(92)(31*8-1 downto 30*8),   w32 => Pw(92)(32*8-1 downto 31*8),  
w33 => Pw(92)(33*8-1 downto 32*8),   w34 => Pw(92)(34*8-1 downto 33*8),   w35 => Pw(92)(35*8-1 downto 34*8),   w36 => Pw(92)(36*8-1 downto 35*8),   w37 => Pw(92)(37*8-1 downto 36*8),   w38 => Pw(92)(38*8-1 downto 37*8),   w39 => Pw(92)(39*8-1 downto 38*8),   w40 => Pw(92)(40*8-1 downto 39*8),  
w41 => Pw(92)(41*8-1 downto 40*8),   w42 => Pw(92)(42*8-1 downto 41*8),   w43 => Pw(92)(43*8-1 downto 42*8),   w44 => Pw(92)(44*8-1 downto 43*8),   w45 => Pw(92)(45*8-1 downto 44*8),   w46 => Pw(92)(46*8-1 downto 45*8),   w47 => Pw(92)(47*8-1 downto 46*8),   w48 => Pw(92)(48*8-1 downto 47*8),  
w49 => Pw(92)(49*8-1 downto 48*8),   w50 => Pw(92)(50*8-1 downto 49*8),   w51 => Pw(92)(51*8-1 downto 50*8),   w52 => Pw(92)(52*8-1 downto 51*8),   w53 => Pw(92)(53*8-1 downto 52*8),   w54 => Pw(92)(54*8-1 downto 53*8),   w55 => Pw(92)(55*8-1 downto 54*8),   w56 => Pw(92)(56*8-1 downto 55*8),  
w57 => Pw(92)(57*8-1 downto 56*8),   w58 => Pw(92)(58*8-1 downto 57*8),   w59 => Pw(92)(59*8-1 downto 58*8),   w60 => Pw(92)(60*8-1 downto 59*8),   w61 => Pw(92)(61*8-1 downto 60*8),   w62 => Pw(92)(62*8-1 downto 61*8),   w63 => Pw(92)(63*8-1 downto 62*8),   w64 => Pw(92)(64*8-1 downto 63*8), 
w65 => Pw(92)( 65*8-1 downto  64*8), w66 => Pw(92)( 66*8-1 downto  65*8), w67 => Pw(92)( 67*8-1 downto  66*8), w68 => Pw(92)( 68*8-1 downto  67*8), w69 => Pw(92)( 69*8-1 downto  68*8), w70 => Pw(92)( 70*8-1 downto  69*8), w71 => Pw(92)( 71*8-1 downto  70*8), w72 => Pw(92)( 72*8-1 downto  71*8), 
w73 => Pw(92)( 73*8-1 downto  72*8), w74 => Pw(92)( 74*8-1 downto  73*8), w75 => Pw(92)( 75*8-1 downto  74*8), w76 => Pw(92)( 76*8-1 downto  75*8), w77 => Pw(92)( 77*8-1 downto  76*8), w78 => Pw(92)( 78*8-1 downto  77*8), w79 => Pw(92)( 79*8-1 downto  78*8), w80 => Pw(92)( 80*8-1 downto  79*8), 
w81 => Pw(92)( 81*8-1 downto  80*8), w82 => Pw(92)( 82*8-1 downto  81*8), w83 => Pw(92)( 83*8-1 downto  82*8), w84 => Pw(92)( 84*8-1 downto  83*8), w85 => Pw(92)( 85*8-1 downto  84*8), w86 => Pw(92)( 86*8-1 downto  85*8), w87 => Pw(92)( 87*8-1 downto  86*8), w88 => Pw(92)( 88*8-1 downto  87*8), 
w89 => Pw(92)( 89*8-1 downto  88*8), w90 => Pw(92)( 90*8-1 downto  89*8), w91 => Pw(92)( 91*8-1 downto  90*8), w92 => Pw(92)( 92*8-1 downto  91*8), w93 => Pw(92)( 93*8-1 downto  92*8), w94 => Pw(92)( 94*8-1 downto  93*8), w95 => Pw(92)( 95*8-1 downto  94*8), w96 => Pw(92)( 96*8-1 downto  95*8), 
w97 => Pw(92)( 97*8-1 downto  96*8), w98 => Pw(92)( 98*8-1 downto  97*8), w99 => Pw(92)( 99*8-1 downto  98*8), w100=> Pw(92)(100*8-1 downto  99*8), w101=> Pw(92)(101*8-1 downto 100*8), w102=> Pw(92)(102*8-1 downto 101*8), w103=> Pw(92)(103*8-1 downto 102*8), w104=> Pw(92)(104*8-1 downto 103*8), 
w105=> Pw(92)(105*8-1 downto 104*8), w106=> Pw(92)(106*8-1 downto 105*8), w107=> Pw(92)(107*8-1 downto 106*8), w108=> Pw(92)(108*8-1 downto 107*8), w109=> Pw(92)(109*8-1 downto 108*8), w110=> Pw(92)(110*8-1 downto 109*8), w111=> Pw(92)(111*8-1 downto 110*8), w112=> Pw(92)(112*8-1 downto 111*8), 
w113=> Pw(92)(113*8-1 downto 112*8), w114=> Pw(92)(114*8-1 downto 113*8), w115=> Pw(92)(115*8-1 downto 114*8), w116=> Pw(92)(116*8-1 downto 115*8), w117=> Pw(92)(117*8-1 downto 116*8), w118=> Pw(92)(118*8-1 downto 117*8), w119=> Pw(92)(119*8-1 downto 118*8), w120=> Pw(92)(120*8-1 downto 119*8), 
w121=> Pw(92)(121*8-1 downto 120*8), w122=> Pw(92)(122*8-1 downto 121*8), w123=> Pw(92)(123*8-1 downto 122*8), w124=> Pw(92)(124*8-1 downto 123*8), w125=> Pw(92)(125*8-1 downto 124*8), w126=> Pw(92)(126*8-1 downto 125*8), w127=> Pw(92)(127*8-1 downto 126*8), w128=> Pw(92)(128*8-1 downto 127*8), 
           d_out   => pca_d92_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_93_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(93)(     7 downto    0),   w02 => Pw(93)( 2*8-1 downto    8),   w03 => Pw(93)( 3*8-1 downto  2*8),   w04 => Pw(93)( 4*8-1 downto  3*8),  w05 => Pw(93)( 5*8-1 downto  4*8),   w06 => Pw(93)( 6*8-1 downto  5*8),   w07 => Pw(93)( 7*8-1 downto  6*8),   w08 => Pw(93)( 8*8-1 downto  7*8),  
w09 => Pw(93)( 9*8-1 downto  8*8),   w10 => Pw(93)(10*8-1 downto  9*8),   w11 => Pw(93)(11*8-1 downto 10*8),   w12 => Pw(93)(12*8-1 downto 11*8),   w13 => Pw(93)(13*8-1 downto 12*8),   w14 => Pw(93)(14*8-1 downto 13*8),   w15 => Pw(93)(15*8-1 downto 14*8),   w16 => Pw(93)(16*8-1 downto 15*8),  
w17 => Pw(93)(17*8-1 downto 16*8),   w18 => Pw(93)(18*8-1 downto 17*8),   w19 => Pw(93)(19*8-1 downto 18*8),   w20 => Pw(93)(20*8-1 downto 19*8),   w21 => Pw(93)(21*8-1 downto 20*8),   w22 => Pw(93)(22*8-1 downto 21*8),   w23 => Pw(93)(23*8-1 downto 22*8),   w24 => Pw(93)(24*8-1 downto 23*8),  
w25 => Pw(93)(25*8-1 downto 24*8),   w26 => Pw(93)(26*8-1 downto 25*8),   w27 => Pw(93)(27*8-1 downto 26*8),   w28 => Pw(93)(28*8-1 downto 27*8),   w29 => Pw(93)(29*8-1 downto 28*8),   w30 => Pw(93)(30*8-1 downto 29*8),   w31 => Pw(93)(31*8-1 downto 30*8),   w32 => Pw(93)(32*8-1 downto 31*8),  
w33 => Pw(93)(33*8-1 downto 32*8),   w34 => Pw(93)(34*8-1 downto 33*8),   w35 => Pw(93)(35*8-1 downto 34*8),   w36 => Pw(93)(36*8-1 downto 35*8),   w37 => Pw(93)(37*8-1 downto 36*8),   w38 => Pw(93)(38*8-1 downto 37*8),   w39 => Pw(93)(39*8-1 downto 38*8),   w40 => Pw(93)(40*8-1 downto 39*8),  
w41 => Pw(93)(41*8-1 downto 40*8),   w42 => Pw(93)(42*8-1 downto 41*8),   w43 => Pw(93)(43*8-1 downto 42*8),   w44 => Pw(93)(44*8-1 downto 43*8),   w45 => Pw(93)(45*8-1 downto 44*8),   w46 => Pw(93)(46*8-1 downto 45*8),   w47 => Pw(93)(47*8-1 downto 46*8),   w48 => Pw(93)(48*8-1 downto 47*8),  
w49 => Pw(93)(49*8-1 downto 48*8),   w50 => Pw(93)(50*8-1 downto 49*8),   w51 => Pw(93)(51*8-1 downto 50*8),   w52 => Pw(93)(52*8-1 downto 51*8),   w53 => Pw(93)(53*8-1 downto 52*8),   w54 => Pw(93)(54*8-1 downto 53*8),   w55 => Pw(93)(55*8-1 downto 54*8),   w56 => Pw(93)(56*8-1 downto 55*8),  
w57 => Pw(93)(57*8-1 downto 56*8),   w58 => Pw(93)(58*8-1 downto 57*8),   w59 => Pw(93)(59*8-1 downto 58*8),   w60 => Pw(93)(60*8-1 downto 59*8),   w61 => Pw(93)(61*8-1 downto 60*8),   w62 => Pw(93)(62*8-1 downto 61*8),   w63 => Pw(93)(63*8-1 downto 62*8),   w64 => Pw(93)(64*8-1 downto 63*8), 
w65 => Pw(93)( 65*8-1 downto  64*8), w66 => Pw(93)( 66*8-1 downto  65*8), w67 => Pw(93)( 67*8-1 downto  66*8), w68 => Pw(93)( 68*8-1 downto  67*8), w69 => Pw(93)( 69*8-1 downto  68*8), w70 => Pw(93)( 70*8-1 downto  69*8), w71 => Pw(93)( 71*8-1 downto  70*8), w72 => Pw(93)( 72*8-1 downto  71*8), 
w73 => Pw(93)( 73*8-1 downto  72*8), w74 => Pw(93)( 74*8-1 downto  73*8), w75 => Pw(93)( 75*8-1 downto  74*8), w76 => Pw(93)( 76*8-1 downto  75*8), w77 => Pw(93)( 77*8-1 downto  76*8), w78 => Pw(93)( 78*8-1 downto  77*8), w79 => Pw(93)( 79*8-1 downto  78*8), w80 => Pw(93)( 80*8-1 downto  79*8), 
w81 => Pw(93)( 81*8-1 downto  80*8), w82 => Pw(93)( 82*8-1 downto  81*8), w83 => Pw(93)( 83*8-1 downto  82*8), w84 => Pw(93)( 84*8-1 downto  83*8), w85 => Pw(93)( 85*8-1 downto  84*8), w86 => Pw(93)( 86*8-1 downto  85*8), w87 => Pw(93)( 87*8-1 downto  86*8), w88 => Pw(93)( 88*8-1 downto  87*8), 
w89 => Pw(93)( 89*8-1 downto  88*8), w90 => Pw(93)( 90*8-1 downto  89*8), w91 => Pw(93)( 91*8-1 downto  90*8), w92 => Pw(93)( 92*8-1 downto  91*8), w93 => Pw(93)( 93*8-1 downto  92*8), w94 => Pw(93)( 94*8-1 downto  93*8), w95 => Pw(93)( 95*8-1 downto  94*8), w96 => Pw(93)( 96*8-1 downto  95*8), 
w97 => Pw(93)( 97*8-1 downto  96*8), w98 => Pw(93)( 98*8-1 downto  97*8), w99 => Pw(93)( 99*8-1 downto  98*8), w100=> Pw(93)(100*8-1 downto  99*8), w101=> Pw(93)(101*8-1 downto 100*8), w102=> Pw(93)(102*8-1 downto 101*8), w103=> Pw(93)(103*8-1 downto 102*8), w104=> Pw(93)(104*8-1 downto 103*8), 
w105=> Pw(93)(105*8-1 downto 104*8), w106=> Pw(93)(106*8-1 downto 105*8), w107=> Pw(93)(107*8-1 downto 106*8), w108=> Pw(93)(108*8-1 downto 107*8), w109=> Pw(93)(109*8-1 downto 108*8), w110=> Pw(93)(110*8-1 downto 109*8), w111=> Pw(93)(111*8-1 downto 110*8), w112=> Pw(93)(112*8-1 downto 111*8), 
w113=> Pw(93)(113*8-1 downto 112*8), w114=> Pw(93)(114*8-1 downto 113*8), w115=> Pw(93)(115*8-1 downto 114*8), w116=> Pw(93)(116*8-1 downto 115*8), w117=> Pw(93)(117*8-1 downto 116*8), w118=> Pw(93)(118*8-1 downto 117*8), w119=> Pw(93)(119*8-1 downto 118*8), w120=> Pw(93)(120*8-1 downto 119*8), 
w121=> Pw(93)(121*8-1 downto 120*8), w122=> Pw(93)(122*8-1 downto 121*8), w123=> Pw(93)(123*8-1 downto 122*8), w124=> Pw(93)(124*8-1 downto 123*8), w125=> Pw(93)(125*8-1 downto 124*8), w126=> Pw(93)(126*8-1 downto 125*8), w127=> Pw(93)(127*8-1 downto 126*8), w128=> Pw(93)(128*8-1 downto 127*8), 
           d_out   => pca_d93_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_94_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(94)(     7 downto    0),   w02 => Pw(94)( 2*8-1 downto    8),   w03 => Pw(94)( 3*8-1 downto  2*8),   w04 => Pw(94)( 4*8-1 downto  3*8),  w05 => Pw(94)( 5*8-1 downto  4*8),   w06 => Pw(94)( 6*8-1 downto  5*8),   w07 => Pw(94)( 7*8-1 downto  6*8),   w08 => Pw(94)( 8*8-1 downto  7*8),  
w09 => Pw(94)( 9*8-1 downto  8*8),   w10 => Pw(94)(10*8-1 downto  9*8),   w11 => Pw(94)(11*8-1 downto 10*8),   w12 => Pw(94)(12*8-1 downto 11*8),   w13 => Pw(94)(13*8-1 downto 12*8),   w14 => Pw(94)(14*8-1 downto 13*8),   w15 => Pw(94)(15*8-1 downto 14*8),   w16 => Pw(94)(16*8-1 downto 15*8),  
w17 => Pw(94)(17*8-1 downto 16*8),   w18 => Pw(94)(18*8-1 downto 17*8),   w19 => Pw(94)(19*8-1 downto 18*8),   w20 => Pw(94)(20*8-1 downto 19*8),   w21 => Pw(94)(21*8-1 downto 20*8),   w22 => Pw(94)(22*8-1 downto 21*8),   w23 => Pw(94)(23*8-1 downto 22*8),   w24 => Pw(94)(24*8-1 downto 23*8),  
w25 => Pw(94)(25*8-1 downto 24*8),   w26 => Pw(94)(26*8-1 downto 25*8),   w27 => Pw(94)(27*8-1 downto 26*8),   w28 => Pw(94)(28*8-1 downto 27*8),   w29 => Pw(94)(29*8-1 downto 28*8),   w30 => Pw(94)(30*8-1 downto 29*8),   w31 => Pw(94)(31*8-1 downto 30*8),   w32 => Pw(94)(32*8-1 downto 31*8),  
w33 => Pw(94)(33*8-1 downto 32*8),   w34 => Pw(94)(34*8-1 downto 33*8),   w35 => Pw(94)(35*8-1 downto 34*8),   w36 => Pw(94)(36*8-1 downto 35*8),   w37 => Pw(94)(37*8-1 downto 36*8),   w38 => Pw(94)(38*8-1 downto 37*8),   w39 => Pw(94)(39*8-1 downto 38*8),   w40 => Pw(94)(40*8-1 downto 39*8),  
w41 => Pw(94)(41*8-1 downto 40*8),   w42 => Pw(94)(42*8-1 downto 41*8),   w43 => Pw(94)(43*8-1 downto 42*8),   w44 => Pw(94)(44*8-1 downto 43*8),   w45 => Pw(94)(45*8-1 downto 44*8),   w46 => Pw(94)(46*8-1 downto 45*8),   w47 => Pw(94)(47*8-1 downto 46*8),   w48 => Pw(94)(48*8-1 downto 47*8),  
w49 => Pw(94)(49*8-1 downto 48*8),   w50 => Pw(94)(50*8-1 downto 49*8),   w51 => Pw(94)(51*8-1 downto 50*8),   w52 => Pw(94)(52*8-1 downto 51*8),   w53 => Pw(94)(53*8-1 downto 52*8),   w54 => Pw(94)(54*8-1 downto 53*8),   w55 => Pw(94)(55*8-1 downto 54*8),   w56 => Pw(94)(56*8-1 downto 55*8),  
w57 => Pw(94)(57*8-1 downto 56*8),   w58 => Pw(94)(58*8-1 downto 57*8),   w59 => Pw(94)(59*8-1 downto 58*8),   w60 => Pw(94)(60*8-1 downto 59*8),   w61 => Pw(94)(61*8-1 downto 60*8),   w62 => Pw(94)(62*8-1 downto 61*8),   w63 => Pw(94)(63*8-1 downto 62*8),   w64 => Pw(94)(64*8-1 downto 63*8), 
w65 => Pw(94)( 65*8-1 downto  64*8), w66 => Pw(94)( 66*8-1 downto  65*8), w67 => Pw(94)( 67*8-1 downto  66*8), w68 => Pw(94)( 68*8-1 downto  67*8), w69 => Pw(94)( 69*8-1 downto  68*8), w70 => Pw(94)( 70*8-1 downto  69*8), w71 => Pw(94)( 71*8-1 downto  70*8), w72 => Pw(94)( 72*8-1 downto  71*8), 
w73 => Pw(94)( 73*8-1 downto  72*8), w74 => Pw(94)( 74*8-1 downto  73*8), w75 => Pw(94)( 75*8-1 downto  74*8), w76 => Pw(94)( 76*8-1 downto  75*8), w77 => Pw(94)( 77*8-1 downto  76*8), w78 => Pw(94)( 78*8-1 downto  77*8), w79 => Pw(94)( 79*8-1 downto  78*8), w80 => Pw(94)( 80*8-1 downto  79*8), 
w81 => Pw(94)( 81*8-1 downto  80*8), w82 => Pw(94)( 82*8-1 downto  81*8), w83 => Pw(94)( 83*8-1 downto  82*8), w84 => Pw(94)( 84*8-1 downto  83*8), w85 => Pw(94)( 85*8-1 downto  84*8), w86 => Pw(94)( 86*8-1 downto  85*8), w87 => Pw(94)( 87*8-1 downto  86*8), w88 => Pw(94)( 88*8-1 downto  87*8), 
w89 => Pw(94)( 89*8-1 downto  88*8), w90 => Pw(94)( 90*8-1 downto  89*8), w91 => Pw(94)( 91*8-1 downto  90*8), w92 => Pw(94)( 92*8-1 downto  91*8), w93 => Pw(94)( 93*8-1 downto  92*8), w94 => Pw(94)( 94*8-1 downto  93*8), w95 => Pw(94)( 95*8-1 downto  94*8), w96 => Pw(94)( 96*8-1 downto  95*8), 
w97 => Pw(94)( 97*8-1 downto  96*8), w98 => Pw(94)( 98*8-1 downto  97*8), w99 => Pw(94)( 99*8-1 downto  98*8), w100=> Pw(94)(100*8-1 downto  99*8), w101=> Pw(94)(101*8-1 downto 100*8), w102=> Pw(94)(102*8-1 downto 101*8), w103=> Pw(94)(103*8-1 downto 102*8), w104=> Pw(94)(104*8-1 downto 103*8), 
w105=> Pw(94)(105*8-1 downto 104*8), w106=> Pw(94)(106*8-1 downto 105*8), w107=> Pw(94)(107*8-1 downto 106*8), w108=> Pw(94)(108*8-1 downto 107*8), w109=> Pw(94)(109*8-1 downto 108*8), w110=> Pw(94)(110*8-1 downto 109*8), w111=> Pw(94)(111*8-1 downto 110*8), w112=> Pw(94)(112*8-1 downto 111*8), 
w113=> Pw(94)(113*8-1 downto 112*8), w114=> Pw(94)(114*8-1 downto 113*8), w115=> Pw(94)(115*8-1 downto 114*8), w116=> Pw(94)(116*8-1 downto 115*8), w117=> Pw(94)(117*8-1 downto 116*8), w118=> Pw(94)(118*8-1 downto 117*8), w119=> Pw(94)(119*8-1 downto 118*8), w120=> Pw(94)(120*8-1 downto 119*8), 
w121=> Pw(94)(121*8-1 downto 120*8), w122=> Pw(94)(122*8-1 downto 121*8), w123=> Pw(94)(123*8-1 downto 122*8), w124=> Pw(94)(124*8-1 downto 123*8), w125=> Pw(94)(125*8-1 downto 124*8), w126=> Pw(94)(126*8-1 downto 125*8), w127=> Pw(94)(127*8-1 downto 126*8), w128=> Pw(94)(128*8-1 downto 127*8), 
           d_out   => pca_d94_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_95_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(95)(     7 downto    0),   w02 => Pw(95)( 2*8-1 downto    8),   w03 => Pw(95)( 3*8-1 downto  2*8),   w04 => Pw(95)( 4*8-1 downto  3*8),   w05 => Pw(95)( 5*8-1 downto  4*8),   w06 => Pw(95)( 6*8-1 downto  5*8),   w07 => Pw(95)( 7*8-1 downto  6*8),   w08 => Pw(95)( 8*8-1 downto  7*8),  
w09 => Pw(95)( 9*8-1 downto  8*8),   w10 => Pw(95)(10*8-1 downto  9*8),   w11 => Pw(95)(11*8-1 downto 10*8),   w12 => Pw(95)(12*8-1 downto 11*8),   w13 => Pw(95)(13*8-1 downto 12*8),   w14 => Pw(95)(14*8-1 downto 13*8),   w15 => Pw(95)(15*8-1 downto 14*8),   w16 => Pw(95)(16*8-1 downto 15*8),  
w17 => Pw(95)(17*8-1 downto 16*8),   w18 => Pw(95)(18*8-1 downto 17*8),   w19 => Pw(95)(19*8-1 downto 18*8),   w20 => Pw(95)(20*8-1 downto 19*8),   w21 => Pw(95)(21*8-1 downto 20*8),   w22 => Pw(95)(22*8-1 downto 21*8),   w23 => Pw(95)(23*8-1 downto 22*8),   w24 => Pw(95)(24*8-1 downto 23*8),  
w25 => Pw(95)(25*8-1 downto 24*8),   w26 => Pw(95)(26*8-1 downto 25*8),   w27 => Pw(95)(27*8-1 downto 26*8),   w28 => Pw(95)(28*8-1 downto 27*8),   w29 => Pw(95)(29*8-1 downto 28*8),   w30 => Pw(95)(30*8-1 downto 29*8),   w31 => Pw(95)(31*8-1 downto 30*8),   w32 => Pw(95)(32*8-1 downto 31*8),  
w33 => Pw(95)(33*8-1 downto 32*8),   w34 => Pw(95)(34*8-1 downto 33*8),   w35 => Pw(95)(35*8-1 downto 34*8),   w36 => Pw(95)(36*8-1 downto 35*8),   w37 => Pw(95)(37*8-1 downto 36*8),   w38 => Pw(95)(38*8-1 downto 37*8),   w39 => Pw(95)(39*8-1 downto 38*8),   w40 => Pw(95)(40*8-1 downto 39*8),  
w41 => Pw(95)(41*8-1 downto 40*8),   w42 => Pw(95)(42*8-1 downto 41*8),   w43 => Pw(95)(43*8-1 downto 42*8),   w44 => Pw(95)(44*8-1 downto 43*8),   w45 => Pw(95)(45*8-1 downto 44*8),   w46 => Pw(95)(46*8-1 downto 45*8),   w47 => Pw(95)(47*8-1 downto 46*8),   w48 => Pw(95)(48*8-1 downto 47*8),  
w49 => Pw(95)(49*8-1 downto 48*8),   w50 => Pw(95)(50*8-1 downto 49*8),   w51 => Pw(95)(51*8-1 downto 50*8),   w52 => Pw(95)(52*8-1 downto 51*8),   w53 => Pw(95)(53*8-1 downto 52*8),   w54 => Pw(95)(54*8-1 downto 53*8),   w55 => Pw(95)(55*8-1 downto 54*8),   w56 => Pw(95)(56*8-1 downto 55*8),  
w57 => Pw(95)(57*8-1 downto 56*8),   w58 => Pw(95)(58*8-1 downto 57*8),   w59 => Pw(95)(59*8-1 downto 58*8),   w60 => Pw(95)(60*8-1 downto 59*8),   w61 => Pw(95)(61*8-1 downto 60*8),   w62 => Pw(95)(62*8-1 downto 61*8),   w63 => Pw(95)(63*8-1 downto 62*8),   w64 => Pw(95)(64*8-1 downto 63*8), 
w65 => Pw(95)( 65*8-1 downto  64*8), w66 => Pw(95)( 66*8-1 downto  65*8), w67 => Pw(95)( 67*8-1 downto  66*8), w68 => Pw(95)( 68*8-1 downto  67*8), w69 => Pw(95)( 69*8-1 downto  68*8), w70 => Pw(95)( 70*8-1 downto  69*8), w71 => Pw(95)( 71*8-1 downto  70*8), w72 => Pw(95)( 72*8-1 downto  71*8), 
w73 => Pw(95)( 73*8-1 downto  72*8), w74 => Pw(95)( 74*8-1 downto  73*8), w75 => Pw(95)( 75*8-1 downto  74*8), w76 => Pw(95)( 76*8-1 downto  75*8), w77 => Pw(95)( 77*8-1 downto  76*8), w78 => Pw(95)( 78*8-1 downto  77*8), w79 => Pw(95)( 79*8-1 downto  78*8), w80 => Pw(95)( 80*8-1 downto  79*8), 
w81 => Pw(95)( 81*8-1 downto  80*8), w82 => Pw(95)( 82*8-1 downto  81*8), w83 => Pw(95)( 83*8-1 downto  82*8), w84 => Pw(95)( 84*8-1 downto  83*8), w85 => Pw(95)( 85*8-1 downto  84*8), w86 => Pw(95)( 86*8-1 downto  85*8), w87 => Pw(95)( 87*8-1 downto  86*8), w88 => Pw(95)( 88*8-1 downto  87*8), 
w89 => Pw(95)( 89*8-1 downto  88*8), w90 => Pw(95)( 90*8-1 downto  89*8), w91 => Pw(95)( 91*8-1 downto  90*8), w92 => Pw(95)( 92*8-1 downto  91*8), w93 => Pw(95)( 93*8-1 downto  92*8), w94 => Pw(95)( 94*8-1 downto  93*8), w95 => Pw(95)( 95*8-1 downto  94*8), w96 => Pw(95)( 96*8-1 downto  95*8), 
w97 => Pw(95)( 97*8-1 downto  96*8), w98 => Pw(95)( 98*8-1 downto  97*8), w99 => Pw(95)( 99*8-1 downto  98*8), w100=> Pw(95)(100*8-1 downto  99*8), w101=> Pw(95)(101*8-1 downto 100*8), w102=> Pw(95)(102*8-1 downto 101*8), w103=> Pw(95)(103*8-1 downto 102*8), w104=> Pw(95)(104*8-1 downto 103*8), 
w105=> Pw(95)(105*8-1 downto 104*8), w106=> Pw(95)(106*8-1 downto 105*8), w107=> Pw(95)(107*8-1 downto 106*8), w108=> Pw(95)(108*8-1 downto 107*8), w109=> Pw(95)(109*8-1 downto 108*8), w110=> Pw(95)(110*8-1 downto 109*8), w111=> Pw(95)(111*8-1 downto 110*8), w112=> Pw(95)(112*8-1 downto 111*8), 
w113=> Pw(95)(113*8-1 downto 112*8), w114=> Pw(95)(114*8-1 downto 113*8), w115=> Pw(95)(115*8-1 downto 114*8), w116=> Pw(95)(116*8-1 downto 115*8), w117=> Pw(95)(117*8-1 downto 116*8), w118=> Pw(95)(118*8-1 downto 117*8), w119=> Pw(95)(119*8-1 downto 118*8), w120=> Pw(95)(120*8-1 downto 119*8), 
w121=> Pw(95)(121*8-1 downto 120*8), w122=> Pw(95)(122*8-1 downto 121*8), w123=> Pw(95)(123*8-1 downto 122*8), w124=> Pw(95)(124*8-1 downto 123*8), w125=> Pw(95)(125*8-1 downto 124*8), w126=> Pw(95)(126*8-1 downto 125*8), w127=> Pw(95)(127*8-1 downto 126*8), w128=> Pw(95)(128*8-1 downto 127*8), 
           d_out   => pca_d95_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_96_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(96)(     7 downto    0),   w02 => Pw(96)( 2*8-1 downto    8),   w03 => Pw(96)( 3*8-1 downto  2*8),   w04 => Pw(96)( 4*8-1 downto  3*8),   w05 => Pw(96)( 5*8-1 downto  4*8),   w06 => Pw(96)( 6*8-1 downto  5*8),   w07 => Pw(96)( 7*8-1 downto  6*8),   w08 => Pw(96)( 8*8-1 downto  7*8),  
w09 => Pw(96)( 9*8-1 downto  8*8),   w10 => Pw(96)(10*8-1 downto  9*8),   w11 => Pw(96)(11*8-1 downto 10*8),   w12 => Pw(96)(12*8-1 downto 11*8),   w13 => Pw(96)(13*8-1 downto 12*8),   w14 => Pw(96)(14*8-1 downto 13*8),   w15 => Pw(96)(15*8-1 downto 14*8),   w16 => Pw(96)(16*8-1 downto 15*8),  
w17 => Pw(96)(17*8-1 downto 16*8),   w18 => Pw(96)(18*8-1 downto 17*8),   w19 => Pw(96)(19*8-1 downto 18*8),   w20 => Pw(96)(20*8-1 downto 19*8),   w21 => Pw(96)(21*8-1 downto 20*8),   w22 => Pw(96)(22*8-1 downto 21*8),   w23 => Pw(96)(23*8-1 downto 22*8),   w24 => Pw(96)(24*8-1 downto 23*8),  
w25 => Pw(96)(25*8-1 downto 24*8),   w26 => Pw(96)(26*8-1 downto 25*8),   w27 => Pw(96)(27*8-1 downto 26*8),   w28 => Pw(96)(28*8-1 downto 27*8),   w29 => Pw(96)(29*8-1 downto 28*8),   w30 => Pw(96)(30*8-1 downto 29*8),   w31 => Pw(96)(31*8-1 downto 30*8),   w32 => Pw(96)(32*8-1 downto 31*8),  
w33 => Pw(96)(33*8-1 downto 32*8),   w34 => Pw(96)(34*8-1 downto 33*8),   w35 => Pw(96)(35*8-1 downto 34*8),   w36 => Pw(96)(36*8-1 downto 35*8),   w37 => Pw(96)(37*8-1 downto 36*8),   w38 => Pw(96)(38*8-1 downto 37*8),   w39 => Pw(96)(39*8-1 downto 38*8),   w40 => Pw(96)(40*8-1 downto 39*8),  
w41 => Pw(96)(41*8-1 downto 40*8),   w42 => Pw(96)(42*8-1 downto 41*8),   w43 => Pw(96)(43*8-1 downto 42*8),   w44 => Pw(96)(44*8-1 downto 43*8),   w45 => Pw(96)(45*8-1 downto 44*8),   w46 => Pw(96)(46*8-1 downto 45*8),   w47 => Pw(96)(47*8-1 downto 46*8),   w48 => Pw(96)(48*8-1 downto 47*8),  
w49 => Pw(96)(49*8-1 downto 48*8),   w50 => Pw(96)(50*8-1 downto 49*8),   w51 => Pw(96)(51*8-1 downto 50*8),   w52 => Pw(96)(52*8-1 downto 51*8),   w53 => Pw(96)(53*8-1 downto 52*8),   w54 => Pw(96)(54*8-1 downto 53*8),   w55 => Pw(96)(55*8-1 downto 54*8),   w56 => Pw(96)(56*8-1 downto 55*8),  
w57 => Pw(96)(57*8-1 downto 56*8),   w58 => Pw(96)(58*8-1 downto 57*8),   w59 => Pw(96)(59*8-1 downto 58*8),   w60 => Pw(96)(60*8-1 downto 59*8),   w61 => Pw(96)(61*8-1 downto 60*8),   w62 => Pw(96)(62*8-1 downto 61*8),   w63 => Pw(96)(63*8-1 downto 62*8),   w64 => Pw(96)(64*8-1 downto 63*8), 
w65 => Pw(96)( 65*8-1 downto  64*8), w66 => Pw(96)( 66*8-1 downto  65*8), w67 => Pw(96)( 67*8-1 downto  66*8), w68 => Pw(96)( 68*8-1 downto  67*8), w69 => Pw(96)( 69*8-1 downto  68*8), w70 => Pw(96)( 70*8-1 downto  69*8), w71 => Pw(96)( 71*8-1 downto  70*8), w72 => Pw(96)( 72*8-1 downto  71*8), 
w73 => Pw(96)( 73*8-1 downto  72*8), w74 => Pw(96)( 74*8-1 downto  73*8), w75 => Pw(96)( 75*8-1 downto  74*8), w76 => Pw(96)( 76*8-1 downto  75*8), w77 => Pw(96)( 77*8-1 downto  76*8), w78 => Pw(96)( 78*8-1 downto  77*8), w79 => Pw(96)( 79*8-1 downto  78*8), w80 => Pw(96)( 80*8-1 downto  79*8), 
w81 => Pw(96)( 81*8-1 downto  80*8), w82 => Pw(96)( 82*8-1 downto  81*8), w83 => Pw(96)( 83*8-1 downto  82*8), w84 => Pw(96)( 84*8-1 downto  83*8), w85 => Pw(96)( 85*8-1 downto  84*8), w86 => Pw(96)( 86*8-1 downto  85*8), w87 => Pw(96)( 87*8-1 downto  86*8), w88 => Pw(96)( 88*8-1 downto  87*8), 
w89 => Pw(96)( 89*8-1 downto  88*8), w90 => Pw(96)( 90*8-1 downto  89*8), w91 => Pw(96)( 91*8-1 downto  90*8), w92 => Pw(96)( 92*8-1 downto  91*8), w93 => Pw(96)( 93*8-1 downto  92*8), w94 => Pw(96)( 94*8-1 downto  93*8), w95 => Pw(96)( 95*8-1 downto  94*8), w96 => Pw(96)( 96*8-1 downto  95*8), 
w97 => Pw(96)( 97*8-1 downto  96*8), w98 => Pw(96)( 98*8-1 downto  97*8), w99 => Pw(96)( 99*8-1 downto  98*8), w100=> Pw(96)(100*8-1 downto  99*8), w101=> Pw(96)(101*8-1 downto 100*8), w102=> Pw(96)(102*8-1 downto 101*8), w103=> Pw(96)(103*8-1 downto 102*8), w104=> Pw(96)(104*8-1 downto 103*8), 
w105=> Pw(96)(105*8-1 downto 104*8), w106=> Pw(96)(106*8-1 downto 105*8), w107=> Pw(96)(107*8-1 downto 106*8), w108=> Pw(96)(108*8-1 downto 107*8), w109=> Pw(96)(109*8-1 downto 108*8), w110=> Pw(96)(110*8-1 downto 109*8), w111=> Pw(96)(111*8-1 downto 110*8), w112=> Pw(96)(112*8-1 downto 111*8), 
w113=> Pw(96)(113*8-1 downto 112*8), w114=> Pw(96)(114*8-1 downto 113*8), w115=> Pw(96)(115*8-1 downto 114*8), w116=> Pw(96)(116*8-1 downto 115*8), w117=> Pw(96)(117*8-1 downto 116*8), w118=> Pw(96)(118*8-1 downto 117*8), w119=> Pw(96)(119*8-1 downto 118*8), w120=> Pw(96)(120*8-1 downto 119*8), 
w121=> Pw(96)(121*8-1 downto 120*8), w122=> Pw(96)(122*8-1 downto 121*8), w123=> Pw(96)(123*8-1 downto 122*8), w124=> Pw(96)(124*8-1 downto 123*8), w125=> Pw(96)(125*8-1 downto 124*8), w126=> Pw(96)(126*8-1 downto 125*8), w127=> Pw(96)(127*8-1 downto 126*8), w128=> Pw(96)(128*8-1 downto 127*8), 
           d_out   => pca_d96_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_97_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(97)(     7 downto    0),   w02 => Pw(97)( 2*8-1 downto    8),   w03 => Pw(97)( 3*8-1 downto  2*8),   w04 => Pw(97)( 4*8-1 downto  3*8),   w05 => Pw(97)( 5*8-1 downto  4*8),   w06 => Pw(97)( 6*8-1 downto  5*8),   w07 => Pw(97)( 7*8-1 downto  6*8),   w08 => Pw(97)( 8*8-1 downto  7*8),  
w09 => Pw(97)( 9*8-1 downto  8*8),   w10 => Pw(97)(10*8-1 downto  9*8),   w11 => Pw(97)(11*8-1 downto 10*8),   w12 => Pw(97)(12*8-1 downto 11*8),   w13 => Pw(97)(13*8-1 downto 12*8),   w14 => Pw(97)(14*8-1 downto 13*8),   w15 => Pw(97)(15*8-1 downto 14*8),   w16 => Pw(97)(16*8-1 downto 15*8),  
w17 => Pw(97)(17*8-1 downto 16*8),   w18 => Pw(97)(18*8-1 downto 17*8),   w19 => Pw(97)(19*8-1 downto 18*8),   w20 => Pw(97)(20*8-1 downto 19*8),   w21 => Pw(97)(21*8-1 downto 20*8),   w22 => Pw(97)(22*8-1 downto 21*8),   w23 => Pw(97)(23*8-1 downto 22*8),   w24 => Pw(97)(24*8-1 downto 23*8),  
w25 => Pw(97)(25*8-1 downto 24*8),   w26 => Pw(97)(26*8-1 downto 25*8),   w27 => Pw(97)(27*8-1 downto 26*8),   w28 => Pw(97)(28*8-1 downto 27*8),   w29 => Pw(97)(29*8-1 downto 28*8),   w30 => Pw(97)(30*8-1 downto 29*8),   w31 => Pw(97)(31*8-1 downto 30*8),   w32 => Pw(97)(32*8-1 downto 31*8),  
w33 => Pw(97)(33*8-1 downto 32*8),   w34 => Pw(97)(34*8-1 downto 33*8),   w35 => Pw(97)(35*8-1 downto 34*8),   w36 => Pw(97)(36*8-1 downto 35*8),   w37 => Pw(97)(37*8-1 downto 36*8),   w38 => Pw(97)(38*8-1 downto 37*8),   w39 => Pw(97)(39*8-1 downto 38*8),   w40 => Pw(97)(40*8-1 downto 39*8),  
w41 => Pw(97)(41*8-1 downto 40*8),   w42 => Pw(97)(42*8-1 downto 41*8),   w43 => Pw(97)(43*8-1 downto 42*8),   w44 => Pw(97)(44*8-1 downto 43*8),   w45 => Pw(97)(45*8-1 downto 44*8),   w46 => Pw(97)(46*8-1 downto 45*8),   w47 => Pw(97)(47*8-1 downto 46*8),   w48 => Pw(97)(48*8-1 downto 47*8),  
w49 => Pw(97)(49*8-1 downto 48*8),   w50 => Pw(97)(50*8-1 downto 49*8),   w51 => Pw(97)(51*8-1 downto 50*8),   w52 => Pw(97)(52*8-1 downto 51*8),   w53 => Pw(97)(53*8-1 downto 52*8),   w54 => Pw(97)(54*8-1 downto 53*8),   w55 => Pw(97)(55*8-1 downto 54*8),   w56 => Pw(97)(56*8-1 downto 55*8),  
w57 => Pw(97)(57*8-1 downto 56*8),   w58 => Pw(97)(58*8-1 downto 57*8),   w59 => Pw(97)(59*8-1 downto 58*8),   w60 => Pw(97)(60*8-1 downto 59*8),   w61 => Pw(97)(61*8-1 downto 60*8),   w62 => Pw(97)(62*8-1 downto 61*8),   w63 => Pw(97)(63*8-1 downto 62*8),   w64 => Pw(97)(64*8-1 downto 63*8), 
w65 => Pw(97)( 65*8-1 downto  64*8), w66 => Pw(97)( 66*8-1 downto  65*8), w67 => Pw(97)( 67*8-1 downto  66*8), w68 => Pw(97)( 68*8-1 downto  67*8), w69 => Pw(97)( 69*8-1 downto  68*8), w70 => Pw(97)( 70*8-1 downto  69*8), w71 => Pw(97)( 71*8-1 downto  70*8), w72 => Pw(97)( 72*8-1 downto  71*8), 
w73 => Pw(97)( 73*8-1 downto  72*8), w74 => Pw(97)( 74*8-1 downto  73*8), w75 => Pw(97)( 75*8-1 downto  74*8), w76 => Pw(97)( 76*8-1 downto  75*8), w77 => Pw(97)( 77*8-1 downto  76*8), w78 => Pw(97)( 78*8-1 downto  77*8), w79 => Pw(97)( 79*8-1 downto  78*8), w80 => Pw(97)( 80*8-1 downto  79*8), 
w81 => Pw(97)( 81*8-1 downto  80*8), w82 => Pw(97)( 82*8-1 downto  81*8), w83 => Pw(97)( 83*8-1 downto  82*8), w84 => Pw(97)( 84*8-1 downto  83*8), w85 => Pw(97)( 85*8-1 downto  84*8), w86 => Pw(97)( 86*8-1 downto  85*8), w87 => Pw(97)( 87*8-1 downto  86*8), w88 => Pw(97)( 88*8-1 downto  87*8), 
w89 => Pw(97)( 89*8-1 downto  88*8), w90 => Pw(97)( 90*8-1 downto  89*8), w91 => Pw(97)( 91*8-1 downto  90*8), w92 => Pw(97)( 92*8-1 downto  91*8), w93 => Pw(97)( 93*8-1 downto  92*8), w94 => Pw(97)( 94*8-1 downto  93*8), w95 => Pw(97)( 95*8-1 downto  94*8), w96 => Pw(97)( 96*8-1 downto  95*8), 
w97 => Pw(97)( 97*8-1 downto  96*8), w98 => Pw(97)( 98*8-1 downto  97*8), w99 => Pw(97)( 99*8-1 downto  98*8), w100=> Pw(97)(100*8-1 downto  99*8), w101=> Pw(97)(101*8-1 downto 100*8), w102=> Pw(97)(102*8-1 downto 101*8), w103=> Pw(97)(103*8-1 downto 102*8), w104=> Pw(97)(104*8-1 downto 103*8), 
w105=> Pw(97)(105*8-1 downto 104*8), w106=> Pw(97)(106*8-1 downto 105*8), w107=> Pw(97)(107*8-1 downto 106*8), w108=> Pw(97)(108*8-1 downto 107*8), w109=> Pw(97)(109*8-1 downto 108*8), w110=> Pw(97)(110*8-1 downto 109*8), w111=> Pw(97)(111*8-1 downto 110*8), w112=> Pw(97)(112*8-1 downto 111*8), 
w113=> Pw(97)(113*8-1 downto 112*8), w114=> Pw(97)(114*8-1 downto 113*8), w115=> Pw(97)(115*8-1 downto 114*8), w116=> Pw(97)(116*8-1 downto 115*8), w117=> Pw(97)(117*8-1 downto 116*8), w118=> Pw(97)(118*8-1 downto 117*8), w119=> Pw(97)(119*8-1 downto 118*8), w120=> Pw(97)(120*8-1 downto 119*8), 
w121=> Pw(97)(121*8-1 downto 120*8), w122=> Pw(97)(122*8-1 downto 121*8), w123=> Pw(97)(123*8-1 downto 122*8), w124=> Pw(97)(124*8-1 downto 123*8), w125=> Pw(97)(125*8-1 downto 124*8), w126=> Pw(97)(126*8-1 downto 125*8), w127=> Pw(97)(127*8-1 downto 126*8), w128=> Pw(97)(128*8-1 downto 127*8), 
           d_out   => pca_d97_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_98_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(98)(     7 downto    0),   w02 => Pw(98)( 2*8-1 downto    8),   w03 => Pw(98)( 3*8-1 downto  2*8),   w04 => Pw(98)( 4*8-1 downto  3*8),   w05 => Pw(98)( 5*8-1 downto  4*8),   w06 => Pw(98)( 6*8-1 downto  5*8),   w07 => Pw(98)( 7*8-1 downto  6*8),   w08 => Pw(98)( 8*8-1 downto  7*8),  
w09 => Pw(98)( 9*8-1 downto  8*8),   w10 => Pw(98)(10*8-1 downto  9*8),   w11 => Pw(98)(11*8-1 downto 10*8),   w12 => Pw(98)(12*8-1 downto 11*8),   w13 => Pw(98)(13*8-1 downto 12*8),   w14 => Pw(98)(14*8-1 downto 13*8),   w15 => Pw(98)(15*8-1 downto 14*8),   w16 => Pw(98)(16*8-1 downto 15*8),  
w17 => Pw(98)(17*8-1 downto 16*8),   w18 => Pw(98)(18*8-1 downto 17*8),   w19 => Pw(98)(19*8-1 downto 18*8),   w20 => Pw(98)(20*8-1 downto 19*8),   w21 => Pw(98)(21*8-1 downto 20*8),   w22 => Pw(98)(22*8-1 downto 21*8),   w23 => Pw(98)(23*8-1 downto 22*8),   w24 => Pw(98)(24*8-1 downto 23*8),  
w25 => Pw(98)(25*8-1 downto 24*8),   w26 => Pw(98)(26*8-1 downto 25*8),   w27 => Pw(98)(27*8-1 downto 26*8),   w28 => Pw(98)(28*8-1 downto 27*8),   w29 => Pw(98)(29*8-1 downto 28*8),   w30 => Pw(98)(30*8-1 downto 29*8),   w31 => Pw(98)(31*8-1 downto 30*8),   w32 => Pw(98)(32*8-1 downto 31*8),  
w33 => Pw(98)(33*8-1 downto 32*8),   w34 => Pw(98)(34*8-1 downto 33*8),   w35 => Pw(98)(35*8-1 downto 34*8),   w36 => Pw(98)(36*8-1 downto 35*8),   w37 => Pw(98)(37*8-1 downto 36*8),   w38 => Pw(98)(38*8-1 downto 37*8),   w39 => Pw(98)(39*8-1 downto 38*8),   w40 => Pw(98)(40*8-1 downto 39*8),  
w41 => Pw(98)(41*8-1 downto 40*8),   w42 => Pw(98)(42*8-1 downto 41*8),   w43 => Pw(98)(43*8-1 downto 42*8),   w44 => Pw(98)(44*8-1 downto 43*8),   w45 => Pw(98)(45*8-1 downto 44*8),   w46 => Pw(98)(46*8-1 downto 45*8),   w47 => Pw(98)(47*8-1 downto 46*8),   w48 => Pw(98)(48*8-1 downto 47*8),  
w49 => Pw(98)(49*8-1 downto 48*8),   w50 => Pw(98)(50*8-1 downto 49*8),   w51 => Pw(98)(51*8-1 downto 50*8),   w52 => Pw(98)(52*8-1 downto 51*8),   w53 => Pw(98)(53*8-1 downto 52*8),   w54 => Pw(98)(54*8-1 downto 53*8),   w55 => Pw(98)(55*8-1 downto 54*8),   w56 => Pw(98)(56*8-1 downto 55*8),  
w57 => Pw(98)(57*8-1 downto 56*8),   w58 => Pw(98)(58*8-1 downto 57*8),   w59 => Pw(98)(59*8-1 downto 58*8),   w60 => Pw(98)(60*8-1 downto 59*8),   w61 => Pw(98)(61*8-1 downto 60*8),   w62 => Pw(98)(62*8-1 downto 61*8),   w63 => Pw(98)(63*8-1 downto 62*8),   w64 => Pw(98)(64*8-1 downto 63*8), 
w65 => Pw(98)( 65*8-1 downto  64*8), w66 => Pw(98)( 66*8-1 downto  65*8), w67 => Pw(98)( 67*8-1 downto  66*8), w68 => Pw(98)( 68*8-1 downto  67*8), w69 => Pw(98)( 69*8-1 downto  68*8), w70 => Pw(98)( 70*8-1 downto  69*8), w71 => Pw(98)( 71*8-1 downto  70*8), w72 => Pw(98)( 72*8-1 downto  71*8), 
w73 => Pw(98)( 73*8-1 downto  72*8), w74 => Pw(98)( 74*8-1 downto  73*8), w75 => Pw(98)( 75*8-1 downto  74*8), w76 => Pw(98)( 76*8-1 downto  75*8), w77 => Pw(98)( 77*8-1 downto  76*8), w78 => Pw(98)( 78*8-1 downto  77*8), w79 => Pw(98)( 79*8-1 downto  78*8), w80 => Pw(98)( 80*8-1 downto  79*8), 
w81 => Pw(98)( 81*8-1 downto  80*8), w82 => Pw(98)( 82*8-1 downto  81*8), w83 => Pw(98)( 83*8-1 downto  82*8), w84 => Pw(98)( 84*8-1 downto  83*8), w85 => Pw(98)( 85*8-1 downto  84*8), w86 => Pw(98)( 86*8-1 downto  85*8), w87 => Pw(98)( 87*8-1 downto  86*8), w88 => Pw(98)( 88*8-1 downto  87*8), 
w89 => Pw(98)( 89*8-1 downto  88*8), w90 => Pw(98)( 90*8-1 downto  89*8), w91 => Pw(98)( 91*8-1 downto  90*8), w92 => Pw(98)( 92*8-1 downto  91*8), w93 => Pw(98)( 93*8-1 downto  92*8), w94 => Pw(98)( 94*8-1 downto  93*8), w95 => Pw(98)( 95*8-1 downto  94*8), w96 => Pw(98)( 96*8-1 downto  95*8), 
w97 => Pw(98)( 97*8-1 downto  96*8), w98 => Pw(98)( 98*8-1 downto  97*8), w99 => Pw(98)( 99*8-1 downto  98*8), w100=> Pw(98)(100*8-1 downto  99*8), w101=> Pw(98)(101*8-1 downto 100*8), w102=> Pw(98)(102*8-1 downto 101*8), w103=> Pw(98)(103*8-1 downto 102*8), w104=> Pw(98)(104*8-1 downto 103*8), 
w105=> Pw(98)(105*8-1 downto 104*8), w106=> Pw(98)(106*8-1 downto 105*8), w107=> Pw(98)(107*8-1 downto 106*8), w108=> Pw(98)(108*8-1 downto 107*8), w109=> Pw(98)(109*8-1 downto 108*8), w110=> Pw(98)(110*8-1 downto 109*8), w111=> Pw(98)(111*8-1 downto 110*8), w112=> Pw(98)(112*8-1 downto 111*8), 
w113=> Pw(98)(113*8-1 downto 112*8), w114=> Pw(98)(114*8-1 downto 113*8), w115=> Pw(98)(115*8-1 downto 114*8), w116=> Pw(98)(116*8-1 downto 115*8), w117=> Pw(98)(117*8-1 downto 116*8), w118=> Pw(98)(118*8-1 downto 117*8), w119=> Pw(98)(119*8-1 downto 118*8), w120=> Pw(98)(120*8-1 downto 119*8), 
w121=> Pw(98)(121*8-1 downto 120*8), w122=> Pw(98)(122*8-1 downto 121*8), w123=> Pw(98)(123*8-1 downto 122*8), w124=> Pw(98)(124*8-1 downto 123*8), w125=> Pw(98)(125*8-1 downto 124*8), w126=> Pw(98)(126*8-1 downto 125*8), w127=> Pw(98)(127*8-1 downto 126*8), w128=> Pw(98)(128*8-1 downto 127*8), 
           d_out   => pca_d98_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_99_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(99)(     7 downto    0),   w02 => Pw(99)( 2*8-1 downto    8),   w03 => Pw(99)( 3*8-1 downto  2*8),   w04 => Pw(99)( 4*8-1 downto  3*8),   w05 => Pw(99)( 5*8-1 downto  4*8),   w06 => Pw(99)( 6*8-1 downto  5*8),   w07 => Pw(99)( 7*8-1 downto  6*8),   w08 => Pw(99)( 8*8-1 downto  7*8),  
w09 => Pw(99)( 9*8-1 downto  8*8),   w10 => Pw(99)(10*8-1 downto  9*8),   w11 => Pw(99)(11*8-1 downto 10*8),   w12 => Pw(99)(12*8-1 downto 11*8),   w13 => Pw(99)(13*8-1 downto 12*8),   w14 => Pw(99)(14*8-1 downto 13*8),   w15 => Pw(99)(15*8-1 downto 14*8),   w16 => Pw(99)(16*8-1 downto 15*8),  
w17 => Pw(99)(17*8-1 downto 16*8),   w18 => Pw(99)(18*8-1 downto 17*8),   w19 => Pw(99)(19*8-1 downto 18*8),   w20 => Pw(99)(20*8-1 downto 19*8),   w21 => Pw(99)(21*8-1 downto 20*8),   w22 => Pw(99)(22*8-1 downto 21*8),   w23 => Pw(99)(23*8-1 downto 22*8),   w24 => Pw(99)(24*8-1 downto 23*8),  
w25 => Pw(99)(25*8-1 downto 24*8),   w26 => Pw(99)(26*8-1 downto 25*8),   w27 => Pw(99)(27*8-1 downto 26*8),   w28 => Pw(99)(28*8-1 downto 27*8),   w29 => Pw(99)(29*8-1 downto 28*8),   w30 => Pw(99)(30*8-1 downto 29*8),   w31 => Pw(99)(31*8-1 downto 30*8),   w32 => Pw(99)(32*8-1 downto 31*8),  
w33 => Pw(99)(33*8-1 downto 32*8),   w34 => Pw(99)(34*8-1 downto 33*8),   w35 => Pw(99)(35*8-1 downto 34*8),   w36 => Pw(99)(36*8-1 downto 35*8),   w37 => Pw(99)(37*8-1 downto 36*8),   w38 => Pw(99)(38*8-1 downto 37*8),   w39 => Pw(99)(39*8-1 downto 38*8),   w40 => Pw(99)(40*8-1 downto 39*8),  
w41 => Pw(99)(41*8-1 downto 40*8),   w42 => Pw(99)(42*8-1 downto 41*8),   w43 => Pw(99)(43*8-1 downto 42*8),   w44 => Pw(99)(44*8-1 downto 43*8),   w45 => Pw(99)(45*8-1 downto 44*8),   w46 => Pw(99)(46*8-1 downto 45*8),   w47 => Pw(99)(47*8-1 downto 46*8),   w48 => Pw(99)(48*8-1 downto 47*8),  
w49 => Pw(99)(49*8-1 downto 48*8),   w50 => Pw(99)(50*8-1 downto 49*8),   w51 => Pw(99)(51*8-1 downto 50*8),   w52 => Pw(99)(52*8-1 downto 51*8),   w53 => Pw(99)(53*8-1 downto 52*8),   w54 => Pw(99)(54*8-1 downto 53*8),   w55 => Pw(99)(55*8-1 downto 54*8),   w56 => Pw(99)(56*8-1 downto 55*8),  
w57 => Pw(99)(57*8-1 downto 56*8),   w58 => Pw(99)(58*8-1 downto 57*8),   w59 => Pw(99)(59*8-1 downto 58*8),   w60 => Pw(99)(60*8-1 downto 59*8),   w61 => Pw(99)(61*8-1 downto 60*8),   w62 => Pw(99)(62*8-1 downto 61*8),   w63 => Pw(99)(63*8-1 downto 62*8),   w64 => Pw(99)(64*8-1 downto 63*8), 
w65 => Pw(99)( 65*8-1 downto  64*8), w66 => Pw(99)( 66*8-1 downto  65*8), w67 => Pw(99)( 67*8-1 downto  66*8), w68 => Pw(99)( 68*8-1 downto  67*8), w69 => Pw(99)( 69*8-1 downto  68*8), w70 => Pw(99)( 70*8-1 downto  69*8), w71 => Pw(99)( 71*8-1 downto  70*8), w72 => Pw(99)( 72*8-1 downto  71*8), 
w73 => Pw(99)( 73*8-1 downto  72*8), w74 => Pw(99)( 74*8-1 downto  73*8), w75 => Pw(99)( 75*8-1 downto  74*8), w76 => Pw(99)( 76*8-1 downto  75*8), w77 => Pw(99)( 77*8-1 downto  76*8), w78 => Pw(99)( 78*8-1 downto  77*8), w79 => Pw(99)( 79*8-1 downto  78*8), w80 => Pw(99)( 80*8-1 downto  79*8), 
w81 => Pw(99)( 81*8-1 downto  80*8), w82 => Pw(99)( 82*8-1 downto  81*8), w83 => Pw(99)( 83*8-1 downto  82*8), w84 => Pw(99)( 84*8-1 downto  83*8), w85 => Pw(99)( 85*8-1 downto  84*8), w86 => Pw(99)( 86*8-1 downto  85*8), w87 => Pw(99)( 87*8-1 downto  86*8), w88 => Pw(99)( 88*8-1 downto  87*8), 
w89 => Pw(99)( 89*8-1 downto  88*8), w90 => Pw(99)( 90*8-1 downto  89*8), w91 => Pw(99)( 91*8-1 downto  90*8), w92 => Pw(99)( 92*8-1 downto  91*8), w93 => Pw(99)( 93*8-1 downto  92*8), w94 => Pw(99)( 94*8-1 downto  93*8), w95 => Pw(99)( 95*8-1 downto  94*8), w96 => Pw(99)( 96*8-1 downto  95*8), 
w97 => Pw(99)( 97*8-1 downto  96*8), w98 => Pw(99)( 98*8-1 downto  97*8), w99 => Pw(99)( 99*8-1 downto  98*8), w100=> Pw(99)(100*8-1 downto  99*8), w101=> Pw(99)(101*8-1 downto 100*8), w102=> Pw(99)(102*8-1 downto 101*8), w103=> Pw(99)(103*8-1 downto 102*8), w104=> Pw(99)(104*8-1 downto 103*8), 
w105=> Pw(99)(105*8-1 downto 104*8), w106=> Pw(99)(106*8-1 downto 105*8), w107=> Pw(99)(107*8-1 downto 106*8), w108=> Pw(99)(108*8-1 downto 107*8), w109=> Pw(99)(109*8-1 downto 108*8), w110=> Pw(99)(110*8-1 downto 109*8), w111=> Pw(99)(111*8-1 downto 110*8), w112=> Pw(99)(112*8-1 downto 111*8), 
w113=> Pw(99)(113*8-1 downto 112*8), w114=> Pw(99)(114*8-1 downto 113*8), w115=> Pw(99)(115*8-1 downto 114*8), w116=> Pw(99)(116*8-1 downto 115*8), w117=> Pw(99)(117*8-1 downto 116*8), w118=> Pw(99)(118*8-1 downto 117*8), w119=> Pw(99)(119*8-1 downto 118*8), w120=> Pw(99)(120*8-1 downto 119*8), 
w121=> Pw(99)(121*8-1 downto 120*8), w122=> Pw(99)(122*8-1 downto 121*8), w123=> Pw(99)(123*8-1 downto 122*8), w124=> Pw(99)(124*8-1 downto 123*8), w125=> Pw(99)(125*8-1 downto 124*8), w126=> Pw(99)(126*8-1 downto 125*8), w127=> Pw(99)(127*8-1 downto 126*8), w128=> Pw(99)(128*8-1 downto 127*8), 
           d_out   => pca_d99_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_100_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(100)(     7 downto    0),   w02 => Pw(100)( 2*8-1 downto    8),   w03 => Pw(100)( 3*8-1 downto  2*8),   w04 => Pw(100)( 4*8-1 downto  3*8),   w05 => Pw(100)( 5*8-1 downto  4*8),   w06 => Pw(100)( 6*8-1 downto  5*8),   w07 => Pw(100)( 7*8-1 downto  6*8),   w08 => Pw(100)( 8*8-1 downto  7*8),  
w09 => Pw(100)( 9*8-1 downto  8*8),   w10 => Pw(100)(10*8-1 downto  9*8),   w11 => Pw(100)(11*8-1 downto 10*8),   w12 => Pw(100)(12*8-1 downto 11*8),   w13 => Pw(100)(13*8-1 downto 12*8),   w14 => Pw(100)(14*8-1 downto 13*8),   w15 => Pw(100)(15*8-1 downto 14*8),   w16 => Pw(100)(16*8-1 downto 15*8),  
w17 => Pw(100)(17*8-1 downto 16*8),   w18 => Pw(100)(18*8-1 downto 17*8),   w19 => Pw(100)(19*8-1 downto 18*8),   w20 => Pw(100)(20*8-1 downto 19*8),   w21 => Pw(100)(21*8-1 downto 20*8),   w22 => Pw(100)(22*8-1 downto 21*8),   w23 => Pw(100)(23*8-1 downto 22*8),   w24 => Pw(100)(24*8-1 downto 23*8),  
w25 => Pw(100)(25*8-1 downto 24*8),   w26 => Pw(100)(26*8-1 downto 25*8),   w27 => Pw(100)(27*8-1 downto 26*8),   w28 => Pw(100)(28*8-1 downto 27*8),   w29 => Pw(100)(29*8-1 downto 28*8),   w30 => Pw(100)(30*8-1 downto 29*8),   w31 => Pw(100)(31*8-1 downto 30*8),   w32 => Pw(100)(32*8-1 downto 31*8),  
w33 => Pw(100)(33*8-1 downto 32*8),   w34 => Pw(100)(34*8-1 downto 33*8),   w35 => Pw(100)(35*8-1 downto 34*8),   w36 => Pw(100)(36*8-1 downto 35*8),   w37 => Pw(100)(37*8-1 downto 36*8),   w38 => Pw(100)(38*8-1 downto 37*8),   w39 => Pw(100)(39*8-1 downto 38*8),   w40 => Pw(100)(40*8-1 downto 39*8),  
w41 => Pw(100)(41*8-1 downto 40*8),   w42 => Pw(100)(42*8-1 downto 41*8),   w43 => Pw(100)(43*8-1 downto 42*8),   w44 => Pw(100)(44*8-1 downto 43*8),   w45 => Pw(100)(45*8-1 downto 44*8),   w46 => Pw(100)(46*8-1 downto 45*8),   w47 => Pw(100)(47*8-1 downto 46*8),   w48 => Pw(100)(48*8-1 downto 47*8),  
w49 => Pw(100)(49*8-1 downto 48*8),   w50 => Pw(100)(50*8-1 downto 49*8),   w51 => Pw(100)(51*8-1 downto 50*8),   w52 => Pw(100)(52*8-1 downto 51*8),   w53 => Pw(100)(53*8-1 downto 52*8),   w54 => Pw(100)(54*8-1 downto 53*8),   w55 => Pw(100)(55*8-1 downto 54*8),   w56 => Pw(100)(56*8-1 downto 55*8),  
w57 => Pw(100)(57*8-1 downto 56*8),   w58 => Pw(100)(58*8-1 downto 57*8),   w59 => Pw(100)(59*8-1 downto 58*8),   w60 => Pw(100)(60*8-1 downto 59*8),   w61 => Pw(100)(61*8-1 downto 60*8),   w62 => Pw(100)(62*8-1 downto 61*8),   w63 => Pw(100)(63*8-1 downto 62*8),   w64 => Pw(100)(64*8-1 downto 63*8), 
w65 => Pw(100)( 65*8-1 downto  64*8), w66 => Pw(100)( 66*8-1 downto  65*8), w67 => Pw(100)( 67*8-1 downto  66*8), w68 => Pw(100)( 68*8-1 downto  67*8), w69 => Pw(100)( 69*8-1 downto  68*8), w70 => Pw(100)( 70*8-1 downto  69*8), w71 => Pw(100)( 71*8-1 downto  70*8), w72 => Pw(100)( 72*8-1 downto  71*8), 
w73 => Pw(100)( 73*8-1 downto  72*8), w74 => Pw(100)( 74*8-1 downto  73*8), w75 => Pw(100)( 75*8-1 downto  74*8), w76 => Pw(100)( 76*8-1 downto  75*8), w77 => Pw(100)( 77*8-1 downto  76*8), w78 => Pw(100)( 78*8-1 downto  77*8), w79 => Pw(100)( 79*8-1 downto  78*8), w80 => Pw(100)( 80*8-1 downto  79*8), 
w81 => Pw(100)( 81*8-1 downto  80*8), w82 => Pw(100)( 82*8-1 downto  81*8), w83 => Pw(100)( 83*8-1 downto  82*8), w84 => Pw(100)( 84*8-1 downto  83*8), w85 => Pw(100)( 85*8-1 downto  84*8), w86 => Pw(100)( 86*8-1 downto  85*8), w87 => Pw(100)( 87*8-1 downto  86*8), w88 => Pw(100)( 88*8-1 downto  87*8), 
w89 => Pw(100)( 89*8-1 downto  88*8), w90 => Pw(100)( 90*8-1 downto  89*8), w91 => Pw(100)( 91*8-1 downto  90*8), w92 => Pw(100)( 92*8-1 downto  91*8), w93 => Pw(100)( 93*8-1 downto  92*8), w94 => Pw(100)( 94*8-1 downto  93*8), w95 => Pw(100)( 95*8-1 downto  94*8), w96 => Pw(100)( 96*8-1 downto  95*8), 
w97 => Pw(100)( 97*8-1 downto  96*8), w98 => Pw(100)( 98*8-1 downto  97*8), w99 => Pw(100)( 99*8-1 downto  98*8), w100=> Pw(100)(100*8-1 downto  99*8), w101=> Pw(100)(101*8-1 downto 100*8), w102=> Pw(100)(102*8-1 downto 101*8), w103=> Pw(100)(103*8-1 downto 102*8), w104=> Pw(100)(104*8-1 downto 103*8), 
w105=> Pw(100)(105*8-1 downto 104*8), w106=> Pw(100)(106*8-1 downto 105*8), w107=> Pw(100)(107*8-1 downto 106*8), w108=> Pw(100)(108*8-1 downto 107*8), w109=> Pw(100)(109*8-1 downto 108*8), w110=> Pw(100)(110*8-1 downto 109*8), w111=> Pw(100)(111*8-1 downto 110*8), w112=> Pw(100)(112*8-1 downto 111*8), 
w113=> Pw(100)(113*8-1 downto 112*8), w114=> Pw(100)(114*8-1 downto 113*8), w115=> Pw(100)(115*8-1 downto 114*8), w116=> Pw(100)(116*8-1 downto 115*8), w117=> Pw(100)(117*8-1 downto 116*8), w118=> Pw(100)(118*8-1 downto 117*8), w119=> Pw(100)(119*8-1 downto 118*8), w120=> Pw(100)(120*8-1 downto 119*8), 
w121=> Pw(100)(121*8-1 downto 120*8), w122=> Pw(100)(122*8-1 downto 121*8), w123=> Pw(100)(123*8-1 downto 122*8), w124=> Pw(100)(124*8-1 downto 123*8), w125=> Pw(100)(125*8-1 downto 124*8), w126=> Pw(100)(126*8-1 downto 125*8), w127=> Pw(100)(127*8-1 downto 126*8), w128=> Pw(100)(128*8-1 downto 127*8), 
           d_out   => pca_d100_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_101_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(101)(     7 downto    0),   w02 => Pw(101)( 2*8-1 downto    8),   w03 => Pw(101)( 3*8-1 downto  2*8),   w04 => Pw(101)( 4*8-1 downto  3*8),   w05 => Pw(101)( 5*8-1 downto  4*8),   w06 => Pw(101)( 6*8-1 downto  5*8),   w07 => Pw(101)( 7*8-1 downto  6*8),   w08 => Pw(101)( 8*8-1 downto  7*8),  
w09 => Pw(101)( 9*8-1 downto  8*8),   w10 => Pw(101)(10*8-1 downto  9*8),   w11 => Pw(101)(11*8-1 downto 10*8),   w12 => Pw(101)(12*8-1 downto 11*8),   w13 => Pw(101)(13*8-1 downto 12*8),   w14 => Pw(101)(14*8-1 downto 13*8),   w15 => Pw(101)(15*8-1 downto 14*8),   w16 => Pw(101)(16*8-1 downto 15*8),  
w17 => Pw(101)(17*8-1 downto 16*8),   w18 => Pw(101)(18*8-1 downto 17*8),   w19 => Pw(101)(19*8-1 downto 18*8),   w20 => Pw(101)(20*8-1 downto 19*8),   w21 => Pw(101)(21*8-1 downto 20*8),   w22 => Pw(101)(22*8-1 downto 21*8),   w23 => Pw(101)(23*8-1 downto 22*8),   w24 => Pw(101)(24*8-1 downto 23*8),  
w25 => Pw(101)(25*8-1 downto 24*8),   w26 => Pw(101)(26*8-1 downto 25*8),   w27 => Pw(101)(27*8-1 downto 26*8),   w28 => Pw(101)(28*8-1 downto 27*8),   w29 => Pw(101)(29*8-1 downto 28*8),   w30 => Pw(101)(30*8-1 downto 29*8),   w31 => Pw(101)(31*8-1 downto 30*8),   w32 => Pw(101)(32*8-1 downto 31*8),  
w33 => Pw(101)(33*8-1 downto 32*8),   w34 => Pw(101)(34*8-1 downto 33*8),   w35 => Pw(101)(35*8-1 downto 34*8),   w36 => Pw(101)(36*8-1 downto 35*8),   w37 => Pw(101)(37*8-1 downto 36*8),   w38 => Pw(101)(38*8-1 downto 37*8),   w39 => Pw(101)(39*8-1 downto 38*8),   w40 => Pw(101)(40*8-1 downto 39*8),  
w41 => Pw(101)(41*8-1 downto 40*8),   w42 => Pw(101)(42*8-1 downto 41*8),   w43 => Pw(101)(43*8-1 downto 42*8),   w44 => Pw(101)(44*8-1 downto 43*8),   w45 => Pw(101)(45*8-1 downto 44*8),   w46 => Pw(101)(46*8-1 downto 45*8),   w47 => Pw(101)(47*8-1 downto 46*8),   w48 => Pw(101)(48*8-1 downto 47*8),  
w49 => Pw(101)(49*8-1 downto 48*8),   w50 => Pw(101)(50*8-1 downto 49*8),   w51 => Pw(101)(51*8-1 downto 50*8),   w52 => Pw(101)(52*8-1 downto 51*8),   w53 => Pw(101)(53*8-1 downto 52*8),   w54 => Pw(101)(54*8-1 downto 53*8),   w55 => Pw(101)(55*8-1 downto 54*8),   w56 => Pw(101)(56*8-1 downto 55*8),  
w57 => Pw(101)(57*8-1 downto 56*8),   w58 => Pw(101)(58*8-1 downto 57*8),   w59 => Pw(101)(59*8-1 downto 58*8),   w60 => Pw(101)(60*8-1 downto 59*8),   w61 => Pw(101)(61*8-1 downto 60*8),   w62 => Pw(101)(62*8-1 downto 61*8),   w63 => Pw(101)(63*8-1 downto 62*8),   w64 => Pw(101)(64*8-1 downto 63*8), 
w65 => Pw(101)( 65*8-1 downto  64*8), w66 => Pw(101)( 66*8-1 downto  65*8), w67 => Pw(101)( 67*8-1 downto  66*8), w68 => Pw(101)( 68*8-1 downto  67*8), w69 => Pw(101)( 69*8-1 downto  68*8), w70 => Pw(101)( 70*8-1 downto  69*8), w71 => Pw(101)( 71*8-1 downto  70*8), w72 => Pw(101)( 72*8-1 downto  71*8), 
w73 => Pw(101)( 73*8-1 downto  72*8), w74 => Pw(101)( 74*8-1 downto  73*8), w75 => Pw(101)( 75*8-1 downto  74*8), w76 => Pw(101)( 76*8-1 downto  75*8), w77 => Pw(101)( 77*8-1 downto  76*8), w78 => Pw(101)( 78*8-1 downto  77*8), w79 => Pw(101)( 79*8-1 downto  78*8), w80 => Pw(101)( 80*8-1 downto  79*8), 
w81 => Pw(101)( 81*8-1 downto  80*8), w82 => Pw(101)( 82*8-1 downto  81*8), w83 => Pw(101)( 83*8-1 downto  82*8), w84 => Pw(101)( 84*8-1 downto  83*8), w85 => Pw(101)( 85*8-1 downto  84*8), w86 => Pw(101)( 86*8-1 downto  85*8), w87 => Pw(101)( 87*8-1 downto  86*8), w88 => Pw(101)( 88*8-1 downto  87*8), 
w89 => Pw(101)( 89*8-1 downto  88*8), w90 => Pw(101)( 90*8-1 downto  89*8), w91 => Pw(101)( 91*8-1 downto  90*8), w92 => Pw(101)( 92*8-1 downto  91*8), w93 => Pw(101)( 93*8-1 downto  92*8), w94 => Pw(101)( 94*8-1 downto  93*8), w95 => Pw(101)( 95*8-1 downto  94*8), w96 => Pw(101)( 96*8-1 downto  95*8), 
w97 => Pw(101)( 97*8-1 downto  96*8), w98 => Pw(101)( 98*8-1 downto  97*8), w99 => Pw(101)( 99*8-1 downto  98*8), w100=> Pw(101)(100*8-1 downto  99*8), w101=> Pw(101)(101*8-1 downto 100*8), w102=> Pw(101)(102*8-1 downto 101*8), w103=> Pw(101)(103*8-1 downto 102*8), w104=> Pw(101)(104*8-1 downto 103*8), 
w105=> Pw(101)(105*8-1 downto 104*8), w106=> Pw(101)(106*8-1 downto 105*8), w107=> Pw(101)(107*8-1 downto 106*8), w108=> Pw(101)(108*8-1 downto 107*8), w109=> Pw(101)(109*8-1 downto 108*8), w110=> Pw(101)(110*8-1 downto 109*8), w111=> Pw(101)(111*8-1 downto 110*8), w112=> Pw(101)(112*8-1 downto 111*8), 
w113=> Pw(101)(113*8-1 downto 112*8), w114=> Pw(101)(114*8-1 downto 113*8), w115=> Pw(101)(115*8-1 downto 114*8), w116=> Pw(101)(116*8-1 downto 115*8), w117=> Pw(101)(117*8-1 downto 116*8), w118=> Pw(101)(118*8-1 downto 117*8), w119=> Pw(101)(119*8-1 downto 118*8), w120=> Pw(101)(120*8-1 downto 119*8), 
w121=> Pw(101)(121*8-1 downto 120*8), w122=> Pw(101)(122*8-1 downto 121*8), w123=> Pw(101)(123*8-1 downto 122*8), w124=> Pw(101)(124*8-1 downto 123*8), w125=> Pw(101)(125*8-1 downto 124*8), w126=> Pw(101)(126*8-1 downto 125*8), w127=> Pw(101)(127*8-1 downto 126*8), w128=> Pw(101)(128*8-1 downto 127*8), 
           d_out   => pca_d101_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_102_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(102)(     7 downto    0),   w02 => Pw(102)( 2*8-1 downto    8),   w03 => Pw(102)( 3*8-1 downto  2*8),   w04 => Pw(102)( 4*8-1 downto  3*8),   w05 => Pw(102)( 5*8-1 downto  4*8),   w06 => Pw(102)( 6*8-1 downto  5*8),   w07 => Pw(102)( 7*8-1 downto  6*8),   w08 => Pw(102)( 8*8-1 downto  7*8),  
w09 => Pw(102)( 9*8-1 downto  8*8),   w10 => Pw(102)(10*8-1 downto  9*8),   w11 => Pw(102)(11*8-1 downto 10*8),   w12 => Pw(102)(12*8-1 downto 11*8),   w13 => Pw(102)(13*8-1 downto 12*8),   w14 => Pw(102)(14*8-1 downto 13*8),   w15 => Pw(102)(15*8-1 downto 14*8),   w16 => Pw(102)(16*8-1 downto 15*8),  
w17 => Pw(102)(17*8-1 downto 16*8),   w18 => Pw(102)(18*8-1 downto 17*8),   w19 => Pw(102)(19*8-1 downto 18*8),   w20 => Pw(102)(20*8-1 downto 19*8),   w21 => Pw(102)(21*8-1 downto 20*8),   w22 => Pw(102)(22*8-1 downto 21*8),   w23 => Pw(102)(23*8-1 downto 22*8),   w24 => Pw(102)(24*8-1 downto 23*8),  
w25 => Pw(102)(25*8-1 downto 24*8),   w26 => Pw(102)(26*8-1 downto 25*8),   w27 => Pw(102)(27*8-1 downto 26*8),   w28 => Pw(102)(28*8-1 downto 27*8),   w29 => Pw(102)(29*8-1 downto 28*8),   w30 => Pw(102)(30*8-1 downto 29*8),   w31 => Pw(102)(31*8-1 downto 30*8),   w32 => Pw(102)(32*8-1 downto 31*8),  
w33 => Pw(102)(33*8-1 downto 32*8),   w34 => Pw(102)(34*8-1 downto 33*8),   w35 => Pw(102)(35*8-1 downto 34*8),   w36 => Pw(102)(36*8-1 downto 35*8),   w37 => Pw(102)(37*8-1 downto 36*8),   w38 => Pw(102)(38*8-1 downto 37*8),   w39 => Pw(102)(39*8-1 downto 38*8),   w40 => Pw(102)(40*8-1 downto 39*8),  
w41 => Pw(102)(41*8-1 downto 40*8),   w42 => Pw(102)(42*8-1 downto 41*8),   w43 => Pw(102)(43*8-1 downto 42*8),   w44 => Pw(102)(44*8-1 downto 43*8),   w45 => Pw(102)(45*8-1 downto 44*8),   w46 => Pw(102)(46*8-1 downto 45*8),   w47 => Pw(102)(47*8-1 downto 46*8),   w48 => Pw(102)(48*8-1 downto 47*8),  
w49 => Pw(102)(49*8-1 downto 48*8),   w50 => Pw(102)(50*8-1 downto 49*8),   w51 => Pw(102)(51*8-1 downto 50*8),   w52 => Pw(102)(52*8-1 downto 51*8),   w53 => Pw(102)(53*8-1 downto 52*8),   w54 => Pw(102)(54*8-1 downto 53*8),   w55 => Pw(102)(55*8-1 downto 54*8),   w56 => Pw(102)(56*8-1 downto 55*8),  
w57 => Pw(102)(57*8-1 downto 56*8),   w58 => Pw(102)(58*8-1 downto 57*8),   w59 => Pw(102)(59*8-1 downto 58*8),   w60 => Pw(102)(60*8-1 downto 59*8),   w61 => Pw(102)(61*8-1 downto 60*8),   w62 => Pw(102)(62*8-1 downto 61*8),   w63 => Pw(102)(63*8-1 downto 62*8),   w64 => Pw(102)(64*8-1 downto 63*8), 
w65 => Pw(102)( 65*8-1 downto  64*8), w66 => Pw(102)( 66*8-1 downto  65*8), w67 => Pw(102)( 67*8-1 downto  66*8), w68 => Pw(102)( 68*8-1 downto  67*8), w69 => Pw(102)( 69*8-1 downto  68*8), w70 => Pw(102)( 70*8-1 downto  69*8), w71 => Pw(102)( 71*8-1 downto  70*8), w72 => Pw(102)( 72*8-1 downto  71*8), 
w73 => Pw(102)( 73*8-1 downto  72*8), w74 => Pw(102)( 74*8-1 downto  73*8), w75 => Pw(102)( 75*8-1 downto  74*8), w76 => Pw(102)( 76*8-1 downto  75*8), w77 => Pw(102)( 77*8-1 downto  76*8), w78 => Pw(102)( 78*8-1 downto  77*8), w79 => Pw(102)( 79*8-1 downto  78*8), w80 => Pw(102)( 80*8-1 downto  79*8), 
w81 => Pw(102)( 81*8-1 downto  80*8), w82 => Pw(102)( 82*8-1 downto  81*8), w83 => Pw(102)( 83*8-1 downto  82*8), w84 => Pw(102)( 84*8-1 downto  83*8), w85 => Pw(102)( 85*8-1 downto  84*8), w86 => Pw(102)( 86*8-1 downto  85*8), w87 => Pw(102)( 87*8-1 downto  86*8), w88 => Pw(102)( 88*8-1 downto  87*8), 
w89 => Pw(102)( 89*8-1 downto  88*8), w90 => Pw(102)( 90*8-1 downto  89*8), w91 => Pw(102)( 91*8-1 downto  90*8), w92 => Pw(102)( 92*8-1 downto  91*8), w93 => Pw(102)( 93*8-1 downto  92*8), w94 => Pw(102)( 94*8-1 downto  93*8), w95 => Pw(102)( 95*8-1 downto  94*8), w96 => Pw(102)( 96*8-1 downto  95*8), 
w97 => Pw(102)( 97*8-1 downto  96*8), w98 => Pw(102)( 98*8-1 downto  97*8), w99 => Pw(102)( 99*8-1 downto  98*8), w100=> Pw(102)(100*8-1 downto  99*8), w101=> Pw(102)(101*8-1 downto 100*8), w102=> Pw(102)(102*8-1 downto 101*8), w103=> Pw(102)(103*8-1 downto 102*8), w104=> Pw(102)(104*8-1 downto 103*8), 
w105=> Pw(102)(105*8-1 downto 104*8), w106=> Pw(102)(106*8-1 downto 105*8), w107=> Pw(102)(107*8-1 downto 106*8), w108=> Pw(102)(108*8-1 downto 107*8), w109=> Pw(102)(109*8-1 downto 108*8), w110=> Pw(102)(110*8-1 downto 109*8), w111=> Pw(102)(111*8-1 downto 110*8), w112=> Pw(102)(112*8-1 downto 111*8), 
w113=> Pw(102)(113*8-1 downto 112*8), w114=> Pw(102)(114*8-1 downto 113*8), w115=> Pw(102)(115*8-1 downto 114*8), w116=> Pw(102)(116*8-1 downto 115*8), w117=> Pw(102)(117*8-1 downto 116*8), w118=> Pw(102)(118*8-1 downto 117*8), w119=> Pw(102)(119*8-1 downto 118*8), w120=> Pw(102)(120*8-1 downto 119*8), 
w121=> Pw(102)(121*8-1 downto 120*8), w122=> Pw(102)(122*8-1 downto 121*8), w123=> Pw(102)(123*8-1 downto 122*8), w124=> Pw(102)(124*8-1 downto 123*8), w125=> Pw(102)(125*8-1 downto 124*8), w126=> Pw(102)(126*8-1 downto 125*8), w127=> Pw(102)(127*8-1 downto 126*8), w128=> Pw(102)(128*8-1 downto 127*8), 
           d_out   => pca_d102_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_103_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(103)(     7 downto    0),   w02 => Pw(103)( 2*8-1 downto    8),   w03 => Pw(103)( 3*8-1 downto  2*8),   w04 => Pw(103)( 4*8-1 downto  3*8),  w05 => Pw(103)( 5*8-1 downto  4*8),   w06 => Pw(103)( 6*8-1 downto  5*8),   w07 => Pw(103)( 7*8-1 downto  6*8),   w08 => Pw(103)( 8*8-1 downto  7*8),  
w09 => Pw(103)( 9*8-1 downto  8*8),   w10 => Pw(103)(10*8-1 downto  9*8),   w11 => Pw(103)(11*8-1 downto 10*8),   w12 => Pw(103)(12*8-1 downto 11*8),  w13 => Pw(103)(13*8-1 downto 12*8),   w14 => Pw(103)(14*8-1 downto 13*8),   w15 => Pw(103)(15*8-1 downto 14*8),   w16 => Pw(103)(16*8-1 downto 15*8),  
w17 => Pw(103)(17*8-1 downto 16*8),   w18 => Pw(103)(18*8-1 downto 17*8),   w19 => Pw(103)(19*8-1 downto 18*8),   w20 => Pw(103)(20*8-1 downto 19*8),  w21 => Pw(103)(21*8-1 downto 20*8),   w22 => Pw(103)(22*8-1 downto 21*8),   w23 => Pw(103)(23*8-1 downto 22*8),   w24 => Pw(103)(24*8-1 downto 23*8),  
w25 => Pw(103)(25*8-1 downto 24*8),   w26 => Pw(103)(26*8-1 downto 25*8),   w27 => Pw(103)(27*8-1 downto 26*8),   w28 => Pw(103)(28*8-1 downto 27*8),  w29 => Pw(103)(29*8-1 downto 28*8),   w30 => Pw(103)(30*8-1 downto 29*8),   w31 => Pw(103)(31*8-1 downto 30*8),   w32 => Pw(103)(32*8-1 downto 31*8),  
w33 => Pw(103)(33*8-1 downto 32*8),   w34 => Pw(103)(34*8-1 downto 33*8),   w35 => Pw(103)(35*8-1 downto 34*8),   w36 => Pw(103)(36*8-1 downto 35*8),   w37 => Pw(103)(37*8-1 downto 36*8),   w38 => Pw(103)(38*8-1 downto 37*8),   w39 => Pw(103)(39*8-1 downto 38*8),   w40 => Pw(103)(40*8-1 downto 39*8),  
w41 => Pw(103)(41*8-1 downto 40*8),   w42 => Pw(103)(42*8-1 downto 41*8),   w43 => Pw(103)(43*8-1 downto 42*8),   w44 => Pw(103)(44*8-1 downto 43*8),   w45 => Pw(103)(45*8-1 downto 44*8),   w46 => Pw(103)(46*8-1 downto 45*8),   w47 => Pw(103)(47*8-1 downto 46*8),   w48 => Pw(103)(48*8-1 downto 47*8),  
w49 => Pw(103)(49*8-1 downto 48*8),   w50 => Pw(103)(50*8-1 downto 49*8),   w51 => Pw(103)(51*8-1 downto 50*8),   w52 => Pw(103)(52*8-1 downto 51*8),   w53 => Pw(103)(53*8-1 downto 52*8),   w54 => Pw(103)(54*8-1 downto 53*8),   w55 => Pw(103)(55*8-1 downto 54*8),   w56 => Pw(103)(56*8-1 downto 55*8),  
w57 => Pw(103)(57*8-1 downto 56*8),   w58 => Pw(103)(58*8-1 downto 57*8),   w59 => Pw(103)(59*8-1 downto 58*8),   w60 => Pw(103)(60*8-1 downto 59*8),   w61 => Pw(103)(61*8-1 downto 60*8),   w62 => Pw(103)(62*8-1 downto 61*8),   w63 => Pw(103)(63*8-1 downto 62*8),   w64 => Pw(103)(64*8-1 downto 63*8), 
w65 => Pw(103)( 65*8-1 downto  64*8), w66 => Pw(103)( 66*8-1 downto  65*8), w67 => Pw(103)( 67*8-1 downto  66*8), w68 => Pw(103)( 68*8-1 downto  67*8), w69 => Pw(103)( 69*8-1 downto  68*8), w70 => Pw(103)( 70*8-1 downto  69*8), w71 => Pw(103)( 71*8-1 downto  70*8), w72 => Pw(103)( 72*8-1 downto  71*8), 
w73 => Pw(103)( 73*8-1 downto  72*8), w74 => Pw(103)( 74*8-1 downto  73*8), w75 => Pw(103)( 75*8-1 downto  74*8), w76 => Pw(103)( 76*8-1 downto  75*8), w77 => Pw(103)( 77*8-1 downto  76*8), w78 => Pw(103)( 78*8-1 downto  77*8), w79 => Pw(103)( 79*8-1 downto  78*8), w80 => Pw(103)( 80*8-1 downto  79*8), 
w81 => Pw(103)( 81*8-1 downto  80*8), w82 => Pw(103)( 82*8-1 downto  81*8), w83 => Pw(103)( 83*8-1 downto  82*8), w84 => Pw(103)( 84*8-1 downto  83*8), w85 => Pw(103)( 85*8-1 downto  84*8), w86 => Pw(103)( 86*8-1 downto  85*8), w87 => Pw(103)( 87*8-1 downto  86*8), w88 => Pw(103)( 88*8-1 downto  87*8), 
w89 => Pw(103)( 89*8-1 downto  88*8), w90 => Pw(103)( 90*8-1 downto  89*8), w91 => Pw(103)( 91*8-1 downto  90*8), w92 => Pw(103)( 92*8-1 downto  91*8), w93 => Pw(103)( 93*8-1 downto  92*8), w94 => Pw(103)( 94*8-1 downto  93*8), w95 => Pw(103)( 95*8-1 downto  94*8), w96 => Pw(103)( 96*8-1 downto  95*8), 
w97 => Pw(103)( 97*8-1 downto  96*8), w98 => Pw(103)( 98*8-1 downto  97*8), w99 => Pw(103)( 99*8-1 downto  98*8), w100=> Pw(103)(100*8-1 downto  99*8), w101=> Pw(103)(101*8-1 downto 100*8), w102=> Pw(103)(102*8-1 downto 101*8), w103=> Pw(103)(103*8-1 downto 102*8), w104=> Pw(103)(104*8-1 downto 103*8), 
w105=> Pw(103)(105*8-1 downto 104*8), w106=> Pw(103)(106*8-1 downto 105*8), w107=> Pw(103)(107*8-1 downto 106*8), w108=> Pw(103)(108*8-1 downto 107*8), w109=> Pw(103)(109*8-1 downto 108*8), w110=> Pw(103)(110*8-1 downto 109*8), w111=> Pw(103)(111*8-1 downto 110*8), w112=> Pw(103)(112*8-1 downto 111*8), 
w113=> Pw(103)(113*8-1 downto 112*8), w114=> Pw(103)(114*8-1 downto 113*8), w115=> Pw(103)(115*8-1 downto 114*8), w116=> Pw(103)(116*8-1 downto 115*8), w117=> Pw(103)(117*8-1 downto 116*8), w118=> Pw(103)(118*8-1 downto 117*8), w119=> Pw(103)(119*8-1 downto 118*8), w120=> Pw(103)(120*8-1 downto 119*8), 
w121=> Pw(103)(121*8-1 downto 120*8), w122=> Pw(103)(122*8-1 downto 121*8), w123=> Pw(103)(123*8-1 downto 122*8), w124=> Pw(103)(124*8-1 downto 123*8), w125=> Pw(103)(125*8-1 downto 124*8), w126=> Pw(103)(126*8-1 downto 125*8), w127=> Pw(103)(127*8-1 downto 126*8), w128=> Pw(103)(128*8-1 downto 127*8), 
           d_out   => pca_d103_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_104_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(104)(     7 downto    0),   w02 => Pw(104)( 2*8-1 downto    8),   w03 => Pw(104)( 3*8-1 downto  2*8),   w04 => Pw(104)( 4*8-1 downto  3*8),   
w05 => Pw(104)( 5*8-1 downto  4*8),   w06 => Pw(104)( 6*8-1 downto  5*8),   w07 => Pw(104)( 7*8-1 downto  6*8),   w08 => Pw(104)( 8*8-1 downto  7*8),  
w09 => Pw(104)( 9*8-1 downto  8*8),   w10 => Pw(104)(10*8-1 downto  9*8),   w11 => Pw(104)(11*8-1 downto 10*8),   w12 => Pw(104)(12*8-1 downto 11*8),   
w13 => Pw(104)(13*8-1 downto 12*8),   w14 => Pw(104)(14*8-1 downto 13*8),   w15 => Pw(104)(15*8-1 downto 14*8),   w16 => Pw(104)(16*8-1 downto 15*8),  
w17 => Pw(104)(17*8-1 downto 16*8),   w18 => Pw(104)(18*8-1 downto 17*8),   w19 => Pw(104)(19*8-1 downto 18*8),   w20 => Pw(104)(20*8-1 downto 19*8),   
w21 => Pw(104)(21*8-1 downto 20*8),   w22 => Pw(104)(22*8-1 downto 21*8),   w23 => Pw(104)(23*8-1 downto 22*8),   w24 => Pw(104)(24*8-1 downto 23*8),  
w25 => Pw(104)(25*8-1 downto 24*8),   w26 => Pw(104)(26*8-1 downto 25*8),   w27 => Pw(104)(27*8-1 downto 26*8),   w28 => Pw(104)(28*8-1 downto 27*8),   
w29 => Pw(104)(29*8-1 downto 28*8),   w30 => Pw(104)(30*8-1 downto 29*8),   w31 => Pw(104)(31*8-1 downto 30*8),   w32 => Pw(104)(32*8-1 downto 31*8),  
w33 => Pw(104)(33*8-1 downto 32*8),   w34 => Pw(104)(34*8-1 downto 33*8),   w35 => Pw(104)(35*8-1 downto 34*8),   w36 => Pw(104)(36*8-1 downto 35*8),   
w37 => Pw(104)(37*8-1 downto 36*8),   w38 => Pw(104)(38*8-1 downto 37*8),   w39 => Pw(104)(39*8-1 downto 38*8),   w40 => Pw(104)(40*8-1 downto 39*8),  
w41 => Pw(104)(41*8-1 downto 40*8),   w42 => Pw(104)(42*8-1 downto 41*8),   w43 => Pw(104)(43*8-1 downto 42*8),   w44 => Pw(104)(44*8-1 downto 43*8),   
w45 => Pw(104)(45*8-1 downto 44*8),   w46 => Pw(104)(46*8-1 downto 45*8),   w47 => Pw(104)(47*8-1 downto 46*8),   w48 => Pw(104)(48*8-1 downto 47*8),  
w49 => Pw(104)(49*8-1 downto 48*8),   w50 => Pw(104)(50*8-1 downto 49*8),   w51 => Pw(104)(51*8-1 downto 50*8),   w52 => Pw(104)(52*8-1 downto 51*8),   
w53 => Pw(104)(53*8-1 downto 52*8),   w54 => Pw(104)(54*8-1 downto 53*8),   w55 => Pw(104)(55*8-1 downto 54*8),   w56 => Pw(104)(56*8-1 downto 55*8),  
w57 => Pw(104)(57*8-1 downto 56*8),   w58 => Pw(104)(58*8-1 downto 57*8),   w59 => Pw(104)(59*8-1 downto 58*8),   w60 => Pw(104)(60*8-1 downto 59*8),   
w61 => Pw(104)(61*8-1 downto 60*8),   w62 => Pw(104)(62*8-1 downto 61*8),   w63 => Pw(104)(63*8-1 downto 62*8),   w64 => Pw(104)(64*8-1 downto 63*8), 
w65 => Pw(104)( 65*8-1 downto  64*8), w66 => Pw(104)( 66*8-1 downto  65*8), w67 => Pw(104)( 67*8-1 downto  66*8), w68 => Pw(104)( 68*8-1 downto  67*8), 
w69 => Pw(104)( 69*8-1 downto  68*8), w70 => Pw(104)( 70*8-1 downto  69*8), w71 => Pw(104)( 71*8-1 downto  70*8), w72 => Pw(104)( 72*8-1 downto  71*8), 
w73 => Pw(104)( 73*8-1 downto  72*8), w74 => Pw(104)( 74*8-1 downto  73*8), w75 => Pw(104)( 75*8-1 downto  74*8), w76 => Pw(104)( 76*8-1 downto  75*8), 
w77 => Pw(104)( 77*8-1 downto  76*8), w78 => Pw(104)( 78*8-1 downto  77*8), w79 => Pw(104)( 79*8-1 downto  78*8), w80 => Pw(104)( 80*8-1 downto  79*8), 
w81 => Pw(104)( 81*8-1 downto  80*8), w82 => Pw(104)( 82*8-1 downto  81*8), w83 => Pw(104)( 83*8-1 downto  82*8), w84 => Pw(104)( 84*8-1 downto  83*8), 
w85 => Pw(104)( 85*8-1 downto  84*8), w86 => Pw(104)( 86*8-1 downto  85*8), w87 => Pw(104)( 87*8-1 downto  86*8), w88 => Pw(104)( 88*8-1 downto  87*8), 
w89 => Pw(104)( 89*8-1 downto  88*8), w90 => Pw(104)( 90*8-1 downto  89*8), w91 => Pw(104)( 91*8-1 downto  90*8), w92 => Pw(104)( 92*8-1 downto  91*8), 
w93 => Pw(104)( 93*8-1 downto  92*8), w94 => Pw(104)( 94*8-1 downto  93*8), w95 => Pw(104)( 95*8-1 downto  94*8), w96 => Pw(104)( 96*8-1 downto  95*8), 
w97 => Pw(104)( 97*8-1 downto  96*8), w98 => Pw(104)( 98*8-1 downto  97*8), w99 => Pw(104)( 99*8-1 downto  98*8), w100=> Pw(104)(100*8-1 downto  99*8), 
w101=> Pw(104)(101*8-1 downto 100*8), w102=> Pw(104)(102*8-1 downto 101*8), w103=> Pw(104)(103*8-1 downto 102*8), w104=> Pw(104)(104*8-1 downto 103*8), 
w105=> Pw(104)(105*8-1 downto 104*8), w106=> Pw(104)(106*8-1 downto 105*8), w107=> Pw(104)(107*8-1 downto 106*8), w108=> Pw(104)(108*8-1 downto 107*8), 
w109=> Pw(104)(109*8-1 downto 108*8), w110=> Pw(104)(110*8-1 downto 109*8), w111=> Pw(104)(111*8-1 downto 110*8), w112=> Pw(104)(112*8-1 downto 111*8), 
w113=> Pw(104)(113*8-1 downto 112*8), w114=> Pw(104)(114*8-1 downto 113*8), w115=> Pw(104)(115*8-1 downto 114*8), w116=> Pw(104)(116*8-1 downto 115*8), 
w117=> Pw(104)(117*8-1 downto 116*8), w118=> Pw(104)(118*8-1 downto 117*8), w119=> Pw(104)(119*8-1 downto 118*8), w120=> Pw(104)(120*8-1 downto 119*8), 
w121=> Pw(104)(121*8-1 downto 120*8), w122=> Pw(104)(122*8-1 downto 121*8), w123=> Pw(104)(123*8-1 downto 122*8), w124=> Pw(104)(124*8-1 downto 123*8), 
w125=> Pw(104)(125*8-1 downto 124*8), w126=> Pw(104)(126*8-1 downto 125*8), w127=> Pw(104)(127*8-1 downto 126*8), w128=> Pw(104)(128*8-1 downto 127*8), 
           d_out   => pca_d104_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_105_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(105)(     7 downto    0),   w02 => Pw(105)( 2*8-1 downto    8),   w03 => Pw(105)( 3*8-1 downto  2*8),   w04 => Pw(105)( 4*8-1 downto  3*8),   
w05 => Pw(105)( 5*8-1 downto  4*8),   w06 => Pw(105)( 6*8-1 downto  5*8),   w07 => Pw(105)( 7*8-1 downto  6*8),   w08 => Pw(105)( 8*8-1 downto  7*8),  
w09 => Pw(105)( 9*8-1 downto  8*8),   w10 => Pw(105)(10*8-1 downto  9*8),   w11 => Pw(105)(11*8-1 downto 10*8),   w12 => Pw(105)(12*8-1 downto 11*8),   
w13 => Pw(105)(13*8-1 downto 12*8),   w14 => Pw(105)(14*8-1 downto 13*8),   w15 => Pw(105)(15*8-1 downto 14*8),   w16 => Pw(105)(16*8-1 downto 15*8),  
w17 => Pw(105)(17*8-1 downto 16*8),   w18 => Pw(105)(18*8-1 downto 17*8),   w19 => Pw(105)(19*8-1 downto 18*8),   w20 => Pw(105)(20*8-1 downto 19*8),   
w21 => Pw(105)(21*8-1 downto 20*8),   w22 => Pw(105)(22*8-1 downto 21*8),   w23 => Pw(105)(23*8-1 downto 22*8),   w24 => Pw(105)(24*8-1 downto 23*8),  
w25 => Pw(105)(25*8-1 downto 24*8),   w26 => Pw(105)(26*8-1 downto 25*8),   w27 => Pw(105)(27*8-1 downto 26*8),   w28 => Pw(105)(28*8-1 downto 27*8),   
w29 => Pw(105)(29*8-1 downto 28*8),   w30 => Pw(105)(30*8-1 downto 29*8),   w31 => Pw(105)(31*8-1 downto 30*8),   w32 => Pw(105)(32*8-1 downto 31*8),  
w33 => Pw(105)(33*8-1 downto 32*8),   w34 => Pw(105)(34*8-1 downto 33*8),   w35 => Pw(105)(35*8-1 downto 34*8),   w36 => Pw(105)(36*8-1 downto 35*8),   
w37 => Pw(105)(37*8-1 downto 36*8),   w38 => Pw(105)(38*8-1 downto 37*8),   w39 => Pw(105)(39*8-1 downto 38*8),   w40 => Pw(105)(40*8-1 downto 39*8),  
w41 => Pw(105)(41*8-1 downto 40*8),   w42 => Pw(105)(42*8-1 downto 41*8),   w43 => Pw(105)(43*8-1 downto 42*8),   w44 => Pw(105)(44*8-1 downto 43*8),   
w45 => Pw(105)(45*8-1 downto 44*8),   w46 => Pw(105)(46*8-1 downto 45*8),   w47 => Pw(105)(47*8-1 downto 46*8),   w48 => Pw(105)(48*8-1 downto 47*8),  
w49 => Pw(105)(49*8-1 downto 48*8),   w50 => Pw(105)(50*8-1 downto 49*8),   w51 => Pw(105)(51*8-1 downto 50*8),   w52 => Pw(105)(52*8-1 downto 51*8),   
w53 => Pw(105)(53*8-1 downto 52*8),   w54 => Pw(105)(54*8-1 downto 53*8),   w55 => Pw(105)(55*8-1 downto 54*8),   w56 => Pw(105)(56*8-1 downto 55*8),  
w57 => Pw(105)(57*8-1 downto 56*8),   w58 => Pw(105)(58*8-1 downto 57*8),   w59 => Pw(105)(59*8-1 downto 58*8),   w60 => Pw(105)(60*8-1 downto 59*8),   
w61 => Pw(105)(61*8-1 downto 60*8),   w62 => Pw(105)(62*8-1 downto 61*8),   w63 => Pw(105)(63*8-1 downto 62*8),   w64 => Pw(105)(64*8-1 downto 63*8), 
w65 => Pw(105)( 65*8-1 downto  64*8), w66 => Pw(105)( 66*8-1 downto  65*8), w67 => Pw(105)( 67*8-1 downto  66*8), w68 => Pw(105)( 68*8-1 downto  67*8), 
w69 => Pw(105)( 69*8-1 downto  68*8), w70 => Pw(105)( 70*8-1 downto  69*8), w71 => Pw(105)( 71*8-1 downto  70*8), w72 => Pw(105)( 72*8-1 downto  71*8), 
w73 => Pw(105)( 73*8-1 downto  72*8), w74 => Pw(105)( 74*8-1 downto  73*8), w75 => Pw(105)( 75*8-1 downto  74*8), w76 => Pw(105)( 76*8-1 downto  75*8), 
w77 => Pw(105)( 77*8-1 downto  76*8), w78 => Pw(105)( 78*8-1 downto  77*8), w79 => Pw(105)( 79*8-1 downto  78*8), w80 => Pw(105)( 80*8-1 downto  79*8), 
w81 => Pw(105)( 81*8-1 downto  80*8), w82 => Pw(105)( 82*8-1 downto  81*8), w83 => Pw(105)( 83*8-1 downto  82*8), w84 => Pw(105)( 84*8-1 downto  83*8), 
w85 => Pw(105)( 85*8-1 downto  84*8), w86 => Pw(105)( 86*8-1 downto  85*8), w87 => Pw(105)( 87*8-1 downto  86*8), w88 => Pw(105)( 88*8-1 downto  87*8), 
w89 => Pw(105)( 89*8-1 downto  88*8), w90 => Pw(105)( 90*8-1 downto  89*8), w91 => Pw(105)( 91*8-1 downto  90*8), w92 => Pw(105)( 92*8-1 downto  91*8), 
w93 => Pw(105)( 93*8-1 downto  92*8), w94 => Pw(105)( 94*8-1 downto  93*8), w95 => Pw(105)( 95*8-1 downto  94*8), w96 => Pw(105)( 96*8-1 downto  95*8), 
w97 => Pw(105)( 97*8-1 downto  96*8), w98 => Pw(105)( 98*8-1 downto  97*8), w99 => Pw(105)( 99*8-1 downto  98*8), w100=> Pw(105)(100*8-1 downto  99*8), 
w101=> Pw(105)(101*8-1 downto 100*8), w102=> Pw(105)(102*8-1 downto 101*8), w103=> Pw(105)(103*8-1 downto 102*8), w104=> Pw(105)(104*8-1 downto 103*8), 
w105=> Pw(105)(105*8-1 downto 104*8), w106=> Pw(105)(106*8-1 downto 105*8), w107=> Pw(105)(107*8-1 downto 106*8), w108=> Pw(105)(108*8-1 downto 107*8), 
w109=> Pw(105)(109*8-1 downto 108*8), w110=> Pw(105)(110*8-1 downto 109*8), w111=> Pw(105)(111*8-1 downto 110*8), w112=> Pw(105)(112*8-1 downto 111*8), 
w113=> Pw(105)(113*8-1 downto 112*8), w114=> Pw(105)(114*8-1 downto 113*8), w115=> Pw(105)(115*8-1 downto 114*8), w116=> Pw(105)(116*8-1 downto 115*8), 
w117=> Pw(105)(117*8-1 downto 116*8), w118=> Pw(105)(118*8-1 downto 117*8), w119=> Pw(105)(119*8-1 downto 118*8), w120=> Pw(105)(120*8-1 downto 119*8), 
w121=> Pw(105)(121*8-1 downto 120*8), w122=> Pw(105)(122*8-1 downto 121*8), w123=> Pw(105)(123*8-1 downto 122*8), w124=> Pw(105)(124*8-1 downto 123*8), 
w125=> Pw(105)(125*8-1 downto 124*8), w126=> Pw(105)(126*8-1 downto 125*8), w127=> Pw(105)(127*8-1 downto 126*8), w128=> Pw(105)(128*8-1 downto 127*8), 
           d_out   => pca_d105_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_106_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(106)(     7 downto    0),   w02 => Pw(106)( 2*8-1 downto    8),   w03 => Pw(106)( 3*8-1 downto  2*8),   w04 => Pw(106)( 4*8-1 downto  3*8),   
w05 => Pw(106)( 5*8-1 downto  4*8),   w06 => Pw(106)( 6*8-1 downto  5*8),   w07 => Pw(106)( 7*8-1 downto  6*8),   w08 => Pw(106)( 8*8-1 downto  7*8),  
w09 => Pw(106)( 9*8-1 downto  8*8),   w10 => Pw(106)(10*8-1 downto  9*8),   w11 => Pw(106)(11*8-1 downto 10*8),   w12 => Pw(106)(12*8-1 downto 11*8),   
w13 => Pw(106)(13*8-1 downto 12*8),   w14 => Pw(106)(14*8-1 downto 13*8),   w15 => Pw(106)(15*8-1 downto 14*8),   w16 => Pw(106)(16*8-1 downto 15*8),  
w17 => Pw(106)(17*8-1 downto 16*8),   w18 => Pw(106)(18*8-1 downto 17*8),   w19 => Pw(106)(19*8-1 downto 18*8),   w20 => Pw(106)(20*8-1 downto 19*8),   
w21 => Pw(106)(21*8-1 downto 20*8),   w22 => Pw(106)(22*8-1 downto 21*8),   w23 => Pw(106)(23*8-1 downto 22*8),   w24 => Pw(106)(24*8-1 downto 23*8),  
w25 => Pw(106)(25*8-1 downto 24*8),   w26 => Pw(106)(26*8-1 downto 25*8),   w27 => Pw(106)(27*8-1 downto 26*8),   w28 => Pw(106)(28*8-1 downto 27*8),   
w29 => Pw(106)(29*8-1 downto 28*8),   w30 => Pw(106)(30*8-1 downto 29*8),   w31 => Pw(106)(31*8-1 downto 30*8),   w32 => Pw(106)(32*8-1 downto 31*8),  
w33 => Pw(106)(33*8-1 downto 32*8),   w34 => Pw(106)(34*8-1 downto 33*8),   w35 => Pw(106)(35*8-1 downto 34*8),   w36 => Pw(106)(36*8-1 downto 35*8),   
w37 => Pw(106)(37*8-1 downto 36*8),   w38 => Pw(106)(38*8-1 downto 37*8),   w39 => Pw(106)(39*8-1 downto 38*8),   w40 => Pw(106)(40*8-1 downto 39*8),  
w41 => Pw(106)(41*8-1 downto 40*8),   w42 => Pw(106)(42*8-1 downto 41*8),   w43 => Pw(106)(43*8-1 downto 42*8),   w44 => Pw(106)(44*8-1 downto 43*8),   
w45 => Pw(106)(45*8-1 downto 44*8),   w46 => Pw(106)(46*8-1 downto 45*8),   w47 => Pw(106)(47*8-1 downto 46*8),   w48 => Pw(106)(48*8-1 downto 47*8),  
w49 => Pw(106)(49*8-1 downto 48*8),   w50 => Pw(106)(50*8-1 downto 49*8),   w51 => Pw(106)(51*8-1 downto 50*8),   w52 => Pw(106)(52*8-1 downto 51*8),   
w53 => Pw(106)(53*8-1 downto 52*8),   w54 => Pw(106)(54*8-1 downto 53*8),   w55 => Pw(106)(55*8-1 downto 54*8),   w56 => Pw(106)(56*8-1 downto 55*8),  
w57 => Pw(106)(57*8-1 downto 56*8),   w58 => Pw(106)(58*8-1 downto 57*8),   w59 => Pw(106)(59*8-1 downto 58*8),   w60 => Pw(106)(60*8-1 downto 59*8),   
w61 => Pw(106)(61*8-1 downto 60*8),   w62 => Pw(106)(62*8-1 downto 61*8),   w63 => Pw(106)(63*8-1 downto 62*8),   w64 => Pw(106)(64*8-1 downto 63*8), 
w65 => Pw(106)( 65*8-1 downto  64*8), w66 => Pw(106)( 66*8-1 downto  65*8), w67 => Pw(106)( 67*8-1 downto  66*8), w68 => Pw(106)( 68*8-1 downto  67*8), 
w69 => Pw(106)( 69*8-1 downto  68*8), w70 => Pw(106)( 70*8-1 downto  69*8), w71 => Pw(106)( 71*8-1 downto  70*8), w72 => Pw(106)( 72*8-1 downto  71*8), 
w73 => Pw(106)( 73*8-1 downto  72*8), w74 => Pw(106)( 74*8-1 downto  73*8), w75 => Pw(106)( 75*8-1 downto  74*8), w76 => Pw(106)( 76*8-1 downto  75*8), 
w77 => Pw(106)( 77*8-1 downto  76*8), w78 => Pw(106)( 78*8-1 downto  77*8), w79 => Pw(106)( 79*8-1 downto  78*8), w80 => Pw(106)( 80*8-1 downto  79*8), 
w81 => Pw(106)( 81*8-1 downto  80*8), w82 => Pw(106)( 82*8-1 downto  81*8), w83 => Pw(106)( 83*8-1 downto  82*8), w84 => Pw(106)( 84*8-1 downto  83*8), 
w85 => Pw(106)( 85*8-1 downto  84*8), w86 => Pw(106)( 86*8-1 downto  85*8), w87 => Pw(106)( 87*8-1 downto  86*8), w88 => Pw(106)( 88*8-1 downto  87*8), 
w89 => Pw(106)( 89*8-1 downto  88*8), w90 => Pw(106)( 90*8-1 downto  89*8), w91 => Pw(106)( 91*8-1 downto  90*8), w92 => Pw(106)( 92*8-1 downto  91*8), 
w93 => Pw(106)( 93*8-1 downto  92*8), w94 => Pw(106)( 94*8-1 downto  93*8), w95 => Pw(106)( 95*8-1 downto  94*8), w96 => Pw(106)( 96*8-1 downto  95*8), 
w97 => Pw(106)( 97*8-1 downto  96*8), w98 => Pw(106)( 98*8-1 downto  97*8), w99 => Pw(106)( 99*8-1 downto  98*8), w100=> Pw(106)(100*8-1 downto  99*8), 
w101=> Pw(106)(101*8-1 downto 100*8), w102=> Pw(106)(102*8-1 downto 101*8), w103=> Pw(106)(103*8-1 downto 102*8), w104=> Pw(106)(104*8-1 downto 103*8), 
w105=> Pw(106)(105*8-1 downto 104*8), w106=> Pw(106)(106*8-1 downto 105*8), w107=> Pw(106)(107*8-1 downto 106*8), w108=> Pw(106)(108*8-1 downto 107*8), 
w109=> Pw(106)(109*8-1 downto 108*8), w110=> Pw(106)(110*8-1 downto 109*8), w111=> Pw(106)(111*8-1 downto 110*8), w112=> Pw(106)(112*8-1 downto 111*8), 
w113=> Pw(106)(113*8-1 downto 112*8), w114=> Pw(106)(114*8-1 downto 113*8), w115=> Pw(106)(115*8-1 downto 114*8), w116=> Pw(106)(116*8-1 downto 115*8), 
w117=> Pw(106)(117*8-1 downto 116*8), w118=> Pw(106)(118*8-1 downto 117*8), w119=> Pw(106)(119*8-1 downto 118*8), w120=> Pw(106)(120*8-1 downto 119*8), 
w121=> Pw(106)(121*8-1 downto 120*8), w122=> Pw(106)(122*8-1 downto 121*8), w123=> Pw(106)(123*8-1 downto 122*8), w124=> Pw(106)(124*8-1 downto 123*8), 
w125=> Pw(106)(125*8-1 downto 124*8), w126=> Pw(106)(126*8-1 downto 125*8), w127=> Pw(106)(127*8-1 downto 126*8), w128=> Pw(106)(128*8-1 downto 127*8), 
           d_out   => pca_d106_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_107_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(107)(     7 downto    0),   w02 => Pw(107)( 2*8-1 downto    8),   w03 => Pw(107)( 3*8-1 downto  2*8),   w04 => Pw(107)( 4*8-1 downto  3*8),   
w05 => Pw(107)( 5*8-1 downto  4*8),   w06 => Pw(107)( 6*8-1 downto  5*8),   w07 => Pw(107)( 7*8-1 downto  6*8),   w08 => Pw(107)( 8*8-1 downto  7*8),  
w09 => Pw(107)( 9*8-1 downto  8*8),   w10 => Pw(107)(10*8-1 downto  9*8),   w11 => Pw(107)(11*8-1 downto 10*8),   w12 => Pw(107)(12*8-1 downto 11*8),   
w13 => Pw(107)(13*8-1 downto 12*8),   w14 => Pw(107)(14*8-1 downto 13*8),   w15 => Pw(107)(15*8-1 downto 14*8),   w16 => Pw(107)(16*8-1 downto 15*8),  
w17 => Pw(107)(17*8-1 downto 16*8),   w18 => Pw(107)(18*8-1 downto 17*8),   w19 => Pw(107)(19*8-1 downto 18*8),   w20 => Pw(107)(20*8-1 downto 19*8),   
w21 => Pw(107)(21*8-1 downto 20*8),   w22 => Pw(107)(22*8-1 downto 21*8),   w23 => Pw(107)(23*8-1 downto 22*8),   w24 => Pw(107)(24*8-1 downto 23*8),  
w25 => Pw(107)(25*8-1 downto 24*8),   w26 => Pw(107)(26*8-1 downto 25*8),   w27 => Pw(107)(27*8-1 downto 26*8),   w28 => Pw(107)(28*8-1 downto 27*8),   
w29 => Pw(107)(29*8-1 downto 28*8),   w30 => Pw(107)(30*8-1 downto 29*8),   w31 => Pw(107)(31*8-1 downto 30*8),   w32 => Pw(107)(32*8-1 downto 31*8),  
w33 => Pw(107)(33*8-1 downto 32*8),   w34 => Pw(107)(34*8-1 downto 33*8),   w35 => Pw(107)(35*8-1 downto 34*8),   w36 => Pw(107)(36*8-1 downto 35*8),   
w37 => Pw(107)(37*8-1 downto 36*8),   w38 => Pw(107)(38*8-1 downto 37*8),   w39 => Pw(107)(39*8-1 downto 38*8),   w40 => Pw(107)(40*8-1 downto 39*8),  
w41 => Pw(107)(41*8-1 downto 40*8),   w42 => Pw(107)(42*8-1 downto 41*8),   w43 => Pw(107)(43*8-1 downto 42*8),   w44 => Pw(107)(44*8-1 downto 43*8),   
w45 => Pw(107)(45*8-1 downto 44*8),   w46 => Pw(107)(46*8-1 downto 45*8),   w47 => Pw(107)(47*8-1 downto 46*8),   w48 => Pw(107)(48*8-1 downto 47*8),  
w49 => Pw(107)(49*8-1 downto 48*8),   w50 => Pw(107)(50*8-1 downto 49*8),   w51 => Pw(107)(51*8-1 downto 50*8),   w52 => Pw(107)(52*8-1 downto 51*8),   
w53 => Pw(107)(53*8-1 downto 52*8),   w54 => Pw(107)(54*8-1 downto 53*8),   w55 => Pw(107)(55*8-1 downto 54*8),   w56 => Pw(107)(56*8-1 downto 55*8),  
w57 => Pw(107)(57*8-1 downto 56*8),   w58 => Pw(107)(58*8-1 downto 57*8),   w59 => Pw(107)(59*8-1 downto 58*8),   w60 => Pw(107)(60*8-1 downto 59*8),   
w61 => Pw(107)(61*8-1 downto 60*8),   w62 => Pw(107)(62*8-1 downto 61*8),   w63 => Pw(107)(63*8-1 downto 62*8),   w64 => Pw(107)(64*8-1 downto 63*8), 
w65 => Pw(107)( 65*8-1 downto  64*8), w66 => Pw(107)( 66*8-1 downto  65*8), w67 => Pw(107)( 67*8-1 downto  66*8), w68 => Pw(107)( 68*8-1 downto  67*8), 
w69 => Pw(107)( 69*8-1 downto  68*8), w70 => Pw(107)( 70*8-1 downto  69*8), w71 => Pw(107)( 71*8-1 downto  70*8), w72 => Pw(107)( 72*8-1 downto  71*8), 
w73 => Pw(107)( 73*8-1 downto  72*8), w74 => Pw(107)( 74*8-1 downto  73*8), w75 => Pw(107)( 75*8-1 downto  74*8), w76 => Pw(107)( 76*8-1 downto  75*8), 
w77 => Pw(107)( 77*8-1 downto  76*8), w78 => Pw(107)( 78*8-1 downto  77*8), w79 => Pw(107)( 79*8-1 downto  78*8), w80 => Pw(107)( 80*8-1 downto  79*8), 
w81 => Pw(107)( 81*8-1 downto  80*8), w82 => Pw(107)( 82*8-1 downto  81*8), w83 => Pw(107)( 83*8-1 downto  82*8), w84 => Pw(107)( 84*8-1 downto  83*8), 
w85 => Pw(107)( 85*8-1 downto  84*8), w86 => Pw(107)( 86*8-1 downto  85*8), w87 => Pw(107)( 87*8-1 downto  86*8), w88 => Pw(107)( 88*8-1 downto  87*8), 
w89 => Pw(107)( 89*8-1 downto  88*8), w90 => Pw(107)( 90*8-1 downto  89*8), w91 => Pw(107)( 91*8-1 downto  90*8), w92 => Pw(107)( 92*8-1 downto  91*8), 
w93 => Pw(107)( 93*8-1 downto  92*8), w94 => Pw(107)( 94*8-1 downto  93*8), w95 => Pw(107)( 95*8-1 downto  94*8), w96 => Pw(107)( 96*8-1 downto  95*8), 
w97 => Pw(107)( 97*8-1 downto  96*8), w98 => Pw(107)( 98*8-1 downto  97*8), w99 => Pw(107)( 99*8-1 downto  98*8), w100=> Pw(107)(100*8-1 downto  99*8), 
w101=> Pw(107)(101*8-1 downto 100*8), w102=> Pw(107)(102*8-1 downto 101*8), w103=> Pw(107)(103*8-1 downto 102*8), w104=> Pw(107)(104*8-1 downto 103*8), 
w105=> Pw(107)(105*8-1 downto 104*8), w106=> Pw(107)(106*8-1 downto 105*8), w107=> Pw(107)(107*8-1 downto 106*8), w108=> Pw(107)(108*8-1 downto 107*8), 
w109=> Pw(107)(109*8-1 downto 108*8), w110=> Pw(107)(110*8-1 downto 109*8), w111=> Pw(107)(111*8-1 downto 110*8), w112=> Pw(107)(112*8-1 downto 111*8), 
w113=> Pw(107)(113*8-1 downto 112*8), w114=> Pw(107)(114*8-1 downto 113*8), w115=> Pw(107)(115*8-1 downto 114*8), w116=> Pw(107)(116*8-1 downto 115*8), 
w117=> Pw(107)(117*8-1 downto 116*8), w118=> Pw(107)(118*8-1 downto 117*8), w119=> Pw(107)(119*8-1 downto 118*8), w120=> Pw(107)(120*8-1 downto 119*8), 
w121=> Pw(107)(121*8-1 downto 120*8), w122=> Pw(107)(122*8-1 downto 121*8), w123=> Pw(107)(123*8-1 downto 122*8), w124=> Pw(107)(124*8-1 downto 123*8), 
w125=> Pw(107)(125*8-1 downto 124*8), w126=> Pw(107)(126*8-1 downto 125*8), w127=> Pw(107)(127*8-1 downto 126*8), w128=> Pw(107)(128*8-1 downto 127*8), 
           d_out   => pca_d107_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_108_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(108)(     7 downto    0),   w02 => Pw(108)( 2*8-1 downto    8),   w03 => Pw(108)( 3*8-1 downto  2*8),   w04 => Pw(108)( 4*8-1 downto  3*8),   
w05 => Pw(108)( 5*8-1 downto  4*8),   w06 => Pw(108)( 6*8-1 downto  5*8),   w07 => Pw(108)( 7*8-1 downto  6*8),   w08 => Pw(108)( 8*8-1 downto  7*8),  
w09 => Pw(108)( 9*8-1 downto  8*8),   w10 => Pw(108)(10*8-1 downto  9*8),   w11 => Pw(108)(11*8-1 downto 10*8),   w12 => Pw(108)(12*8-1 downto 11*8),   
w13 => Pw(108)(13*8-1 downto 12*8),   w14 => Pw(108)(14*8-1 downto 13*8),   w15 => Pw(108)(15*8-1 downto 14*8),   w16 => Pw(108)(16*8-1 downto 15*8),  
w17 => Pw(108)(17*8-1 downto 16*8),   w18 => Pw(108)(18*8-1 downto 17*8),   w19 => Pw(108)(19*8-1 downto 18*8),   w20 => Pw(108)(20*8-1 downto 19*8),   
w21 => Pw(108)(21*8-1 downto 20*8),   w22 => Pw(108)(22*8-1 downto 21*8),   w23 => Pw(108)(23*8-1 downto 22*8),   w24 => Pw(108)(24*8-1 downto 23*8),  
w25 => Pw(108)(25*8-1 downto 24*8),   w26 => Pw(108)(26*8-1 downto 25*8),   w27 => Pw(108)(27*8-1 downto 26*8),   w28 => Pw(108)(28*8-1 downto 27*8),   
w29 => Pw(108)(29*8-1 downto 28*8),   w30 => Pw(108)(30*8-1 downto 29*8),   w31 => Pw(108)(31*8-1 downto 30*8),   w32 => Pw(108)(32*8-1 downto 31*8),  
w33 => Pw(108)(33*8-1 downto 32*8),   w34 => Pw(108)(34*8-1 downto 33*8),   w35 => Pw(108)(35*8-1 downto 34*8),   w36 => Pw(108)(36*8-1 downto 35*8),   
w37 => Pw(108)(37*8-1 downto 36*8),   w38 => Pw(108)(38*8-1 downto 37*8),   w39 => Pw(108)(39*8-1 downto 38*8),   w40 => Pw(108)(40*8-1 downto 39*8),  
w41 => Pw(108)(41*8-1 downto 40*8),   w42 => Pw(108)(42*8-1 downto 41*8),   w43 => Pw(108)(43*8-1 downto 42*8),   w44 => Pw(108)(44*8-1 downto 43*8),   
w45 => Pw(108)(45*8-1 downto 44*8),   w46 => Pw(108)(46*8-1 downto 45*8),   w47 => Pw(108)(47*8-1 downto 46*8),   w48 => Pw(108)(48*8-1 downto 47*8),  
w49 => Pw(108)(49*8-1 downto 48*8),   w50 => Pw(108)(50*8-1 downto 49*8),   w51 => Pw(108)(51*8-1 downto 50*8),   w52 => Pw(108)(52*8-1 downto 51*8),   
w53 => Pw(108)(53*8-1 downto 52*8),   w54 => Pw(108)(54*8-1 downto 53*8),   w55 => Pw(108)(55*8-1 downto 54*8),   w56 => Pw(108)(56*8-1 downto 55*8),  
w57 => Pw(108)(57*8-1 downto 56*8),   w58 => Pw(108)(58*8-1 downto 57*8),   w59 => Pw(108)(59*8-1 downto 58*8),   w60 => Pw(108)(60*8-1 downto 59*8),   
w61 => Pw(108)(61*8-1 downto 60*8),   w62 => Pw(108)(62*8-1 downto 61*8),   w63 => Pw(108)(63*8-1 downto 62*8),   w64 => Pw(108)(64*8-1 downto 63*8), 
w65 => Pw(108)( 65*8-1 downto  64*8), w66 => Pw(108)( 66*8-1 downto  65*8), w67 => Pw(108)( 67*8-1 downto  66*8), w68 => Pw(108)( 68*8-1 downto  67*8), 
w69 => Pw(108)( 69*8-1 downto  68*8), w70 => Pw(108)( 70*8-1 downto  69*8), w71 => Pw(108)( 71*8-1 downto  70*8), w72 => Pw(108)( 72*8-1 downto  71*8), 
w73 => Pw(108)( 73*8-1 downto  72*8), w74 => Pw(108)( 74*8-1 downto  73*8), w75 => Pw(108)( 75*8-1 downto  74*8), w76 => Pw(108)( 76*8-1 downto  75*8), 
w77 => Pw(108)( 77*8-1 downto  76*8), w78 => Pw(108)( 78*8-1 downto  77*8), w79 => Pw(108)( 79*8-1 downto  78*8), w80 => Pw(108)( 80*8-1 downto  79*8), 
w81 => Pw(108)( 81*8-1 downto  80*8), w82 => Pw(108)( 82*8-1 downto  81*8), w83 => Pw(108)( 83*8-1 downto  82*8), w84 => Pw(108)( 84*8-1 downto  83*8), 
w85 => Pw(108)( 85*8-1 downto  84*8), w86 => Pw(108)( 86*8-1 downto  85*8), w87 => Pw(108)( 87*8-1 downto  86*8), w88 => Pw(108)( 88*8-1 downto  87*8), 
w89 => Pw(108)( 89*8-1 downto  88*8), w90 => Pw(108)( 90*8-1 downto  89*8), w91 => Pw(108)( 91*8-1 downto  90*8), w92 => Pw(108)( 92*8-1 downto  91*8), 
w93 => Pw(108)( 93*8-1 downto  92*8), w94 => Pw(108)( 94*8-1 downto  93*8), w95 => Pw(108)( 95*8-1 downto  94*8), w96 => Pw(108)( 96*8-1 downto  95*8), 
w97 => Pw(108)( 97*8-1 downto  96*8), w98 => Pw(108)( 98*8-1 downto  97*8), w99 => Pw(108)( 99*8-1 downto  98*8), w100=> Pw(108)(100*8-1 downto  99*8), 
w101=> Pw(108)(101*8-1 downto 100*8), w102=> Pw(108)(102*8-1 downto 101*8), w103=> Pw(108)(103*8-1 downto 102*8), w104=> Pw(108)(104*8-1 downto 103*8), 
w105=> Pw(108)(105*8-1 downto 104*8), w106=> Pw(108)(106*8-1 downto 105*8), w107=> Pw(108)(107*8-1 downto 106*8), w108=> Pw(108)(108*8-1 downto 107*8), 
w109=> Pw(108)(109*8-1 downto 108*8), w110=> Pw(108)(110*8-1 downto 109*8), w111=> Pw(108)(111*8-1 downto 110*8), w112=> Pw(108)(112*8-1 downto 111*8), 
w113=> Pw(108)(113*8-1 downto 112*8), w114=> Pw(108)(114*8-1 downto 113*8), w115=> Pw(108)(115*8-1 downto 114*8), w116=> Pw(108)(116*8-1 downto 115*8), 
w117=> Pw(108)(117*8-1 downto 116*8), w118=> Pw(108)(118*8-1 downto 117*8), w119=> Pw(108)(119*8-1 downto 118*8), w120=> Pw(108)(120*8-1 downto 119*8), 
w121=> Pw(108)(121*8-1 downto 120*8), w122=> Pw(108)(122*8-1 downto 121*8), w123=> Pw(108)(123*8-1 downto 122*8), w124=> Pw(108)(124*8-1 downto 123*8), 
w125=> Pw(108)(125*8-1 downto 124*8), w126=> Pw(108)(126*8-1 downto 125*8), w127=> Pw(108)(127*8-1 downto 126*8), w128=> Pw(108)(128*8-1 downto 127*8), 
           d_out   => pca_d108_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_109_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(109)(     7 downto    0),   w02 => Pw(109)( 2*8-1 downto    8),   w03 => Pw(109)( 3*8-1 downto  2*8),   w04 => Pw(109)( 4*8-1 downto  3*8),   
w05 => Pw(109)( 5*8-1 downto  4*8),   w06 => Pw(109)( 6*8-1 downto  5*8),   w07 => Pw(109)( 7*8-1 downto  6*8),   w08 => Pw(109)( 8*8-1 downto  7*8),  
w09 => Pw(109)( 9*8-1 downto  8*8),   w10 => Pw(109)(10*8-1 downto  9*8),   w11 => Pw(109)(11*8-1 downto 10*8),   w12 => Pw(109)(12*8-1 downto 11*8),   
w13 => Pw(109)(13*8-1 downto 12*8),   w14 => Pw(109)(14*8-1 downto 13*8),   w15 => Pw(109)(15*8-1 downto 14*8),   w16 => Pw(109)(16*8-1 downto 15*8),  
w17 => Pw(109)(17*8-1 downto 16*8),   w18 => Pw(109)(18*8-1 downto 17*8),   w19 => Pw(109)(19*8-1 downto 18*8),   w20 => Pw(109)(20*8-1 downto 19*8),   
w21 => Pw(109)(21*8-1 downto 20*8),   w22 => Pw(109)(22*8-1 downto 21*8),   w23 => Pw(109)(23*8-1 downto 22*8),   w24 => Pw(109)(24*8-1 downto 23*8),  
w25 => Pw(109)(25*8-1 downto 24*8),   w26 => Pw(109)(26*8-1 downto 25*8),   w27 => Pw(109)(27*8-1 downto 26*8),   w28 => Pw(109)(28*8-1 downto 27*8),   
w29 => Pw(109)(29*8-1 downto 28*8),   w30 => Pw(109)(30*8-1 downto 29*8),   w31 => Pw(109)(31*8-1 downto 30*8),   w32 => Pw(109)(32*8-1 downto 31*8),  
w33 => Pw(109)(33*8-1 downto 32*8),   w34 => Pw(109)(34*8-1 downto 33*8),   w35 => Pw(109)(35*8-1 downto 34*8),   w36 => Pw(109)(36*8-1 downto 35*8),   
w37 => Pw(109)(37*8-1 downto 36*8),   w38 => Pw(109)(38*8-1 downto 37*8),   w39 => Pw(109)(39*8-1 downto 38*8),   w40 => Pw(109)(40*8-1 downto 39*8),  
w41 => Pw(109)(41*8-1 downto 40*8),   w42 => Pw(109)(42*8-1 downto 41*8),   w43 => Pw(109)(43*8-1 downto 42*8),   w44 => Pw(109)(44*8-1 downto 43*8),   
w45 => Pw(109)(45*8-1 downto 44*8),   w46 => Pw(109)(46*8-1 downto 45*8),   w47 => Pw(109)(47*8-1 downto 46*8),   w48 => Pw(109)(48*8-1 downto 47*8),  
w49 => Pw(109)(49*8-1 downto 48*8),   w50 => Pw(109)(50*8-1 downto 49*8),   w51 => Pw(109)(51*8-1 downto 50*8),   w52 => Pw(109)(52*8-1 downto 51*8),   
w53 => Pw(109)(53*8-1 downto 52*8),   w54 => Pw(109)(54*8-1 downto 53*8),   w55 => Pw(109)(55*8-1 downto 54*8),   w56 => Pw(109)(56*8-1 downto 55*8),  
w57 => Pw(109)(57*8-1 downto 56*8),   w58 => Pw(109)(58*8-1 downto 57*8),   w59 => Pw(109)(59*8-1 downto 58*8),   w60 => Pw(109)(60*8-1 downto 59*8),   
w61 => Pw(109)(61*8-1 downto 60*8),   w62 => Pw(109)(62*8-1 downto 61*8),   w63 => Pw(109)(63*8-1 downto 62*8),   w64 => Pw(109)(64*8-1 downto 63*8), 
w65 => Pw(109)( 65*8-1 downto  64*8), w66 => Pw(109)( 66*8-1 downto  65*8), w67 => Pw(109)( 67*8-1 downto  66*8), w68 => Pw(109)( 68*8-1 downto  67*8), 
w69 => Pw(109)( 69*8-1 downto  68*8), w70 => Pw(109)( 70*8-1 downto  69*8), w71 => Pw(109)( 71*8-1 downto  70*8), w72 => Pw(109)( 72*8-1 downto  71*8), 
w73 => Pw(109)( 73*8-1 downto  72*8), w74 => Pw(109)( 74*8-1 downto  73*8), w75 => Pw(109)( 75*8-1 downto  74*8), w76 => Pw(109)( 76*8-1 downto  75*8), 
w77 => Pw(109)( 77*8-1 downto  76*8), w78 => Pw(109)( 78*8-1 downto  77*8), w79 => Pw(109)( 79*8-1 downto  78*8), w80 => Pw(109)( 80*8-1 downto  79*8), 
w81 => Pw(109)( 81*8-1 downto  80*8), w82 => Pw(109)( 82*8-1 downto  81*8), w83 => Pw(109)( 83*8-1 downto  82*8), w84 => Pw(109)( 84*8-1 downto  83*8), 
w85 => Pw(109)( 85*8-1 downto  84*8), w86 => Pw(109)( 86*8-1 downto  85*8), w87 => Pw(109)( 87*8-1 downto  86*8), w88 => Pw(109)( 88*8-1 downto  87*8), 
w89 => Pw(109)( 89*8-1 downto  88*8), w90 => Pw(109)( 90*8-1 downto  89*8), w91 => Pw(109)( 91*8-1 downto  90*8), w92 => Pw(109)( 92*8-1 downto  91*8), 
w93 => Pw(109)( 93*8-1 downto  92*8), w94 => Pw(109)( 94*8-1 downto  93*8), w95 => Pw(109)( 95*8-1 downto  94*8), w96 => Pw(109)( 96*8-1 downto  95*8), 
w97 => Pw(109)( 97*8-1 downto  96*8), w98 => Pw(109)( 98*8-1 downto  97*8), w99 => Pw(109)( 99*8-1 downto  98*8), w100=> Pw(109)(100*8-1 downto  99*8), 
w101=> Pw(109)(101*8-1 downto 100*8), w102=> Pw(109)(102*8-1 downto 101*8), w103=> Pw(109)(103*8-1 downto 102*8), w104=> Pw(109)(104*8-1 downto 103*8), 
w105=> Pw(109)(105*8-1 downto 104*8), w106=> Pw(109)(106*8-1 downto 105*8), w107=> Pw(109)(107*8-1 downto 106*8), w108=> Pw(109)(108*8-1 downto 107*8), 
w109=> Pw(109)(109*8-1 downto 108*8), w110=> Pw(109)(110*8-1 downto 109*8), w111=> Pw(109)(111*8-1 downto 110*8), w112=> Pw(109)(112*8-1 downto 111*8), 
w113=> Pw(109)(113*8-1 downto 112*8), w114=> Pw(109)(114*8-1 downto 113*8), w115=> Pw(109)(115*8-1 downto 114*8), w116=> Pw(109)(116*8-1 downto 115*8), 
w117=> Pw(109)(117*8-1 downto 116*8), w118=> Pw(109)(118*8-1 downto 117*8), w119=> Pw(109)(119*8-1 downto 118*8), w120=> Pw(109)(120*8-1 downto 119*8), 
w121=> Pw(109)(121*8-1 downto 120*8), w122=> Pw(109)(122*8-1 downto 121*8), w123=> Pw(109)(123*8-1 downto 122*8), w124=> Pw(109)(124*8-1 downto 123*8), 
w125=> Pw(109)(125*8-1 downto 124*8), w126=> Pw(109)(126*8-1 downto 125*8), w127=> Pw(109)(127*8-1 downto 126*8), w128=> Pw(109)(128*8-1 downto 127*8), 
           d_out   => pca_d109_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_110_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(110)(     7 downto    0),   w02 => Pw(110)( 2*8-1 downto    8),   w03 => Pw(110)( 3*8-1 downto  2*8),   w04 => Pw(110)( 4*8-1 downto  3*8),   
w05 => Pw(110)( 5*8-1 downto  4*8),   w06 => Pw(110)( 6*8-1 downto  5*8),   w07 => Pw(110)( 7*8-1 downto  6*8),   w08 => Pw(110)( 8*8-1 downto  7*8),  
w09 => Pw(110)( 9*8-1 downto  8*8),   w10 => Pw(110)(10*8-1 downto  9*8),   w11 => Pw(110)(11*8-1 downto 10*8),   w12 => Pw(110)(12*8-1 downto 11*8),   
w13 => Pw(110)(13*8-1 downto 12*8),   w14 => Pw(110)(14*8-1 downto 13*8),   w15 => Pw(110)(15*8-1 downto 14*8),   w16 => Pw(110)(16*8-1 downto 15*8),  
w17 => Pw(110)(17*8-1 downto 16*8),   w18 => Pw(110)(18*8-1 downto 17*8),   w19 => Pw(110)(19*8-1 downto 18*8),   w20 => Pw(110)(20*8-1 downto 19*8),   
w21 => Pw(110)(21*8-1 downto 20*8),   w22 => Pw(110)(22*8-1 downto 21*8),   w23 => Pw(110)(23*8-1 downto 22*8),   w24 => Pw(110)(24*8-1 downto 23*8),  
w25 => Pw(110)(25*8-1 downto 24*8),   w26 => Pw(110)(26*8-1 downto 25*8),   w27 => Pw(110)(27*8-1 downto 26*8),   w28 => Pw(110)(28*8-1 downto 27*8),   
w29 => Pw(110)(29*8-1 downto 28*8),   w30 => Pw(110)(30*8-1 downto 29*8),   w31 => Pw(110)(31*8-1 downto 30*8),   w32 => Pw(110)(32*8-1 downto 31*8),  
w33 => Pw(110)(33*8-1 downto 32*8),   w34 => Pw(110)(34*8-1 downto 33*8),   w35 => Pw(110)(35*8-1 downto 34*8),   w36 => Pw(110)(36*8-1 downto 35*8),   
w37 => Pw(110)(37*8-1 downto 36*8),   w38 => Pw(110)(38*8-1 downto 37*8),   w39 => Pw(110)(39*8-1 downto 38*8),   w40 => Pw(110)(40*8-1 downto 39*8),  
w41 => Pw(110)(41*8-1 downto 40*8),   w42 => Pw(110)(42*8-1 downto 41*8),   w43 => Pw(110)(43*8-1 downto 42*8),   w44 => Pw(110)(44*8-1 downto 43*8),   
w45 => Pw(110)(45*8-1 downto 44*8),   w46 => Pw(110)(46*8-1 downto 45*8),   w47 => Pw(110)(47*8-1 downto 46*8),   w48 => Pw(110)(48*8-1 downto 47*8),  
w49 => Pw(110)(49*8-1 downto 48*8),   w50 => Pw(110)(50*8-1 downto 49*8),   w51 => Pw(110)(51*8-1 downto 50*8),   w52 => Pw(110)(52*8-1 downto 51*8),   
w53 => Pw(110)(53*8-1 downto 52*8),   w54 => Pw(110)(54*8-1 downto 53*8),   w55 => Pw(110)(55*8-1 downto 54*8),   w56 => Pw(110)(56*8-1 downto 55*8),  
w57 => Pw(110)(57*8-1 downto 56*8),   w58 => Pw(110)(58*8-1 downto 57*8),   w59 => Pw(110)(59*8-1 downto 58*8),   w60 => Pw(110)(60*8-1 downto 59*8),   
w61 => Pw(110)(61*8-1 downto 60*8),   w62 => Pw(110)(62*8-1 downto 61*8),   w63 => Pw(110)(63*8-1 downto 62*8),   w64 => Pw(110)(64*8-1 downto 63*8), 
w65 => Pw(110)( 65*8-1 downto  64*8), w66 => Pw(110)( 66*8-1 downto  65*8), w67 => Pw(110)( 67*8-1 downto  66*8), w68 => Pw(110)( 68*8-1 downto  67*8), 
w69 => Pw(110)( 69*8-1 downto  68*8), w70 => Pw(110)( 70*8-1 downto  69*8), w71 => Pw(110)( 71*8-1 downto  70*8), w72 => Pw(110)( 72*8-1 downto  71*8), 
w73 => Pw(110)( 73*8-1 downto  72*8), w74 => Pw(110)( 74*8-1 downto  73*8), w75 => Pw(110)( 75*8-1 downto  74*8), w76 => Pw(110)( 76*8-1 downto  75*8), 
w77 => Pw(110)( 77*8-1 downto  76*8), w78 => Pw(110)( 78*8-1 downto  77*8), w79 => Pw(110)( 79*8-1 downto  78*8), w80 => Pw(110)( 80*8-1 downto  79*8), 
w81 => Pw(110)( 81*8-1 downto  80*8), w82 => Pw(110)( 82*8-1 downto  81*8), w83 => Pw(110)( 83*8-1 downto  82*8), w84 => Pw(110)( 84*8-1 downto  83*8), 
w85 => Pw(110)( 85*8-1 downto  84*8), w86 => Pw(110)( 86*8-1 downto  85*8), w87 => Pw(110)( 87*8-1 downto  86*8), w88 => Pw(110)( 88*8-1 downto  87*8), 
w89 => Pw(110)( 89*8-1 downto  88*8), w90 => Pw(110)( 90*8-1 downto  89*8), w91 => Pw(110)( 91*8-1 downto  90*8), w92 => Pw(110)( 92*8-1 downto  91*8), 
w93 => Pw(110)( 93*8-1 downto  92*8), w94 => Pw(110)( 94*8-1 downto  93*8), w95 => Pw(110)( 95*8-1 downto  94*8), w96 => Pw(110)( 96*8-1 downto  95*8), 
w97 => Pw(110)( 97*8-1 downto  96*8), w98 => Pw(110)( 98*8-1 downto  97*8), w99 => Pw(110)( 99*8-1 downto  98*8), w100=> Pw(110)(100*8-1 downto  99*8), 
w101=> Pw(110)(101*8-1 downto 100*8), w102=> Pw(110)(102*8-1 downto 101*8), w103=> Pw(110)(103*8-1 downto 102*8), w104=> Pw(110)(104*8-1 downto 103*8), 
w105=> Pw(110)(105*8-1 downto 104*8), w106=> Pw(110)(106*8-1 downto 105*8), w107=> Pw(110)(107*8-1 downto 106*8), w108=> Pw(110)(108*8-1 downto 107*8), 
w109=> Pw(110)(109*8-1 downto 108*8), w110=> Pw(110)(110*8-1 downto 109*8), w111=> Pw(110)(111*8-1 downto 110*8), w112=> Pw(110)(112*8-1 downto 111*8), 
w113=> Pw(110)(113*8-1 downto 112*8), w114=> Pw(110)(114*8-1 downto 113*8), w115=> Pw(110)(115*8-1 downto 114*8), w116=> Pw(110)(116*8-1 downto 115*8), 
w117=> Pw(110)(117*8-1 downto 116*8), w118=> Pw(110)(118*8-1 downto 117*8), w119=> Pw(110)(119*8-1 downto 118*8), w120=> Pw(110)(120*8-1 downto 119*8), 
w121=> Pw(110)(121*8-1 downto 120*8), w122=> Pw(110)(122*8-1 downto 121*8), w123=> Pw(110)(123*8-1 downto 122*8), w124=> Pw(110)(124*8-1 downto 123*8), 
w125=> Pw(110)(125*8-1 downto 124*8), w126=> Pw(110)(126*8-1 downto 125*8), w127=> Pw(110)(127*8-1 downto 126*8), w128=> Pw(110)(128*8-1 downto 127*8), 
           d_out   => pca_d110_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_111_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(111)(     7 downto    0),   w02 => Pw(111)( 2*8-1 downto    8),   w03 => Pw(111)( 3*8-1 downto  2*8),   w04 => Pw(111)( 4*8-1 downto  3*8),   
w05 => Pw(111)( 5*8-1 downto  4*8),   w06 => Pw(111)( 6*8-1 downto  5*8),   w07 => Pw(111)( 7*8-1 downto  6*8),   w08 => Pw(111)( 8*8-1 downto  7*8),  
w09 => Pw(111)( 9*8-1 downto  8*8),   w10 => Pw(111)(10*8-1 downto  9*8),   w11 => Pw(111)(11*8-1 downto 10*8),   w12 => Pw(111)(12*8-1 downto 11*8),   
w13 => Pw(111)(13*8-1 downto 12*8),   w14 => Pw(111)(14*8-1 downto 13*8),   w15 => Pw(111)(15*8-1 downto 14*8),   w16 => Pw(111)(16*8-1 downto 15*8),  
w17 => Pw(111)(17*8-1 downto 16*8),   w18 => Pw(111)(18*8-1 downto 17*8),   w19 => Pw(111)(19*8-1 downto 18*8),   w20 => Pw(111)(20*8-1 downto 19*8),   
w21 => Pw(111)(21*8-1 downto 20*8),   w22 => Pw(111)(22*8-1 downto 21*8),   w23 => Pw(111)(23*8-1 downto 22*8),   w24 => Pw(111)(24*8-1 downto 23*8),  
w25 => Pw(111)(25*8-1 downto 24*8),   w26 => Pw(111)(26*8-1 downto 25*8),   w27 => Pw(111)(27*8-1 downto 26*8),   w28 => Pw(111)(28*8-1 downto 27*8),   
w29 => Pw(111)(29*8-1 downto 28*8),   w30 => Pw(111)(30*8-1 downto 29*8),   w31 => Pw(111)(31*8-1 downto 30*8),   w32 => Pw(111)(32*8-1 downto 31*8),  
w33 => Pw(111)(33*8-1 downto 32*8),   w34 => Pw(111)(34*8-1 downto 33*8),   w35 => Pw(111)(35*8-1 downto 34*8),   w36 => Pw(111)(36*8-1 downto 35*8),   
w37 => Pw(111)(37*8-1 downto 36*8),   w38 => Pw(111)(38*8-1 downto 37*8),   w39 => Pw(111)(39*8-1 downto 38*8),   w40 => Pw(111)(40*8-1 downto 39*8),  
w41 => Pw(111)(41*8-1 downto 40*8),   w42 => Pw(111)(42*8-1 downto 41*8),   w43 => Pw(111)(43*8-1 downto 42*8),   w44 => Pw(111)(44*8-1 downto 43*8),   
w45 => Pw(111)(45*8-1 downto 44*8),   w46 => Pw(111)(46*8-1 downto 45*8),   w47 => Pw(111)(47*8-1 downto 46*8),   w48 => Pw(111)(48*8-1 downto 47*8),  
w49 => Pw(111)(49*8-1 downto 48*8),   w50 => Pw(111)(50*8-1 downto 49*8),   w51 => Pw(111)(51*8-1 downto 50*8),   w52 => Pw(111)(52*8-1 downto 51*8),   
w53 => Pw(111)(53*8-1 downto 52*8),   w54 => Pw(111)(54*8-1 downto 53*8),   w55 => Pw(111)(55*8-1 downto 54*8),   w56 => Pw(111)(56*8-1 downto 55*8),  
w57 => Pw(111)(57*8-1 downto 56*8),   w58 => Pw(111)(58*8-1 downto 57*8),   w59 => Pw(111)(59*8-1 downto 58*8),   w60 => Pw(111)(60*8-1 downto 59*8),   
w61 => Pw(111)(61*8-1 downto 60*8),   w62 => Pw(111)(62*8-1 downto 61*8),   w63 => Pw(111)(63*8-1 downto 62*8),   w64 => Pw(111)(64*8-1 downto 63*8), 
w65 => Pw(111)( 65*8-1 downto  64*8), w66 => Pw(111)( 66*8-1 downto  65*8), w67 => Pw(111)( 67*8-1 downto  66*8), w68 => Pw(111)( 68*8-1 downto  67*8), 
w69 => Pw(111)( 69*8-1 downto  68*8), w70 => Pw(111)( 70*8-1 downto  69*8), w71 => Pw(111)( 71*8-1 downto  70*8), w72 => Pw(111)( 72*8-1 downto  71*8), 
w73 => Pw(111)( 73*8-1 downto  72*8), w74 => Pw(111)( 74*8-1 downto  73*8), w75 => Pw(111)( 75*8-1 downto  74*8), w76 => Pw(111)( 76*8-1 downto  75*8), 
w77 => Pw(111)( 77*8-1 downto  76*8), w78 => Pw(111)( 78*8-1 downto  77*8), w79 => Pw(111)( 79*8-1 downto  78*8), w80 => Pw(111)( 80*8-1 downto  79*8), 
w81 => Pw(111)( 81*8-1 downto  80*8), w82 => Pw(111)( 82*8-1 downto  81*8), w83 => Pw(111)( 83*8-1 downto  82*8), w84 => Pw(111)( 84*8-1 downto  83*8), 
w85 => Pw(111)( 85*8-1 downto  84*8), w86 => Pw(111)( 86*8-1 downto  85*8), w87 => Pw(111)( 87*8-1 downto  86*8), w88 => Pw(111)( 88*8-1 downto  87*8), 
w89 => Pw(111)( 89*8-1 downto  88*8), w90 => Pw(111)( 90*8-1 downto  89*8), w91 => Pw(111)( 91*8-1 downto  90*8), w92 => Pw(111)( 92*8-1 downto  91*8), 
w93 => Pw(111)( 93*8-1 downto  92*8), w94 => Pw(111)( 94*8-1 downto  93*8), w95 => Pw(111)( 95*8-1 downto  94*8), w96 => Pw(111)( 96*8-1 downto  95*8), 
w97 => Pw(111)( 97*8-1 downto  96*8), w98 => Pw(111)( 98*8-1 downto  97*8), w99 => Pw(111)( 99*8-1 downto  98*8), w100=> Pw(111)(100*8-1 downto  99*8), 
w101=> Pw(111)(101*8-1 downto 100*8), w102=> Pw(111)(102*8-1 downto 101*8), w103=> Pw(111)(103*8-1 downto 102*8), w104=> Pw(111)(104*8-1 downto 103*8), 
w105=> Pw(111)(105*8-1 downto 104*8), w106=> Pw(111)(106*8-1 downto 105*8), w107=> Pw(111)(107*8-1 downto 106*8), w108=> Pw(111)(108*8-1 downto 107*8), 
w109=> Pw(111)(109*8-1 downto 108*8), w110=> Pw(111)(110*8-1 downto 109*8), w111=> Pw(111)(111*8-1 downto 110*8), w112=> Pw(111)(112*8-1 downto 111*8), 
w113=> Pw(111)(113*8-1 downto 112*8), w114=> Pw(111)(114*8-1 downto 113*8), w115=> Pw(111)(115*8-1 downto 114*8), w116=> Pw(111)(116*8-1 downto 115*8), 
w117=> Pw(111)(117*8-1 downto 116*8), w118=> Pw(111)(118*8-1 downto 117*8), w119=> Pw(111)(119*8-1 downto 118*8), w120=> Pw(111)(120*8-1 downto 119*8), 
w121=> Pw(111)(121*8-1 downto 120*8), w122=> Pw(111)(122*8-1 downto 121*8), w123=> Pw(111)(123*8-1 downto 122*8), w124=> Pw(111)(124*8-1 downto 123*8), 
w125=> Pw(111)(125*8-1 downto 124*8), w126=> Pw(111)(126*8-1 downto 125*8), w127=> Pw(111)(127*8-1 downto 126*8), w128=> Pw(111)(128*8-1 downto 127*8), 
           d_out   => pca_d111_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_112_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(112)(     7 downto    0),   w02 => Pw(112)( 2*8-1 downto    8),   w03 => Pw(112)( 3*8-1 downto  2*8),   w04 => Pw(112)( 4*8-1 downto  3*8),   
w05 => Pw(112)( 5*8-1 downto  4*8),   w06 => Pw(112)( 6*8-1 downto  5*8),   w07 => Pw(112)( 7*8-1 downto  6*8),   w08 => Pw(112)( 8*8-1 downto  7*8),  
w09 => Pw(112)( 9*8-1 downto  8*8),   w10 => Pw(112)(10*8-1 downto  9*8),   w11 => Pw(112)(11*8-1 downto 10*8),   w12 => Pw(112)(12*8-1 downto 11*8),   
w13 => Pw(112)(13*8-1 downto 12*8),   w14 => Pw(112)(14*8-1 downto 13*8),   w15 => Pw(112)(15*8-1 downto 14*8),   w16 => Pw(112)(16*8-1 downto 15*8),  
w17 => Pw(112)(17*8-1 downto 16*8),   w18 => Pw(112)(18*8-1 downto 17*8),   w19 => Pw(112)(19*8-1 downto 18*8),   w20 => Pw(112)(20*8-1 downto 19*8),   
w21 => Pw(112)(21*8-1 downto 20*8),   w22 => Pw(112)(22*8-1 downto 21*8),   w23 => Pw(112)(23*8-1 downto 22*8),   w24 => Pw(112)(24*8-1 downto 23*8),  
w25 => Pw(112)(25*8-1 downto 24*8),   w26 => Pw(112)(26*8-1 downto 25*8),   w27 => Pw(112)(27*8-1 downto 26*8),   w28 => Pw(112)(28*8-1 downto 27*8),   
w29 => Pw(112)(29*8-1 downto 28*8),   w30 => Pw(112)(30*8-1 downto 29*8),   w31 => Pw(112)(31*8-1 downto 30*8),   w32 => Pw(112)(32*8-1 downto 31*8),  
w33 => Pw(112)(33*8-1 downto 32*8),   w34 => Pw(112)(34*8-1 downto 33*8),   w35 => Pw(112)(35*8-1 downto 34*8),   w36 => Pw(112)(36*8-1 downto 35*8),   
w37 => Pw(112)(37*8-1 downto 36*8),   w38 => Pw(112)(38*8-1 downto 37*8),   w39 => Pw(112)(39*8-1 downto 38*8),   w40 => Pw(112)(40*8-1 downto 39*8),  
w41 => Pw(112)(41*8-1 downto 40*8),   w42 => Pw(112)(42*8-1 downto 41*8),   w43 => Pw(112)(43*8-1 downto 42*8),   w44 => Pw(112)(44*8-1 downto 43*8),   
w45 => Pw(112)(45*8-1 downto 44*8),   w46 => Pw(112)(46*8-1 downto 45*8),   w47 => Pw(112)(47*8-1 downto 46*8),   w48 => Pw(112)(48*8-1 downto 47*8),  
w49 => Pw(112)(49*8-1 downto 48*8),   w50 => Pw(112)(50*8-1 downto 49*8),   w51 => Pw(112)(51*8-1 downto 50*8),   w52 => Pw(112)(52*8-1 downto 51*8),   
w53 => Pw(112)(53*8-1 downto 52*8),   w54 => Pw(112)(54*8-1 downto 53*8),   w55 => Pw(112)(55*8-1 downto 54*8),   w56 => Pw(112)(56*8-1 downto 55*8),  
w57 => Pw(112)(57*8-1 downto 56*8),   w58 => Pw(112)(58*8-1 downto 57*8),   w59 => Pw(112)(59*8-1 downto 58*8),   w60 => Pw(112)(60*8-1 downto 59*8),   
w61 => Pw(112)(61*8-1 downto 60*8),   w62 => Pw(112)(62*8-1 downto 61*8),   w63 => Pw(112)(63*8-1 downto 62*8),   w64 => Pw(112)(64*8-1 downto 63*8), 
w65 => Pw(112)( 65*8-1 downto  64*8), w66 => Pw(112)( 66*8-1 downto  65*8), w67 => Pw(112)( 67*8-1 downto  66*8), w68 => Pw(112)( 68*8-1 downto  67*8), 
w69 => Pw(112)( 69*8-1 downto  68*8), w70 => Pw(112)( 70*8-1 downto  69*8), w71 => Pw(112)( 71*8-1 downto  70*8), w72 => Pw(112)( 72*8-1 downto  71*8), 
w73 => Pw(112)( 73*8-1 downto  72*8), w74 => Pw(112)( 74*8-1 downto  73*8), w75 => Pw(112)( 75*8-1 downto  74*8), w76 => Pw(112)( 76*8-1 downto  75*8), 
w77 => Pw(112)( 77*8-1 downto  76*8), w78 => Pw(112)( 78*8-1 downto  77*8), w79 => Pw(112)( 79*8-1 downto  78*8), w80 => Pw(112)( 80*8-1 downto  79*8), 
w81 => Pw(112)( 81*8-1 downto  80*8), w82 => Pw(112)( 82*8-1 downto  81*8), w83 => Pw(112)( 83*8-1 downto  82*8), w84 => Pw(112)( 84*8-1 downto  83*8), 
w85 => Pw(112)( 85*8-1 downto  84*8), w86 => Pw(112)( 86*8-1 downto  85*8), w87 => Pw(112)( 87*8-1 downto  86*8), w88 => Pw(112)( 88*8-1 downto  87*8), 
w89 => Pw(112)( 89*8-1 downto  88*8), w90 => Pw(112)( 90*8-1 downto  89*8), w91 => Pw(112)( 91*8-1 downto  90*8), w92 => Pw(112)( 92*8-1 downto  91*8), 
w93 => Pw(112)( 93*8-1 downto  92*8), w94 => Pw(112)( 94*8-1 downto  93*8), w95 => Pw(112)( 95*8-1 downto  94*8), w96 => Pw(112)( 96*8-1 downto  95*8), 
w97 => Pw(112)( 97*8-1 downto  96*8), w98 => Pw(112)( 98*8-1 downto  97*8), w99 => Pw(112)( 99*8-1 downto  98*8), w100=> Pw(112)(100*8-1 downto  99*8), 
w101=> Pw(112)(101*8-1 downto 100*8), w102=> Pw(112)(102*8-1 downto 101*8), w103=> Pw(112)(103*8-1 downto 102*8), w104=> Pw(112)(104*8-1 downto 103*8), 
w105=> Pw(112)(105*8-1 downto 104*8), w106=> Pw(112)(106*8-1 downto 105*8), w107=> Pw(112)(107*8-1 downto 106*8), w108=> Pw(112)(108*8-1 downto 107*8), 
w109=> Pw(112)(109*8-1 downto 108*8), w110=> Pw(112)(110*8-1 downto 109*8), w111=> Pw(112)(111*8-1 downto 110*8), w112=> Pw(112)(112*8-1 downto 111*8), 
w113=> Pw(112)(113*8-1 downto 112*8), w114=> Pw(112)(114*8-1 downto 113*8), w115=> Pw(112)(115*8-1 downto 114*8), w116=> Pw(112)(116*8-1 downto 115*8), 
w117=> Pw(112)(117*8-1 downto 116*8), w118=> Pw(112)(118*8-1 downto 117*8), w119=> Pw(112)(119*8-1 downto 118*8), w120=> Pw(112)(120*8-1 downto 119*8), 
w121=> Pw(112)(121*8-1 downto 120*8), w122=> Pw(112)(122*8-1 downto 121*8), w123=> Pw(112)(123*8-1 downto 122*8), w124=> Pw(112)(124*8-1 downto 123*8), 
w125=> Pw(112)(125*8-1 downto 124*8), w126=> Pw(112)(126*8-1 downto 125*8), w127=> Pw(112)(127*8-1 downto 126*8), w128=> Pw(112)(128*8-1 downto 127*8), 
           d_out   => pca_d112_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_113_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(113)(     7 downto    0),   w02 => Pw(113)( 2*8-1 downto    8),   w03 => Pw(113)( 3*8-1 downto  2*8),   w04 => Pw(113)( 4*8-1 downto  3*8),   
w05 => Pw(113)( 5*8-1 downto  4*8),   w06 => Pw(113)( 6*8-1 downto  5*8),   w07 => Pw(113)( 7*8-1 downto  6*8),   w08 => Pw(113)( 8*8-1 downto  7*8),  
w09 => Pw(113)( 9*8-1 downto  8*8),   w10 => Pw(113)(10*8-1 downto  9*8),   w11 => Pw(113)(11*8-1 downto 10*8),   w12 => Pw(113)(12*8-1 downto 11*8),   
w13 => Pw(113)(13*8-1 downto 12*8),   w14 => Pw(113)(14*8-1 downto 13*8),   w15 => Pw(113)(15*8-1 downto 14*8),   w16 => Pw(113)(16*8-1 downto 15*8),  
w17 => Pw(113)(17*8-1 downto 16*8),   w18 => Pw(113)(18*8-1 downto 17*8),   w19 => Pw(113)(19*8-1 downto 18*8),   w20 => Pw(113)(20*8-1 downto 19*8),   
w21 => Pw(113)(21*8-1 downto 20*8),   w22 => Pw(113)(22*8-1 downto 21*8),   w23 => Pw(113)(23*8-1 downto 22*8),   w24 => Pw(113)(24*8-1 downto 23*8),  
w25 => Pw(113)(25*8-1 downto 24*8),   w26 => Pw(113)(26*8-1 downto 25*8),   w27 => Pw(113)(27*8-1 downto 26*8),   w28 => Pw(113)(28*8-1 downto 27*8),   
w29 => Pw(113)(29*8-1 downto 28*8),   w30 => Pw(113)(30*8-1 downto 29*8),   w31 => Pw(113)(31*8-1 downto 30*8),   w32 => Pw(113)(32*8-1 downto 31*8),  
w33 => Pw(113)(33*8-1 downto 32*8),   w34 => Pw(113)(34*8-1 downto 33*8),   w35 => Pw(113)(35*8-1 downto 34*8),   w36 => Pw(113)(36*8-1 downto 35*8),   
w37 => Pw(113)(37*8-1 downto 36*8),   w38 => Pw(113)(38*8-1 downto 37*8),   w39 => Pw(113)(39*8-1 downto 38*8),   w40 => Pw(113)(40*8-1 downto 39*8),  
w41 => Pw(113)(41*8-1 downto 40*8),   w42 => Pw(113)(42*8-1 downto 41*8),   w43 => Pw(113)(43*8-1 downto 42*8),   w44 => Pw(113)(44*8-1 downto 43*8),   
w45 => Pw(113)(45*8-1 downto 44*8),   w46 => Pw(113)(46*8-1 downto 45*8),   w47 => Pw(113)(47*8-1 downto 46*8),   w48 => Pw(113)(48*8-1 downto 47*8),  
w49 => Pw(113)(49*8-1 downto 48*8),   w50 => Pw(113)(50*8-1 downto 49*8),   w51 => Pw(113)(51*8-1 downto 50*8),   w52 => Pw(113)(52*8-1 downto 51*8),   
w53 => Pw(113)(53*8-1 downto 52*8),   w54 => Pw(113)(54*8-1 downto 53*8),   w55 => Pw(113)(55*8-1 downto 54*8),   w56 => Pw(113)(56*8-1 downto 55*8),  
w57 => Pw(113)(57*8-1 downto 56*8),   w58 => Pw(113)(58*8-1 downto 57*8),   w59 => Pw(113)(59*8-1 downto 58*8),   w60 => Pw(113)(60*8-1 downto 59*8),   
w61 => Pw(113)(61*8-1 downto 60*8),   w62 => Pw(113)(62*8-1 downto 61*8),   w63 => Pw(113)(63*8-1 downto 62*8),   w64 => Pw(113)(64*8-1 downto 63*8), 
w65 => Pw(113)( 65*8-1 downto  64*8), w66 => Pw(113)( 66*8-1 downto  65*8), w67 => Pw(113)( 67*8-1 downto  66*8), w68 => Pw(113)( 68*8-1 downto  67*8), 
w69 => Pw(113)( 69*8-1 downto  68*8), w70 => Pw(113)( 70*8-1 downto  69*8), w71 => Pw(113)( 71*8-1 downto  70*8), w72 => Pw(113)( 72*8-1 downto  71*8), 
w73 => Pw(113)( 73*8-1 downto  72*8), w74 => Pw(113)( 74*8-1 downto  73*8), w75 => Pw(113)( 75*8-1 downto  74*8), w76 => Pw(113)( 76*8-1 downto  75*8), 
w77 => Pw(113)( 77*8-1 downto  76*8), w78 => Pw(113)( 78*8-1 downto  77*8), w79 => Pw(113)( 79*8-1 downto  78*8), w80 => Pw(113)( 80*8-1 downto  79*8), 
w81 => Pw(113)( 81*8-1 downto  80*8), w82 => Pw(113)( 82*8-1 downto  81*8), w83 => Pw(113)( 83*8-1 downto  82*8), w84 => Pw(113)( 84*8-1 downto  83*8), 
w85 => Pw(113)( 85*8-1 downto  84*8), w86 => Pw(113)( 86*8-1 downto  85*8), w87 => Pw(113)( 87*8-1 downto  86*8), w88 => Pw(113)( 88*8-1 downto  87*8), 
w89 => Pw(113)( 89*8-1 downto  88*8), w90 => Pw(113)( 90*8-1 downto  89*8), w91 => Pw(113)( 91*8-1 downto  90*8), w92 => Pw(113)( 92*8-1 downto  91*8), 
w93 => Pw(113)( 93*8-1 downto  92*8), w94 => Pw(113)( 94*8-1 downto  93*8), w95 => Pw(113)( 95*8-1 downto  94*8), w96 => Pw(113)( 96*8-1 downto  95*8), 
w97 => Pw(113)( 97*8-1 downto  96*8), w98 => Pw(113)( 98*8-1 downto  97*8), w99 => Pw(113)( 99*8-1 downto  98*8), w100=> Pw(113)(100*8-1 downto  99*8), 
w101=> Pw(113)(101*8-1 downto 100*8), w102=> Pw(113)(102*8-1 downto 101*8), w103=> Pw(113)(103*8-1 downto 102*8), w104=> Pw(113)(104*8-1 downto 103*8), 
w105=> Pw(113)(105*8-1 downto 104*8), w106=> Pw(113)(106*8-1 downto 105*8), w107=> Pw(113)(107*8-1 downto 106*8), w108=> Pw(113)(108*8-1 downto 107*8), 
w109=> Pw(113)(109*8-1 downto 108*8), w110=> Pw(113)(110*8-1 downto 109*8), w111=> Pw(113)(111*8-1 downto 110*8), w112=> Pw(113)(112*8-1 downto 111*8), 
w113=> Pw(113)(113*8-1 downto 112*8), w114=> Pw(113)(114*8-1 downto 113*8), w115=> Pw(113)(115*8-1 downto 114*8), w116=> Pw(113)(116*8-1 downto 115*8), 
w117=> Pw(113)(117*8-1 downto 116*8), w118=> Pw(113)(118*8-1 downto 117*8), w119=> Pw(113)(119*8-1 downto 118*8), w120=> Pw(113)(120*8-1 downto 119*8), 
w121=> Pw(113)(121*8-1 downto 120*8), w122=> Pw(113)(122*8-1 downto 121*8), w123=> Pw(113)(123*8-1 downto 122*8), w124=> Pw(113)(124*8-1 downto 123*8), 
w125=> Pw(113)(125*8-1 downto 124*8), w126=> Pw(113)(126*8-1 downto 125*8), w127=> Pw(113)(127*8-1 downto 126*8), w128=> Pw(113)(128*8-1 downto 127*8), 
           d_out   => pca_d113_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_114_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(114)(     7 downto    0),   w02 => Pw(114)( 2*8-1 downto    8),   w03 => Pw(114)( 3*8-1 downto  2*8),   w04 => Pw(114)( 4*8-1 downto  3*8),   
w05 => Pw(114)( 5*8-1 downto  4*8),   w06 => Pw(114)( 6*8-1 downto  5*8),   w07 => Pw(114)( 7*8-1 downto  6*8),   w08 => Pw(114)( 8*8-1 downto  7*8),  
w09 => Pw(114)( 9*8-1 downto  8*8),   w10 => Pw(114)(10*8-1 downto  9*8),   w11 => Pw(114)(11*8-1 downto 10*8),   w12 => Pw(114)(12*8-1 downto 11*8),   
w13 => Pw(114)(13*8-1 downto 12*8),   w14 => Pw(114)(14*8-1 downto 13*8),   w15 => Pw(114)(15*8-1 downto 14*8),   w16 => Pw(114)(16*8-1 downto 15*8),  
w17 => Pw(114)(17*8-1 downto 16*8),   w18 => Pw(114)(18*8-1 downto 17*8),   w19 => Pw(114)(19*8-1 downto 18*8),   w20 => Pw(114)(20*8-1 downto 19*8),   
w21 => Pw(114)(21*8-1 downto 20*8),   w22 => Pw(114)(22*8-1 downto 21*8),   w23 => Pw(114)(23*8-1 downto 22*8),   w24 => Pw(114)(24*8-1 downto 23*8),  
w25 => Pw(114)(25*8-1 downto 24*8),   w26 => Pw(114)(26*8-1 downto 25*8),   w27 => Pw(114)(27*8-1 downto 26*8),   w28 => Pw(114)(28*8-1 downto 27*8),   
w29 => Pw(114)(29*8-1 downto 28*8),   w30 => Pw(114)(30*8-1 downto 29*8),   w31 => Pw(114)(31*8-1 downto 30*8),   w32 => Pw(114)(32*8-1 downto 31*8),  
w33 => Pw(114)(33*8-1 downto 32*8),   w34 => Pw(114)(34*8-1 downto 33*8),   w35 => Pw(114)(35*8-1 downto 34*8),   w36 => Pw(114)(36*8-1 downto 35*8),   
w37 => Pw(114)(37*8-1 downto 36*8),   w38 => Pw(114)(38*8-1 downto 37*8),   w39 => Pw(114)(39*8-1 downto 38*8),   w40 => Pw(114)(40*8-1 downto 39*8),  
w41 => Pw(114)(41*8-1 downto 40*8),   w42 => Pw(114)(42*8-1 downto 41*8),   w43 => Pw(114)(43*8-1 downto 42*8),   w44 => Pw(114)(44*8-1 downto 43*8),   
w45 => Pw(114)(45*8-1 downto 44*8),   w46 => Pw(114)(46*8-1 downto 45*8),   w47 => Pw(114)(47*8-1 downto 46*8),   w48 => Pw(114)(48*8-1 downto 47*8),  
w49 => Pw(114)(49*8-1 downto 48*8),   w50 => Pw(114)(50*8-1 downto 49*8),   w51 => Pw(114)(51*8-1 downto 50*8),   w52 => Pw(114)(52*8-1 downto 51*8),   
w53 => Pw(114)(53*8-1 downto 52*8),   w54 => Pw(114)(54*8-1 downto 53*8),   w55 => Pw(114)(55*8-1 downto 54*8),   w56 => Pw(114)(56*8-1 downto 55*8),  
w57 => Pw(114)(57*8-1 downto 56*8),   w58 => Pw(114)(58*8-1 downto 57*8),   w59 => Pw(114)(59*8-1 downto 58*8),   w60 => Pw(114)(60*8-1 downto 59*8),   
w61 => Pw(114)(61*8-1 downto 60*8),   w62 => Pw(114)(62*8-1 downto 61*8),   w63 => Pw(114)(63*8-1 downto 62*8),   w64 => Pw(114)(64*8-1 downto 63*8), 
w65 => Pw(114)( 65*8-1 downto  64*8), w66 => Pw(114)( 66*8-1 downto  65*8), w67 => Pw(114)( 67*8-1 downto  66*8), w68 => Pw(114)( 68*8-1 downto  67*8), 
w69 => Pw(114)( 69*8-1 downto  68*8), w70 => Pw(114)( 70*8-1 downto  69*8), w71 => Pw(114)( 71*8-1 downto  70*8), w72 => Pw(114)( 72*8-1 downto  71*8), 
w73 => Pw(114)( 73*8-1 downto  72*8), w74 => Pw(114)( 74*8-1 downto  73*8), w75 => Pw(114)( 75*8-1 downto  74*8), w76 => Pw(114)( 76*8-1 downto  75*8), 
w77 => Pw(114)( 77*8-1 downto  76*8), w78 => Pw(114)( 78*8-1 downto  77*8), w79 => Pw(114)( 79*8-1 downto  78*8), w80 => Pw(114)( 80*8-1 downto  79*8), 
w81 => Pw(114)( 81*8-1 downto  80*8), w82 => Pw(114)( 82*8-1 downto  81*8), w83 => Pw(114)( 83*8-1 downto  82*8), w84 => Pw(114)( 84*8-1 downto  83*8), 
w85 => Pw(114)( 85*8-1 downto  84*8), w86 => Pw(114)( 86*8-1 downto  85*8), w87 => Pw(114)( 87*8-1 downto  86*8), w88 => Pw(114)( 88*8-1 downto  87*8), 
w89 => Pw(114)( 89*8-1 downto  88*8), w90 => Pw(114)( 90*8-1 downto  89*8), w91 => Pw(114)( 91*8-1 downto  90*8), w92 => Pw(114)( 92*8-1 downto  91*8), 
w93 => Pw(114)( 93*8-1 downto  92*8), w94 => Pw(114)( 94*8-1 downto  93*8), w95 => Pw(114)( 95*8-1 downto  94*8), w96 => Pw(114)( 96*8-1 downto  95*8), 
w97 => Pw(114)( 97*8-1 downto  96*8), w98 => Pw(114)( 98*8-1 downto  97*8), w99 => Pw(114)( 99*8-1 downto  98*8), w100=> Pw(114)(100*8-1 downto  99*8), 
w101=> Pw(114)(101*8-1 downto 100*8), w102=> Pw(114)(102*8-1 downto 101*8), w103=> Pw(114)(103*8-1 downto 102*8), w104=> Pw(114)(104*8-1 downto 103*8), 
w105=> Pw(114)(105*8-1 downto 104*8), w106=> Pw(114)(106*8-1 downto 105*8), w107=> Pw(114)(107*8-1 downto 106*8), w108=> Pw(114)(108*8-1 downto 107*8), 
w109=> Pw(114)(109*8-1 downto 108*8), w110=> Pw(114)(110*8-1 downto 109*8), w111=> Pw(114)(111*8-1 downto 110*8), w112=> Pw(114)(112*8-1 downto 111*8), 
w113=> Pw(114)(113*8-1 downto 112*8), w114=> Pw(114)(114*8-1 downto 113*8), w115=> Pw(114)(115*8-1 downto 114*8), w116=> Pw(114)(116*8-1 downto 115*8), 
w117=> Pw(114)(117*8-1 downto 116*8), w118=> Pw(114)(118*8-1 downto 117*8), w119=> Pw(114)(119*8-1 downto 118*8), w120=> Pw(114)(120*8-1 downto 119*8), 
w121=> Pw(114)(121*8-1 downto 120*8), w122=> Pw(114)(122*8-1 downto 121*8), w123=> Pw(114)(123*8-1 downto 122*8), w124=> Pw(114)(124*8-1 downto 123*8), 
w125=> Pw(114)(125*8-1 downto 124*8), w126=> Pw(114)(126*8-1 downto 125*8), w127=> Pw(114)(127*8-1 downto 126*8), w128=> Pw(114)(128*8-1 downto 127*8), 
           d_out   => pca_d114_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_115_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(115)(     7 downto    0),   w02 => Pw(115)( 2*8-1 downto    8),   w03 => Pw(115)( 3*8-1 downto  2*8),   w04 => Pw(115)( 4*8-1 downto  3*8),   
w05 => Pw(115)( 5*8-1 downto  4*8),   w06 => Pw(115)( 6*8-1 downto  5*8),   w07 => Pw(115)( 7*8-1 downto  6*8),   w08 => Pw(115)( 8*8-1 downto  7*8),  
w09 => Pw(115)( 9*8-1 downto  8*8),   w10 => Pw(115)(10*8-1 downto  9*8),   w11 => Pw(115)(11*8-1 downto 10*8),   w12 => Pw(115)(12*8-1 downto 11*8),   
w13 => Pw(115)(13*8-1 downto 12*8),   w14 => Pw(115)(14*8-1 downto 13*8),   w15 => Pw(115)(15*8-1 downto 14*8),   w16 => Pw(115)(16*8-1 downto 15*8),  
w17 => Pw(115)(17*8-1 downto 16*8),   w18 => Pw(115)(18*8-1 downto 17*8),   w19 => Pw(115)(19*8-1 downto 18*8),   w20 => Pw(115)(20*8-1 downto 19*8),   
w21 => Pw(115)(21*8-1 downto 20*8),   w22 => Pw(115)(22*8-1 downto 21*8),   w23 => Pw(115)(23*8-1 downto 22*8),   w24 => Pw(115)(24*8-1 downto 23*8),  
w25 => Pw(115)(25*8-1 downto 24*8),   w26 => Pw(115)(26*8-1 downto 25*8),   w27 => Pw(115)(27*8-1 downto 26*8),   w28 => Pw(115)(28*8-1 downto 27*8),   
w29 => Pw(115)(29*8-1 downto 28*8),   w30 => Pw(115)(30*8-1 downto 29*8),   w31 => Pw(115)(31*8-1 downto 30*8),   w32 => Pw(115)(32*8-1 downto 31*8),  
w33 => Pw(115)(33*8-1 downto 32*8),   w34 => Pw(115)(34*8-1 downto 33*8),   w35 => Pw(115)(35*8-1 downto 34*8),   w36 => Pw(115)(36*8-1 downto 35*8),   
w37 => Pw(115)(37*8-1 downto 36*8),   w38 => Pw(115)(38*8-1 downto 37*8),   w39 => Pw(115)(39*8-1 downto 38*8),   w40 => Pw(115)(40*8-1 downto 39*8),  
w41 => Pw(115)(41*8-1 downto 40*8),   w42 => Pw(115)(42*8-1 downto 41*8),   w43 => Pw(115)(43*8-1 downto 42*8),   w44 => Pw(115)(44*8-1 downto 43*8),   
w45 => Pw(115)(45*8-1 downto 44*8),   w46 => Pw(115)(46*8-1 downto 45*8),   w47 => Pw(115)(47*8-1 downto 46*8),   w48 => Pw(115)(48*8-1 downto 47*8),  
w49 => Pw(115)(49*8-1 downto 48*8),   w50 => Pw(115)(50*8-1 downto 49*8),   w51 => Pw(115)(51*8-1 downto 50*8),   w52 => Pw(115)(52*8-1 downto 51*8),   
w53 => Pw(115)(53*8-1 downto 52*8),   w54 => Pw(115)(54*8-1 downto 53*8),   w55 => Pw(115)(55*8-1 downto 54*8),   w56 => Pw(115)(56*8-1 downto 55*8),  
w57 => Pw(115)(57*8-1 downto 56*8),   w58 => Pw(115)(58*8-1 downto 57*8),   w59 => Pw(115)(59*8-1 downto 58*8),   w60 => Pw(115)(60*8-1 downto 59*8),   
w61 => Pw(115)(61*8-1 downto 60*8),   w62 => Pw(115)(62*8-1 downto 61*8),   w63 => Pw(115)(63*8-1 downto 62*8),   w64 => Pw(115)(64*8-1 downto 63*8), 
w65 => Pw(115)( 65*8-1 downto  64*8), w66 => Pw(115)( 66*8-1 downto  65*8), w67 => Pw(115)( 67*8-1 downto  66*8), w68 => Pw(115)( 68*8-1 downto  67*8), 
w69 => Pw(115)( 69*8-1 downto  68*8), w70 => Pw(115)( 70*8-1 downto  69*8), w71 => Pw(115)( 71*8-1 downto  70*8), w72 => Pw(115)( 72*8-1 downto  71*8), 
w73 => Pw(115)( 73*8-1 downto  72*8), w74 => Pw(115)( 74*8-1 downto  73*8), w75 => Pw(115)( 75*8-1 downto  74*8), w76 => Pw(115)( 76*8-1 downto  75*8), 
w77 => Pw(115)( 77*8-1 downto  76*8), w78 => Pw(115)( 78*8-1 downto  77*8), w79 => Pw(115)( 79*8-1 downto  78*8), w80 => Pw(115)( 80*8-1 downto  79*8), 
w81 => Pw(115)( 81*8-1 downto  80*8), w82 => Pw(115)( 82*8-1 downto  81*8), w83 => Pw(115)( 83*8-1 downto  82*8), w84 => Pw(115)( 84*8-1 downto  83*8), 
w85 => Pw(115)( 85*8-1 downto  84*8), w86 => Pw(115)( 86*8-1 downto  85*8), w87 => Pw(115)( 87*8-1 downto  86*8), w88 => Pw(115)( 88*8-1 downto  87*8), 
w89 => Pw(115)( 89*8-1 downto  88*8), w90 => Pw(115)( 90*8-1 downto  89*8), w91 => Pw(115)( 91*8-1 downto  90*8), w92 => Pw(115)( 92*8-1 downto  91*8), 
w93 => Pw(115)( 93*8-1 downto  92*8), w94 => Pw(115)( 94*8-1 downto  93*8), w95 => Pw(115)( 95*8-1 downto  94*8), w96 => Pw(115)( 96*8-1 downto  95*8), 
w97 => Pw(115)( 97*8-1 downto  96*8), w98 => Pw(115)( 98*8-1 downto  97*8), w99 => Pw(115)( 99*8-1 downto  98*8), w100=> Pw(115)(100*8-1 downto  99*8), 
w101=> Pw(115)(101*8-1 downto 100*8), w102=> Pw(115)(102*8-1 downto 101*8), w103=> Pw(115)(103*8-1 downto 102*8), w104=> Pw(115)(104*8-1 downto 103*8), 
w105=> Pw(115)(105*8-1 downto 104*8), w106=> Pw(115)(106*8-1 downto 105*8), w107=> Pw(115)(107*8-1 downto 106*8), w108=> Pw(115)(108*8-1 downto 107*8), 
w109=> Pw(115)(109*8-1 downto 108*8), w110=> Pw(115)(110*8-1 downto 109*8), w111=> Pw(115)(111*8-1 downto 110*8), w112=> Pw(115)(112*8-1 downto 111*8), 
w113=> Pw(115)(113*8-1 downto 112*8), w114=> Pw(115)(114*8-1 downto 113*8), w115=> Pw(115)(115*8-1 downto 114*8), w116=> Pw(115)(116*8-1 downto 115*8), 
w117=> Pw(115)(117*8-1 downto 116*8), w118=> Pw(115)(118*8-1 downto 117*8), w119=> Pw(115)(119*8-1 downto 118*8), w120=> Pw(115)(120*8-1 downto 119*8), 
w121=> Pw(115)(121*8-1 downto 120*8), w122=> Pw(115)(122*8-1 downto 121*8), w123=> Pw(115)(123*8-1 downto 122*8), w124=> Pw(115)(124*8-1 downto 123*8), 
w125=> Pw(115)(125*8-1 downto 124*8), w126=> Pw(115)(126*8-1 downto 125*8), w127=> Pw(115)(127*8-1 downto 126*8), w128=> Pw(115)(128*8-1 downto 127*8), 
           d_out   => pca_d115_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_116_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(116)(     7 downto    0),   w02 => Pw(116)( 2*8-1 downto    8),   w03 => Pw(116)( 3*8-1 downto  2*8),   w04 => Pw(116)( 4*8-1 downto  3*8),   
w05 => Pw(116)( 5*8-1 downto  4*8),   w06 => Pw(116)( 6*8-1 downto  5*8),   w07 => Pw(116)( 7*8-1 downto  6*8),   w08 => Pw(116)( 8*8-1 downto  7*8),  
w09 => Pw(116)( 9*8-1 downto  8*8),   w10 => Pw(116)(10*8-1 downto  9*8),   w11 => Pw(116)(11*8-1 downto 10*8),   w12 => Pw(116)(12*8-1 downto 11*8),   
w13 => Pw(116)(13*8-1 downto 12*8),   w14 => Pw(116)(14*8-1 downto 13*8),   w15 => Pw(116)(15*8-1 downto 14*8),   w16 => Pw(116)(16*8-1 downto 15*8),  
w17 => Pw(116)(17*8-1 downto 16*8),   w18 => Pw(116)(18*8-1 downto 17*8),   w19 => Pw(116)(19*8-1 downto 18*8),   w20 => Pw(116)(20*8-1 downto 19*8),   
w21 => Pw(116)(21*8-1 downto 20*8),   w22 => Pw(116)(22*8-1 downto 21*8),   w23 => Pw(116)(23*8-1 downto 22*8),   w24 => Pw(116)(24*8-1 downto 23*8),  
w25 => Pw(116)(25*8-1 downto 24*8),   w26 => Pw(116)(26*8-1 downto 25*8),   w27 => Pw(116)(27*8-1 downto 26*8),   w28 => Pw(116)(28*8-1 downto 27*8),   
w29 => Pw(116)(29*8-1 downto 28*8),   w30 => Pw(116)(30*8-1 downto 29*8),   w31 => Pw(116)(31*8-1 downto 30*8),   w32 => Pw(116)(32*8-1 downto 31*8),  
w33 => Pw(116)(33*8-1 downto 32*8),   w34 => Pw(116)(34*8-1 downto 33*8),   w35 => Pw(116)(35*8-1 downto 34*8),   w36 => Pw(116)(36*8-1 downto 35*8),   
w37 => Pw(116)(37*8-1 downto 36*8),   w38 => Pw(116)(38*8-1 downto 37*8),   w39 => Pw(116)(39*8-1 downto 38*8),   w40 => Pw(116)(40*8-1 downto 39*8),  
w41 => Pw(116)(41*8-1 downto 40*8),   w42 => Pw(116)(42*8-1 downto 41*8),   w43 => Pw(116)(43*8-1 downto 42*8),   w44 => Pw(116)(44*8-1 downto 43*8),   
w45 => Pw(116)(45*8-1 downto 44*8),   w46 => Pw(116)(46*8-1 downto 45*8),   w47 => Pw(116)(47*8-1 downto 46*8),   w48 => Pw(116)(48*8-1 downto 47*8),  
w49 => Pw(116)(49*8-1 downto 48*8),   w50 => Pw(116)(50*8-1 downto 49*8),   w51 => Pw(116)(51*8-1 downto 50*8),   w52 => Pw(116)(52*8-1 downto 51*8),   
w53 => Pw(116)(53*8-1 downto 52*8),   w54 => Pw(116)(54*8-1 downto 53*8),   w55 => Pw(116)(55*8-1 downto 54*8),   w56 => Pw(116)(56*8-1 downto 55*8),  
w57 => Pw(116)(57*8-1 downto 56*8),   w58 => Pw(116)(58*8-1 downto 57*8),   w59 => Pw(116)(59*8-1 downto 58*8),   w60 => Pw(116)(60*8-1 downto 59*8),   
w61 => Pw(116)(61*8-1 downto 60*8),   w62 => Pw(116)(62*8-1 downto 61*8),   w63 => Pw(116)(63*8-1 downto 62*8),   w64 => Pw(116)(64*8-1 downto 63*8), 
w65 => Pw(116)( 65*8-1 downto  64*8), w66 => Pw(116)( 66*8-1 downto  65*8), w67 => Pw(116)( 67*8-1 downto  66*8), w68 => Pw(116)( 68*8-1 downto  67*8), 
w69 => Pw(116)( 69*8-1 downto  68*8), w70 => Pw(116)( 70*8-1 downto  69*8), w71 => Pw(116)( 71*8-1 downto  70*8), w72 => Pw(116)( 72*8-1 downto  71*8), 
w73 => Pw(116)( 73*8-1 downto  72*8), w74 => Pw(116)( 74*8-1 downto  73*8), w75 => Pw(116)( 75*8-1 downto  74*8), w76 => Pw(116)( 76*8-1 downto  75*8), 
w77 => Pw(116)( 77*8-1 downto  76*8), w78 => Pw(116)( 78*8-1 downto  77*8), w79 => Pw(116)( 79*8-1 downto  78*8), w80 => Pw(116)( 80*8-1 downto  79*8), 
w81 => Pw(116)( 81*8-1 downto  80*8), w82 => Pw(116)( 82*8-1 downto  81*8), w83 => Pw(116)( 83*8-1 downto  82*8), w84 => Pw(116)( 84*8-1 downto  83*8), 
w85 => Pw(116)( 85*8-1 downto  84*8), w86 => Pw(116)( 86*8-1 downto  85*8), w87 => Pw(116)( 87*8-1 downto  86*8), w88 => Pw(116)( 88*8-1 downto  87*8), 
w89 => Pw(116)( 89*8-1 downto  88*8), w90 => Pw(116)( 90*8-1 downto  89*8), w91 => Pw(116)( 91*8-1 downto  90*8), w92 => Pw(116)( 92*8-1 downto  91*8), 
w93 => Pw(116)( 93*8-1 downto  92*8), w94 => Pw(116)( 94*8-1 downto  93*8), w95 => Pw(116)( 95*8-1 downto  94*8), w96 => Pw(116)( 96*8-1 downto  95*8), 
w97 => Pw(116)( 97*8-1 downto  96*8), w98 => Pw(116)( 98*8-1 downto  97*8), w99 => Pw(116)( 99*8-1 downto  98*8), w100=> Pw(116)(100*8-1 downto  99*8), 
w101=> Pw(116)(101*8-1 downto 100*8), w102=> Pw(116)(102*8-1 downto 101*8), w103=> Pw(116)(103*8-1 downto 102*8), w104=> Pw(116)(104*8-1 downto 103*8), 
w105=> Pw(116)(105*8-1 downto 104*8), w106=> Pw(116)(106*8-1 downto 105*8), w107=> Pw(116)(107*8-1 downto 106*8), w108=> Pw(116)(108*8-1 downto 107*8), 
w109=> Pw(116)(109*8-1 downto 108*8), w110=> Pw(116)(110*8-1 downto 109*8), w111=> Pw(116)(111*8-1 downto 110*8), w112=> Pw(116)(112*8-1 downto 111*8), 
w113=> Pw(116)(113*8-1 downto 112*8), w114=> Pw(116)(114*8-1 downto 113*8), w115=> Pw(116)(115*8-1 downto 114*8), w116=> Pw(116)(116*8-1 downto 115*8), 
w117=> Pw(116)(117*8-1 downto 116*8), w118=> Pw(116)(118*8-1 downto 117*8), w119=> Pw(116)(119*8-1 downto 118*8), w120=> Pw(116)(120*8-1 downto 119*8), 
w121=> Pw(116)(121*8-1 downto 120*8), w122=> Pw(116)(122*8-1 downto 121*8), w123=> Pw(116)(123*8-1 downto 122*8), w124=> Pw(116)(124*8-1 downto 123*8), 
w125=> Pw(116)(125*8-1 downto 124*8), w126=> Pw(116)(126*8-1 downto 125*8), w127=> Pw(116)(127*8-1 downto 126*8), w128=> Pw(116)(128*8-1 downto 127*8), 
           d_out   => pca_d116_out   ,
           en_out  => open  ,
           sof_out => open );



  PCA128_117_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(117)(     7 downto    0),   w02 => Pw(117)( 2*8-1 downto    8),   w03 => Pw(117)( 3*8-1 downto  2*8),   w04 => Pw(117)( 4*8-1 downto  3*8),   
w05 => Pw(117)( 5*8-1 downto  4*8),   w06 => Pw(117)( 6*8-1 downto  5*8),   w07 => Pw(117)( 7*8-1 downto  6*8),   w08 => Pw(117)( 8*8-1 downto  7*8),  
w09 => Pw(117)( 9*8-1 downto  8*8),   w10 => Pw(117)(10*8-1 downto  9*8),   w11 => Pw(117)(11*8-1 downto 10*8),   w12 => Pw(117)(12*8-1 downto 11*8),   
w13 => Pw(117)(13*8-1 downto 12*8),   w14 => Pw(117)(14*8-1 downto 13*8),   w15 => Pw(117)(15*8-1 downto 14*8),   w16 => Pw(117)(16*8-1 downto 15*8),  
w17 => Pw(117)(17*8-1 downto 16*8),   w18 => Pw(117)(18*8-1 downto 17*8),   w19 => Pw(117)(19*8-1 downto 18*8),   w20 => Pw(117)(20*8-1 downto 19*8),   
w21 => Pw(117)(21*8-1 downto 20*8),   w22 => Pw(117)(22*8-1 downto 21*8),   w23 => Pw(117)(23*8-1 downto 22*8),   w24 => Pw(117)(24*8-1 downto 23*8),  
w25 => Pw(117)(25*8-1 downto 24*8),   w26 => Pw(117)(26*8-1 downto 25*8),   w27 => Pw(117)(27*8-1 downto 26*8),   w28 => Pw(117)(28*8-1 downto 27*8),   
w29 => Pw(117)(29*8-1 downto 28*8),   w30 => Pw(117)(30*8-1 downto 29*8),   w31 => Pw(117)(31*8-1 downto 30*8),   w32 => Pw(117)(32*8-1 downto 31*8),  
w33 => Pw(117)(33*8-1 downto 32*8),   w34 => Pw(117)(34*8-1 downto 33*8),   w35 => Pw(117)(35*8-1 downto 34*8),   w36 => Pw(117)(36*8-1 downto 35*8),   
w37 => Pw(117)(37*8-1 downto 36*8),   w38 => Pw(117)(38*8-1 downto 37*8),   w39 => Pw(117)(39*8-1 downto 38*8),   w40 => Pw(117)(40*8-1 downto 39*8),  
w41 => Pw(117)(41*8-1 downto 40*8),   w42 => Pw(117)(42*8-1 downto 41*8),   w43 => Pw(117)(43*8-1 downto 42*8),   w44 => Pw(117)(44*8-1 downto 43*8),   
w45 => Pw(117)(45*8-1 downto 44*8),   w46 => Pw(117)(46*8-1 downto 45*8),   w47 => Pw(117)(47*8-1 downto 46*8),   w48 => Pw(117)(48*8-1 downto 47*8),  
w49 => Pw(117)(49*8-1 downto 48*8),   w50 => Pw(117)(50*8-1 downto 49*8),   w51 => Pw(117)(51*8-1 downto 50*8),   w52 => Pw(117)(52*8-1 downto 51*8),   
w53 => Pw(117)(53*8-1 downto 52*8),   w54 => Pw(117)(54*8-1 downto 53*8),   w55 => Pw(117)(55*8-1 downto 54*8),   w56 => Pw(117)(56*8-1 downto 55*8),  
w57 => Pw(117)(57*8-1 downto 56*8),   w58 => Pw(117)(58*8-1 downto 57*8),   w59 => Pw(117)(59*8-1 downto 58*8),   w60 => Pw(117)(60*8-1 downto 59*8),   
w61 => Pw(117)(61*8-1 downto 60*8),   w62 => Pw(117)(62*8-1 downto 61*8),   w63 => Pw(117)(63*8-1 downto 62*8),   w64 => Pw(117)(64*8-1 downto 63*8), 
w65 => Pw(117)( 65*8-1 downto  64*8), w66 => Pw(117)( 66*8-1 downto  65*8), w67 => Pw(117)( 67*8-1 downto  66*8), w68 => Pw(117)( 68*8-1 downto  67*8), 
w69 => Pw(117)( 69*8-1 downto  68*8), w70 => Pw(117)( 70*8-1 downto  69*8), w71 => Pw(117)( 71*8-1 downto  70*8), w72 => Pw(117)( 72*8-1 downto  71*8), 
w73 => Pw(117)( 73*8-1 downto  72*8), w74 => Pw(117)( 74*8-1 downto  73*8), w75 => Pw(117)( 75*8-1 downto  74*8), w76 => Pw(117)( 76*8-1 downto  75*8), 
w77 => Pw(117)( 77*8-1 downto  76*8), w78 => Pw(117)( 78*8-1 downto  77*8), w79 => Pw(117)( 79*8-1 downto  78*8), w80 => Pw(117)( 80*8-1 downto  79*8), 
w81 => Pw(117)( 81*8-1 downto  80*8), w82 => Pw(117)( 82*8-1 downto  81*8), w83 => Pw(117)( 83*8-1 downto  82*8), w84 => Pw(117)( 84*8-1 downto  83*8), 
w85 => Pw(117)( 85*8-1 downto  84*8), w86 => Pw(117)( 86*8-1 downto  85*8), w87 => Pw(117)( 87*8-1 downto  86*8), w88 => Pw(117)( 88*8-1 downto  87*8), 
w89 => Pw(117)( 89*8-1 downto  88*8), w90 => Pw(117)( 90*8-1 downto  89*8), w91 => Pw(117)( 91*8-1 downto  90*8), w92 => Pw(117)( 92*8-1 downto  91*8), 
w93 => Pw(117)( 93*8-1 downto  92*8), w94 => Pw(117)( 94*8-1 downto  93*8), w95 => Pw(117)( 95*8-1 downto  94*8), w96 => Pw(117)( 96*8-1 downto  95*8), 
w97 => Pw(117)( 97*8-1 downto  96*8), w98 => Pw(117)( 98*8-1 downto  97*8), w99 => Pw(117)( 99*8-1 downto  98*8), w100=> Pw(117)(100*8-1 downto  99*8), 
w101=> Pw(117)(101*8-1 downto 100*8), w102=> Pw(117)(102*8-1 downto 101*8), w103=> Pw(117)(103*8-1 downto 102*8), w104=> Pw(117)(104*8-1 downto 103*8), 
w105=> Pw(117)(105*8-1 downto 104*8), w106=> Pw(117)(106*8-1 downto 105*8), w107=> Pw(117)(107*8-1 downto 106*8), w108=> Pw(117)(108*8-1 downto 107*8), 
w109=> Pw(117)(109*8-1 downto 108*8), w110=> Pw(117)(110*8-1 downto 109*8), w111=> Pw(117)(111*8-1 downto 110*8), w112=> Pw(117)(112*8-1 downto 111*8), 
w113=> Pw(117)(113*8-1 downto 112*8), w114=> Pw(117)(114*8-1 downto 113*8), w115=> Pw(117)(115*8-1 downto 114*8), w116=> Pw(117)(116*8-1 downto 115*8), 
w117=> Pw(117)(117*8-1 downto 116*8), w118=> Pw(117)(118*8-1 downto 117*8), w119=> Pw(117)(119*8-1 downto 118*8), w120=> Pw(117)(120*8-1 downto 119*8), 
w121=> Pw(117)(121*8-1 downto 120*8), w122=> Pw(117)(122*8-1 downto 121*8), w123=> Pw(117)(123*8-1 downto 122*8), w124=> Pw(117)(124*8-1 downto 123*8), 
w125=> Pw(117)(125*8-1 downto 124*8), w126=> Pw(117)(126*8-1 downto 125*8), w127=> Pw(117)(127*8-1 downto 126*8), w128=> Pw(117)(128*8-1 downto 127*8), 
           d_out   => pca_d117_out   ,
           en_out  => open  ,
           sof_out => open );





  PCA128_118_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(118)(     7 downto    0),   w02 => Pw(118)( 2*8-1 downto    8),   w03 => Pw(118)( 3*8-1 downto  2*8),   w04 => Pw(118)( 4*8-1 downto  3*8),   
w05 => Pw(118)( 5*8-1 downto  4*8),   w06 => Pw(118)( 6*8-1 downto  5*8),   w07 => Pw(118)( 7*8-1 downto  6*8),   w08 => Pw(118)( 8*8-1 downto  7*8),  
w09 => Pw(118)( 9*8-1 downto  8*8),   w10 => Pw(118)(10*8-1 downto  9*8),   w11 => Pw(118)(11*8-1 downto 10*8),   w12 => Pw(118)(12*8-1 downto 11*8),   
w13 => Pw(118)(13*8-1 downto 12*8),   w14 => Pw(118)(14*8-1 downto 13*8),   w15 => Pw(118)(15*8-1 downto 14*8),   w16 => Pw(118)(16*8-1 downto 15*8),  
w17 => Pw(118)(17*8-1 downto 16*8),   w18 => Pw(118)(18*8-1 downto 17*8),   w19 => Pw(118)(19*8-1 downto 18*8),   w20 => Pw(118)(20*8-1 downto 19*8),   
w21 => Pw(118)(21*8-1 downto 20*8),   w22 => Pw(118)(22*8-1 downto 21*8),   w23 => Pw(118)(23*8-1 downto 22*8),   w24 => Pw(118)(24*8-1 downto 23*8),  
w25 => Pw(118)(25*8-1 downto 24*8),   w26 => Pw(118)(26*8-1 downto 25*8),   w27 => Pw(118)(27*8-1 downto 26*8),   w28 => Pw(118)(28*8-1 downto 27*8),   
w29 => Pw(118)(29*8-1 downto 28*8),   w30 => Pw(118)(30*8-1 downto 29*8),   w31 => Pw(118)(31*8-1 downto 30*8),   w32 => Pw(118)(32*8-1 downto 31*8),  
w33 => Pw(118)(33*8-1 downto 32*8),   w34 => Pw(118)(34*8-1 downto 33*8),   w35 => Pw(118)(35*8-1 downto 34*8),   w36 => Pw(118)(36*8-1 downto 35*8),   
w37 => Pw(118)(37*8-1 downto 36*8),   w38 => Pw(118)(38*8-1 downto 37*8),   w39 => Pw(118)(39*8-1 downto 38*8),   w40 => Pw(118)(40*8-1 downto 39*8),  
w41 => Pw(118)(41*8-1 downto 40*8),   w42 => Pw(118)(42*8-1 downto 41*8),   w43 => Pw(118)(43*8-1 downto 42*8),   w44 => Pw(118)(44*8-1 downto 43*8),   
w45 => Pw(118)(45*8-1 downto 44*8),   w46 => Pw(118)(46*8-1 downto 45*8),   w47 => Pw(118)(47*8-1 downto 46*8),   w48 => Pw(118)(48*8-1 downto 47*8),  
w49 => Pw(118)(49*8-1 downto 48*8),   w50 => Pw(118)(50*8-1 downto 49*8),   w51 => Pw(118)(51*8-1 downto 50*8),   w52 => Pw(118)(52*8-1 downto 51*8),   
w53 => Pw(118)(53*8-1 downto 52*8),   w54 => Pw(118)(54*8-1 downto 53*8),   w55 => Pw(118)(55*8-1 downto 54*8),   w56 => Pw(118)(56*8-1 downto 55*8),  
w57 => Pw(118)(57*8-1 downto 56*8),   w58 => Pw(118)(58*8-1 downto 57*8),   w59 => Pw(118)(59*8-1 downto 58*8),   w60 => Pw(118)(60*8-1 downto 59*8),   
w61 => Pw(118)(61*8-1 downto 60*8),   w62 => Pw(118)(62*8-1 downto 61*8),   w63 => Pw(118)(63*8-1 downto 62*8),   w64 => Pw(118)(64*8-1 downto 63*8), 
w65 => Pw(118)( 65*8-1 downto  64*8), w66 => Pw(118)( 66*8-1 downto  65*8), w67 => Pw(118)( 67*8-1 downto  66*8), w68 => Pw(118)( 68*8-1 downto  67*8), 
w69 => Pw(118)( 69*8-1 downto  68*8), w70 => Pw(118)( 70*8-1 downto  69*8), w71 => Pw(118)( 71*8-1 downto  70*8), w72 => Pw(118)( 72*8-1 downto  71*8), 
w73 => Pw(118)( 73*8-1 downto  72*8), w74 => Pw(118)( 74*8-1 downto  73*8), w75 => Pw(118)( 75*8-1 downto  74*8), w76 => Pw(118)( 76*8-1 downto  75*8), 
w77 => Pw(118)( 77*8-1 downto  76*8), w78 => Pw(118)( 78*8-1 downto  77*8), w79 => Pw(118)( 79*8-1 downto  78*8), w80 => Pw(118)( 80*8-1 downto  79*8), 
w81 => Pw(118)( 81*8-1 downto  80*8), w82 => Pw(118)( 82*8-1 downto  81*8), w83 => Pw(118)( 83*8-1 downto  82*8), w84 => Pw(118)( 84*8-1 downto  83*8), 
w85 => Pw(118)( 85*8-1 downto  84*8), w86 => Pw(118)( 86*8-1 downto  85*8), w87 => Pw(118)( 87*8-1 downto  86*8), w88 => Pw(118)( 88*8-1 downto  87*8), 
w89 => Pw(118)( 89*8-1 downto  88*8), w90 => Pw(118)( 90*8-1 downto  89*8), w91 => Pw(118)( 91*8-1 downto  90*8), w92 => Pw(118)( 92*8-1 downto  91*8), 
w93 => Pw(118)( 93*8-1 downto  92*8), w94 => Pw(118)( 94*8-1 downto  93*8), w95 => Pw(118)( 95*8-1 downto  94*8), w96 => Pw(118)( 96*8-1 downto  95*8), 
w97 => Pw(118)( 97*8-1 downto  96*8), w98 => Pw(118)( 98*8-1 downto  97*8), w99 => Pw(118)( 99*8-1 downto  98*8), w100=> Pw(118)(100*8-1 downto  99*8), 
w101=> Pw(118)(101*8-1 downto 100*8), w102=> Pw(118)(102*8-1 downto 101*8), w103=> Pw(118)(103*8-1 downto 102*8), w104=> Pw(118)(104*8-1 downto 103*8), 
w105=> Pw(118)(105*8-1 downto 104*8), w106=> Pw(118)(106*8-1 downto 105*8), w107=> Pw(118)(107*8-1 downto 106*8), w108=> Pw(118)(108*8-1 downto 107*8), 
w109=> Pw(118)(109*8-1 downto 108*8), w110=> Pw(118)(110*8-1 downto 109*8), w111=> Pw(118)(111*8-1 downto 110*8), w112=> Pw(118)(112*8-1 downto 111*8), 
w113=> Pw(118)(113*8-1 downto 112*8), w114=> Pw(118)(114*8-1 downto 113*8), w115=> Pw(118)(115*8-1 downto 114*8), w116=> Pw(118)(116*8-1 downto 115*8), 
w117=> Pw(118)(117*8-1 downto 116*8), w118=> Pw(118)(118*8-1 downto 117*8), w119=> Pw(118)(119*8-1 downto 118*8), w120=> Pw(118)(120*8-1 downto 119*8), 
w121=> Pw(118)(121*8-1 downto 120*8), w122=> Pw(118)(122*8-1 downto 121*8), w123=> Pw(118)(123*8-1 downto 122*8), w124=> Pw(118)(124*8-1 downto 123*8), 
w125=> Pw(118)(125*8-1 downto 124*8), w126=> Pw(118)(126*8-1 downto 125*8), w127=> Pw(118)(127*8-1 downto 126*8), w128=> Pw(118)(128*8-1 downto 127*8), 
           d_out   => pca_d118_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_119_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(119)(     7 downto    0),   w02 => Pw(119)( 2*8-1 downto    8),   w03 => Pw(119)( 3*8-1 downto  2*8),   w04 => Pw(119)( 4*8-1 downto  3*8),   
w05 => Pw(119)( 5*8-1 downto  4*8),   w06 => Pw(119)( 6*8-1 downto  5*8),   w07 => Pw(119)( 7*8-1 downto  6*8),   w08 => Pw(119)( 8*8-1 downto  7*8),  
w09 => Pw(119)( 9*8-1 downto  8*8),   w10 => Pw(119)(10*8-1 downto  9*8),   w11 => Pw(119)(11*8-1 downto 10*8),   w12 => Pw(119)(12*8-1 downto 11*8),   
w13 => Pw(119)(13*8-1 downto 12*8),   w14 => Pw(119)(14*8-1 downto 13*8),   w15 => Pw(119)(15*8-1 downto 14*8),   w16 => Pw(119)(16*8-1 downto 15*8),  
w17 => Pw(119)(17*8-1 downto 16*8),   w18 => Pw(119)(18*8-1 downto 17*8),   w19 => Pw(119)(19*8-1 downto 18*8),   w20 => Pw(119)(20*8-1 downto 19*8),   
w21 => Pw(119)(21*8-1 downto 20*8),   w22 => Pw(119)(22*8-1 downto 21*8),   w23 => Pw(119)(23*8-1 downto 22*8),   w24 => Pw(119)(24*8-1 downto 23*8),  
w25 => Pw(119)(25*8-1 downto 24*8),   w26 => Pw(119)(26*8-1 downto 25*8),   w27 => Pw(119)(27*8-1 downto 26*8),   w28 => Pw(119)(28*8-1 downto 27*8),   
w29 => Pw(119)(29*8-1 downto 28*8),   w30 => Pw(119)(30*8-1 downto 29*8),   w31 => Pw(119)(31*8-1 downto 30*8),   w32 => Pw(119)(32*8-1 downto 31*8),  
w33 => Pw(119)(33*8-1 downto 32*8),   w34 => Pw(119)(34*8-1 downto 33*8),   w35 => Pw(119)(35*8-1 downto 34*8),   w36 => Pw(119)(36*8-1 downto 35*8),   
w37 => Pw(119)(37*8-1 downto 36*8),   w38 => Pw(119)(38*8-1 downto 37*8),   w39 => Pw(119)(39*8-1 downto 38*8),   w40 => Pw(119)(40*8-1 downto 39*8),  
w41 => Pw(119)(41*8-1 downto 40*8),   w42 => Pw(119)(42*8-1 downto 41*8),   w43 => Pw(119)(43*8-1 downto 42*8),   w44 => Pw(119)(44*8-1 downto 43*8),   
w45 => Pw(119)(45*8-1 downto 44*8),   w46 => Pw(119)(46*8-1 downto 45*8),   w47 => Pw(119)(47*8-1 downto 46*8),   w48 => Pw(119)(48*8-1 downto 47*8),  
w49 => Pw(119)(49*8-1 downto 48*8),   w50 => Pw(119)(50*8-1 downto 49*8),   w51 => Pw(119)(51*8-1 downto 50*8),   w52 => Pw(119)(52*8-1 downto 51*8),   
w53 => Pw(119)(53*8-1 downto 52*8),   w54 => Pw(119)(54*8-1 downto 53*8),   w55 => Pw(119)(55*8-1 downto 54*8),   w56 => Pw(119)(56*8-1 downto 55*8),  
w57 => Pw(119)(57*8-1 downto 56*8),   w58 => Pw(119)(58*8-1 downto 57*8),   w59 => Pw(119)(59*8-1 downto 58*8),   w60 => Pw(119)(60*8-1 downto 59*8),   
w61 => Pw(119)(61*8-1 downto 60*8),   w62 => Pw(119)(62*8-1 downto 61*8),   w63 => Pw(119)(63*8-1 downto 62*8),   w64 => Pw(119)(64*8-1 downto 63*8), 
w65 => Pw(119)( 65*8-1 downto  64*8), w66 => Pw(119)( 66*8-1 downto  65*8), w67 => Pw(119)( 67*8-1 downto  66*8), w68 => Pw(119)( 68*8-1 downto  67*8), 
w69 => Pw(119)( 69*8-1 downto  68*8), w70 => Pw(119)( 70*8-1 downto  69*8), w71 => Pw(119)( 71*8-1 downto  70*8), w72 => Pw(119)( 72*8-1 downto  71*8), 
w73 => Pw(119)( 73*8-1 downto  72*8), w74 => Pw(119)( 74*8-1 downto  73*8), w75 => Pw(119)( 75*8-1 downto  74*8), w76 => Pw(119)( 76*8-1 downto  75*8), 
w77 => Pw(119)( 77*8-1 downto  76*8), w78 => Pw(119)( 78*8-1 downto  77*8), w79 => Pw(119)( 79*8-1 downto  78*8), w80 => Pw(119)( 80*8-1 downto  79*8), 
w81 => Pw(119)( 81*8-1 downto  80*8), w82 => Pw(119)( 82*8-1 downto  81*8), w83 => Pw(119)( 83*8-1 downto  82*8), w84 => Pw(119)( 84*8-1 downto  83*8), 
w85 => Pw(119)( 85*8-1 downto  84*8), w86 => Pw(119)( 86*8-1 downto  85*8), w87 => Pw(119)( 87*8-1 downto  86*8), w88 => Pw(119)( 88*8-1 downto  87*8), 
w89 => Pw(119)( 89*8-1 downto  88*8), w90 => Pw(119)( 90*8-1 downto  89*8), w91 => Pw(119)( 91*8-1 downto  90*8), w92 => Pw(119)( 92*8-1 downto  91*8), 
w93 => Pw(119)( 93*8-1 downto  92*8), w94 => Pw(119)( 94*8-1 downto  93*8), w95 => Pw(119)( 95*8-1 downto  94*8), w96 => Pw(119)( 96*8-1 downto  95*8), 
w97 => Pw(119)( 97*8-1 downto  96*8), w98 => Pw(119)( 98*8-1 downto  97*8), w99 => Pw(119)( 99*8-1 downto  98*8), w100=> Pw(119)(100*8-1 downto  99*8), 
w101=> Pw(119)(101*8-1 downto 100*8), w102=> Pw(119)(102*8-1 downto 101*8), w103=> Pw(119)(103*8-1 downto 102*8), w104=> Pw(119)(104*8-1 downto 103*8), 
w105=> Pw(119)(105*8-1 downto 104*8), w106=> Pw(119)(106*8-1 downto 105*8), w107=> Pw(119)(107*8-1 downto 106*8), w108=> Pw(119)(108*8-1 downto 107*8), 
w109=> Pw(119)(109*8-1 downto 108*8), w110=> Pw(119)(110*8-1 downto 109*8), w111=> Pw(119)(111*8-1 downto 110*8), w112=> Pw(119)(112*8-1 downto 111*8), 
w113=> Pw(119)(113*8-1 downto 112*8), w114=> Pw(119)(114*8-1 downto 113*8), w115=> Pw(119)(115*8-1 downto 114*8), w116=> Pw(119)(116*8-1 downto 115*8), 
w117=> Pw(119)(117*8-1 downto 116*8), w118=> Pw(119)(118*8-1 downto 117*8), w119=> Pw(119)(119*8-1 downto 118*8), w120=> Pw(119)(120*8-1 downto 119*8), 
w121=> Pw(119)(121*8-1 downto 120*8), w122=> Pw(119)(122*8-1 downto 121*8), w123=> Pw(119)(123*8-1 downto 122*8), w124=> Pw(119)(124*8-1 downto 123*8), 
w125=> Pw(119)(125*8-1 downto 124*8), w126=> Pw(119)(126*8-1 downto 125*8), w127=> Pw(119)(127*8-1 downto 126*8), w128=> Pw(119)(128*8-1 downto 127*8), 
           d_out   => pca_d119_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_120_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(120)(     7 downto    0),   w02 => Pw(120)( 2*8-1 downto    8),   w03 => Pw(120)( 3*8-1 downto  2*8),   w04 => Pw(120)( 4*8-1 downto  3*8),   
w05 => Pw(120)( 5*8-1 downto  4*8),   w06 => Pw(120)( 6*8-1 downto  5*8),   w07 => Pw(120)( 7*8-1 downto  6*8),   w08 => Pw(120)( 8*8-1 downto  7*8),  
w09 => Pw(120)( 9*8-1 downto  8*8),   w10 => Pw(120)(10*8-1 downto  9*8),   w11 => Pw(120)(11*8-1 downto 10*8),   w12 => Pw(120)(12*8-1 downto 11*8),   
w13 => Pw(120)(13*8-1 downto 12*8),   w14 => Pw(120)(14*8-1 downto 13*8),   w15 => Pw(120)(15*8-1 downto 14*8),   w16 => Pw(120)(16*8-1 downto 15*8),  
w17 => Pw(120)(17*8-1 downto 16*8),   w18 => Pw(120)(18*8-1 downto 17*8),   w19 => Pw(120)(19*8-1 downto 18*8),   w20 => Pw(120)(20*8-1 downto 19*8),   
w21 => Pw(120)(21*8-1 downto 20*8),   w22 => Pw(120)(22*8-1 downto 21*8),   w23 => Pw(120)(23*8-1 downto 22*8),   w24 => Pw(120)(24*8-1 downto 23*8),  
w25 => Pw(120)(25*8-1 downto 24*8),   w26 => Pw(120)(26*8-1 downto 25*8),   w27 => Pw(120)(27*8-1 downto 26*8),   w28 => Pw(120)(28*8-1 downto 27*8),   
w29 => Pw(120)(29*8-1 downto 28*8),   w30 => Pw(120)(30*8-1 downto 29*8),   w31 => Pw(120)(31*8-1 downto 30*8),   w32 => Pw(120)(32*8-1 downto 31*8),  
w33 => Pw(120)(33*8-1 downto 32*8),   w34 => Pw(120)(34*8-1 downto 33*8),   w35 => Pw(120)(35*8-1 downto 34*8),   w36 => Pw(120)(36*8-1 downto 35*8),   
w37 => Pw(120)(37*8-1 downto 36*8),   w38 => Pw(120)(38*8-1 downto 37*8),   w39 => Pw(120)(39*8-1 downto 38*8),   w40 => Pw(120)(40*8-1 downto 39*8),  
w41 => Pw(120)(41*8-1 downto 40*8),   w42 => Pw(120)(42*8-1 downto 41*8),   w43 => Pw(120)(43*8-1 downto 42*8),   w44 => Pw(120)(44*8-1 downto 43*8),   
w45 => Pw(120)(45*8-1 downto 44*8),   w46 => Pw(120)(46*8-1 downto 45*8),   w47 => Pw(120)(47*8-1 downto 46*8),   w48 => Pw(120)(48*8-1 downto 47*8),  
w49 => Pw(120)(49*8-1 downto 48*8),   w50 => Pw(120)(50*8-1 downto 49*8),   w51 => Pw(120)(51*8-1 downto 50*8),   w52 => Pw(120)(52*8-1 downto 51*8),   
w53 => Pw(120)(53*8-1 downto 52*8),   w54 => Pw(120)(54*8-1 downto 53*8),   w55 => Pw(120)(55*8-1 downto 54*8),   w56 => Pw(120)(56*8-1 downto 55*8),  
w57 => Pw(120)(57*8-1 downto 56*8),   w58 => Pw(120)(58*8-1 downto 57*8),   w59 => Pw(120)(59*8-1 downto 58*8),   w60 => Pw(120)(60*8-1 downto 59*8),   
w61 => Pw(120)(61*8-1 downto 60*8),   w62 => Pw(120)(62*8-1 downto 61*8),   w63 => Pw(120)(63*8-1 downto 62*8),   w64 => Pw(120)(64*8-1 downto 63*8), 
w65 => Pw(120)( 65*8-1 downto  64*8), w66 => Pw(120)( 66*8-1 downto  65*8), w67 => Pw(120)( 67*8-1 downto  66*8), w68 => Pw(120)( 68*8-1 downto  67*8), 
w69 => Pw(120)( 69*8-1 downto  68*8), w70 => Pw(120)( 70*8-1 downto  69*8), w71 => Pw(120)( 71*8-1 downto  70*8), w72 => Pw(120)( 72*8-1 downto  71*8), 
w73 => Pw(120)( 73*8-1 downto  72*8), w74 => Pw(120)( 74*8-1 downto  73*8), w75 => Pw(120)( 75*8-1 downto  74*8), w76 => Pw(120)( 76*8-1 downto  75*8), 
w77 => Pw(120)( 77*8-1 downto  76*8), w78 => Pw(120)( 78*8-1 downto  77*8), w79 => Pw(120)( 79*8-1 downto  78*8), w80 => Pw(120)( 80*8-1 downto  79*8), 
w81 => Pw(120)( 81*8-1 downto  80*8), w82 => Pw(120)( 82*8-1 downto  81*8), w83 => Pw(120)( 83*8-1 downto  82*8), w84 => Pw(120)( 84*8-1 downto  83*8), 
w85 => Pw(120)( 85*8-1 downto  84*8), w86 => Pw(120)( 86*8-1 downto  85*8), w87 => Pw(120)( 87*8-1 downto  86*8), w88 => Pw(120)( 88*8-1 downto  87*8), 
w89 => Pw(120)( 89*8-1 downto  88*8), w90 => Pw(120)( 90*8-1 downto  89*8), w91 => Pw(120)( 91*8-1 downto  90*8), w92 => Pw(120)( 92*8-1 downto  91*8), 
w93 => Pw(120)( 93*8-1 downto  92*8), w94 => Pw(120)( 94*8-1 downto  93*8), w95 => Pw(120)( 95*8-1 downto  94*8), w96 => Pw(120)( 96*8-1 downto  95*8), 
w97 => Pw(120)( 97*8-1 downto  96*8), w98 => Pw(120)( 98*8-1 downto  97*8), w99 => Pw(120)( 99*8-1 downto  98*8), w100=> Pw(120)(100*8-1 downto  99*8), 
w101=> Pw(120)(101*8-1 downto 100*8), w102=> Pw(120)(102*8-1 downto 101*8), w103=> Pw(120)(103*8-1 downto 102*8), w104=> Pw(120)(104*8-1 downto 103*8), 
w105=> Pw(120)(105*8-1 downto 104*8), w106=> Pw(120)(106*8-1 downto 105*8), w107=> Pw(120)(107*8-1 downto 106*8), w108=> Pw(120)(108*8-1 downto 107*8), 
w109=> Pw(120)(109*8-1 downto 108*8), w110=> Pw(120)(110*8-1 downto 109*8), w111=> Pw(120)(111*8-1 downto 110*8), w112=> Pw(120)(112*8-1 downto 111*8), 
w113=> Pw(120)(113*8-1 downto 112*8), w114=> Pw(120)(114*8-1 downto 113*8), w115=> Pw(120)(115*8-1 downto 114*8), w116=> Pw(120)(116*8-1 downto 115*8), 
w117=> Pw(120)(117*8-1 downto 116*8), w118=> Pw(120)(118*8-1 downto 117*8), w119=> Pw(120)(119*8-1 downto 118*8), w120=> Pw(120)(120*8-1 downto 119*8), 
w121=> Pw(120)(121*8-1 downto 120*8), w122=> Pw(120)(122*8-1 downto 121*8), w123=> Pw(120)(123*8-1 downto 122*8), w124=> Pw(120)(124*8-1 downto 123*8), 
w125=> Pw(120)(125*8-1 downto 124*8), w126=> Pw(120)(126*8-1 downto 125*8), w127=> Pw(120)(127*8-1 downto 126*8), w128=> Pw(120)(128*8-1 downto 127*8), 
           d_out   => pca_d120_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_121_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(121)(     7 downto    0),   w02 => Pw(121)( 2*8-1 downto    8),   w03 => Pw(121)( 3*8-1 downto  2*8),   w04 => Pw(121)( 4*8-1 downto  3*8),   
w05 => Pw(121)( 5*8-1 downto  4*8),   w06 => Pw(121)( 6*8-1 downto  5*8),   w07 => Pw(121)( 7*8-1 downto  6*8),   w08 => Pw(121)( 8*8-1 downto  7*8),  
w09 => Pw(121)( 9*8-1 downto  8*8),   w10 => Pw(121)(10*8-1 downto  9*8),   w11 => Pw(121)(11*8-1 downto 10*8),   w12 => Pw(121)(12*8-1 downto 11*8),   
w13 => Pw(121)(13*8-1 downto 12*8),   w14 => Pw(121)(14*8-1 downto 13*8),   w15 => Pw(121)(15*8-1 downto 14*8),   w16 => Pw(121)(16*8-1 downto 15*8),  
w17 => Pw(121)(17*8-1 downto 16*8),   w18 => Pw(121)(18*8-1 downto 17*8),   w19 => Pw(121)(19*8-1 downto 18*8),   w20 => Pw(121)(20*8-1 downto 19*8),   
w21 => Pw(121)(21*8-1 downto 20*8),   w22 => Pw(121)(22*8-1 downto 21*8),   w23 => Pw(121)(23*8-1 downto 22*8),   w24 => Pw(121)(24*8-1 downto 23*8),  
w25 => Pw(121)(25*8-1 downto 24*8),   w26 => Pw(121)(26*8-1 downto 25*8),   w27 => Pw(121)(27*8-1 downto 26*8),   w28 => Pw(121)(28*8-1 downto 27*8),   
w29 => Pw(121)(29*8-1 downto 28*8),   w30 => Pw(121)(30*8-1 downto 29*8),   w31 => Pw(121)(31*8-1 downto 30*8),   w32 => Pw(121)(32*8-1 downto 31*8),  
w33 => Pw(121)(33*8-1 downto 32*8),   w34 => Pw(121)(34*8-1 downto 33*8),   w35 => Pw(121)(35*8-1 downto 34*8),   w36 => Pw(121)(36*8-1 downto 35*8),   
w37 => Pw(121)(37*8-1 downto 36*8),   w38 => Pw(121)(38*8-1 downto 37*8),   w39 => Pw(121)(39*8-1 downto 38*8),   w40 => Pw(121)(40*8-1 downto 39*8),  
w41 => Pw(121)(41*8-1 downto 40*8),   w42 => Pw(121)(42*8-1 downto 41*8),   w43 => Pw(121)(43*8-1 downto 42*8),   w44 => Pw(121)(44*8-1 downto 43*8),   
w45 => Pw(121)(45*8-1 downto 44*8),   w46 => Pw(121)(46*8-1 downto 45*8),   w47 => Pw(121)(47*8-1 downto 46*8),   w48 => Pw(121)(48*8-1 downto 47*8),  
w49 => Pw(121)(49*8-1 downto 48*8),   w50 => Pw(121)(50*8-1 downto 49*8),   w51 => Pw(121)(51*8-1 downto 50*8),   w52 => Pw(121)(52*8-1 downto 51*8),   
w53 => Pw(121)(53*8-1 downto 52*8),   w54 => Pw(121)(54*8-1 downto 53*8),   w55 => Pw(121)(55*8-1 downto 54*8),   w56 => Pw(121)(56*8-1 downto 55*8),  
w57 => Pw(121)(57*8-1 downto 56*8),   w58 => Pw(121)(58*8-1 downto 57*8),   w59 => Pw(121)(59*8-1 downto 58*8),   w60 => Pw(121)(60*8-1 downto 59*8),   
w61 => Pw(121)(61*8-1 downto 60*8),   w62 => Pw(121)(62*8-1 downto 61*8),   w63 => Pw(121)(63*8-1 downto 62*8),   w64 => Pw(121)(64*8-1 downto 63*8), 
w65 => Pw(121)( 65*8-1 downto  64*8), w66 => Pw(121)( 66*8-1 downto  65*8), w67 => Pw(121)( 67*8-1 downto  66*8), w68 => Pw(121)( 68*8-1 downto  67*8), 
w69 => Pw(121)( 69*8-1 downto  68*8), w70 => Pw(121)( 70*8-1 downto  69*8), w71 => Pw(121)( 71*8-1 downto  70*8), w72 => Pw(121)( 72*8-1 downto  71*8), 
w73 => Pw(121)( 73*8-1 downto  72*8), w74 => Pw(121)( 74*8-1 downto  73*8), w75 => Pw(121)( 75*8-1 downto  74*8), w76 => Pw(121)( 76*8-1 downto  75*8), 
w77 => Pw(121)( 77*8-1 downto  76*8), w78 => Pw(121)( 78*8-1 downto  77*8), w79 => Pw(121)( 79*8-1 downto  78*8), w80 => Pw(121)( 80*8-1 downto  79*8), 
w81 => Pw(121)( 81*8-1 downto  80*8), w82 => Pw(121)( 82*8-1 downto  81*8), w83 => Pw(121)( 83*8-1 downto  82*8), w84 => Pw(121)( 84*8-1 downto  83*8), 
w85 => Pw(121)( 85*8-1 downto  84*8), w86 => Pw(121)( 86*8-1 downto  85*8), w87 => Pw(121)( 87*8-1 downto  86*8), w88 => Pw(121)( 88*8-1 downto  87*8), 
w89 => Pw(121)( 89*8-1 downto  88*8), w90 => Pw(121)( 90*8-1 downto  89*8), w91 => Pw(121)( 91*8-1 downto  90*8), w92 => Pw(121)( 92*8-1 downto  91*8), 
w93 => Pw(121)( 93*8-1 downto  92*8), w94 => Pw(121)( 94*8-1 downto  93*8), w95 => Pw(121)( 95*8-1 downto  94*8), w96 => Pw(121)( 96*8-1 downto  95*8), 
w97 => Pw(121)( 97*8-1 downto  96*8), w98 => Pw(121)( 98*8-1 downto  97*8), w99 => Pw(121)( 99*8-1 downto  98*8), w100=> Pw(121)(100*8-1 downto  99*8), 
w101=> Pw(121)(101*8-1 downto 100*8), w102=> Pw(121)(102*8-1 downto 101*8), w103=> Pw(121)(103*8-1 downto 102*8), w104=> Pw(121)(104*8-1 downto 103*8), 
w105=> Pw(121)(105*8-1 downto 104*8), w106=> Pw(121)(106*8-1 downto 105*8), w107=> Pw(121)(107*8-1 downto 106*8), w108=> Pw(121)(108*8-1 downto 107*8), 
w109=> Pw(121)(109*8-1 downto 108*8), w110=> Pw(121)(110*8-1 downto 109*8), w111=> Pw(121)(111*8-1 downto 110*8), w112=> Pw(121)(112*8-1 downto 111*8), 
w113=> Pw(121)(113*8-1 downto 112*8), w114=> Pw(121)(114*8-1 downto 113*8), w115=> Pw(121)(115*8-1 downto 114*8), w116=> Pw(121)(116*8-1 downto 115*8), 
w117=> Pw(121)(117*8-1 downto 116*8), w118=> Pw(121)(118*8-1 downto 117*8), w119=> Pw(121)(119*8-1 downto 118*8), w120=> Pw(121)(120*8-1 downto 119*8), 
w121=> Pw(121)(121*8-1 downto 120*8), w122=> Pw(121)(122*8-1 downto 121*8), w123=> Pw(121)(123*8-1 downto 122*8), w124=> Pw(121)(124*8-1 downto 123*8), 
w125=> Pw(121)(125*8-1 downto 124*8), w126=> Pw(121)(126*8-1 downto 125*8), w127=> Pw(121)(127*8-1 downto 126*8), w128=> Pw(121)(128*8-1 downto 127*8), 
           d_out   => pca_d121_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_122_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(122)(     7 downto    0),   w02 => Pw(122)( 2*8-1 downto    8),   w03 => Pw(122)( 3*8-1 downto  2*8),   w04 => Pw(122)( 4*8-1 downto  3*8),   
w05 => Pw(122)( 5*8-1 downto  4*8),   w06 => Pw(122)( 6*8-1 downto  5*8),   w07 => Pw(122)( 7*8-1 downto  6*8),   w08 => Pw(122)( 8*8-1 downto  7*8),  
w09 => Pw(122)( 9*8-1 downto  8*8),   w10 => Pw(122)(10*8-1 downto  9*8),   w11 => Pw(122)(11*8-1 downto 10*8),   w12 => Pw(122)(12*8-1 downto 11*8),   
w13 => Pw(122)(13*8-1 downto 12*8),   w14 => Pw(122)(14*8-1 downto 13*8),   w15 => Pw(122)(15*8-1 downto 14*8),   w16 => Pw(122)(16*8-1 downto 15*8),  
w17 => Pw(122)(17*8-1 downto 16*8),   w18 => Pw(122)(18*8-1 downto 17*8),   w19 => Pw(122)(19*8-1 downto 18*8),   w20 => Pw(122)(20*8-1 downto 19*8),   
w21 => Pw(122)(21*8-1 downto 20*8),   w22 => Pw(122)(22*8-1 downto 21*8),   w23 => Pw(122)(23*8-1 downto 22*8),   w24 => Pw(122)(24*8-1 downto 23*8),  
w25 => Pw(122)(25*8-1 downto 24*8),   w26 => Pw(122)(26*8-1 downto 25*8),   w27 => Pw(122)(27*8-1 downto 26*8),   w28 => Pw(122)(28*8-1 downto 27*8),   
w29 => Pw(122)(29*8-1 downto 28*8),   w30 => Pw(122)(30*8-1 downto 29*8),   w31 => Pw(122)(31*8-1 downto 30*8),   w32 => Pw(122)(32*8-1 downto 31*8),  
w33 => Pw(122)(33*8-1 downto 32*8),   w34 => Pw(122)(34*8-1 downto 33*8),   w35 => Pw(122)(35*8-1 downto 34*8),   w36 => Pw(122)(36*8-1 downto 35*8),   
w37 => Pw(122)(37*8-1 downto 36*8),   w38 => Pw(122)(38*8-1 downto 37*8),   w39 => Pw(122)(39*8-1 downto 38*8),   w40 => Pw(122)(40*8-1 downto 39*8),  
w41 => Pw(122)(41*8-1 downto 40*8),   w42 => Pw(122)(42*8-1 downto 41*8),   w43 => Pw(122)(43*8-1 downto 42*8),   w44 => Pw(122)(44*8-1 downto 43*8),   
w45 => Pw(122)(45*8-1 downto 44*8),   w46 => Pw(122)(46*8-1 downto 45*8),   w47 => Pw(122)(47*8-1 downto 46*8),   w48 => Pw(122)(48*8-1 downto 47*8),  
w49 => Pw(122)(49*8-1 downto 48*8),   w50 => Pw(122)(50*8-1 downto 49*8),   w51 => Pw(122)(51*8-1 downto 50*8),   w52 => Pw(122)(52*8-1 downto 51*8),   
w53 => Pw(122)(53*8-1 downto 52*8),   w54 => Pw(122)(54*8-1 downto 53*8),   w55 => Pw(122)(55*8-1 downto 54*8),   w56 => Pw(122)(56*8-1 downto 55*8),  
w57 => Pw(122)(57*8-1 downto 56*8),   w58 => Pw(122)(58*8-1 downto 57*8),   w59 => Pw(122)(59*8-1 downto 58*8),   w60 => Pw(122)(60*8-1 downto 59*8),   
w61 => Pw(122)(61*8-1 downto 60*8),   w62 => Pw(122)(62*8-1 downto 61*8),   w63 => Pw(122)(63*8-1 downto 62*8),   w64 => Pw(122)(64*8-1 downto 63*8), 
w65 => Pw(122)( 65*8-1 downto  64*8), w66 => Pw(122)( 66*8-1 downto  65*8), w67 => Pw(122)( 67*8-1 downto  66*8), w68 => Pw(122)( 68*8-1 downto  67*8), 
w69 => Pw(122)( 69*8-1 downto  68*8), w70 => Pw(122)( 70*8-1 downto  69*8), w71 => Pw(122)( 71*8-1 downto  70*8), w72 => Pw(122)( 72*8-1 downto  71*8), 
w73 => Pw(122)( 73*8-1 downto  72*8), w74 => Pw(122)( 74*8-1 downto  73*8), w75 => Pw(122)( 75*8-1 downto  74*8), w76 => Pw(122)( 76*8-1 downto  75*8), 
w77 => Pw(122)( 77*8-1 downto  76*8), w78 => Pw(122)( 78*8-1 downto  77*8), w79 => Pw(122)( 79*8-1 downto  78*8), w80 => Pw(122)( 80*8-1 downto  79*8), 
w81 => Pw(122)( 81*8-1 downto  80*8), w82 => Pw(122)( 82*8-1 downto  81*8), w83 => Pw(122)( 83*8-1 downto  82*8), w84 => Pw(122)( 84*8-1 downto  83*8), 
w85 => Pw(122)( 85*8-1 downto  84*8), w86 => Pw(122)( 86*8-1 downto  85*8), w87 => Pw(122)( 87*8-1 downto  86*8), w88 => Pw(122)( 88*8-1 downto  87*8), 
w89 => Pw(122)( 89*8-1 downto  88*8), w90 => Pw(122)( 90*8-1 downto  89*8), w91 => Pw(122)( 91*8-1 downto  90*8), w92 => Pw(122)( 92*8-1 downto  91*8), 
w93 => Pw(122)( 93*8-1 downto  92*8), w94 => Pw(122)( 94*8-1 downto  93*8), w95 => Pw(122)( 95*8-1 downto  94*8), w96 => Pw(122)( 96*8-1 downto  95*8), 
w97 => Pw(122)( 97*8-1 downto  96*8), w98 => Pw(122)( 98*8-1 downto  97*8), w99 => Pw(122)( 99*8-1 downto  98*8), w100=> Pw(122)(100*8-1 downto  99*8), 
w101=> Pw(122)(101*8-1 downto 100*8), w102=> Pw(122)(102*8-1 downto 101*8), w103=> Pw(122)(103*8-1 downto 102*8), w104=> Pw(122)(104*8-1 downto 103*8), 
w105=> Pw(122)(105*8-1 downto 104*8), w106=> Pw(122)(106*8-1 downto 105*8), w107=> Pw(122)(107*8-1 downto 106*8), w108=> Pw(122)(108*8-1 downto 107*8), 
w109=> Pw(122)(109*8-1 downto 108*8), w110=> Pw(122)(110*8-1 downto 109*8), w111=> Pw(122)(111*8-1 downto 110*8), w112=> Pw(122)(112*8-1 downto 111*8), 
w113=> Pw(122)(113*8-1 downto 112*8), w114=> Pw(122)(114*8-1 downto 113*8), w115=> Pw(122)(115*8-1 downto 114*8), w116=> Pw(122)(116*8-1 downto 115*8), 
w117=> Pw(122)(117*8-1 downto 116*8), w118=> Pw(122)(118*8-1 downto 117*8), w119=> Pw(122)(119*8-1 downto 118*8), w120=> Pw(122)(120*8-1 downto 119*8), 
w121=> Pw(122)(121*8-1 downto 120*8), w122=> Pw(122)(122*8-1 downto 121*8), w123=> Pw(122)(123*8-1 downto 122*8), w124=> Pw(122)(124*8-1 downto 123*8), 
w125=> Pw(122)(125*8-1 downto 124*8), w126=> Pw(122)(126*8-1 downto 125*8), w127=> Pw(122)(127*8-1 downto 126*8), w128=> Pw(122)(128*8-1 downto 127*8), 
           d_out   => pca_d122_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_123_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(123)(     7 downto    0),   w02 => Pw(123)( 2*8-1 downto    8),   w03 => Pw(123)( 3*8-1 downto  2*8),   w04 => Pw(123)( 4*8-1 downto  3*8),   
w05 => Pw(123)( 5*8-1 downto  4*8),   w06 => Pw(123)( 6*8-1 downto  5*8),   w07 => Pw(123)( 7*8-1 downto  6*8),   w08 => Pw(123)( 8*8-1 downto  7*8),  
w09 => Pw(123)( 9*8-1 downto  8*8),   w10 => Pw(123)(10*8-1 downto  9*8),   w11 => Pw(123)(11*8-1 downto 10*8),   w12 => Pw(123)(12*8-1 downto 11*8),   
w13 => Pw(123)(13*8-1 downto 12*8),   w14 => Pw(123)(14*8-1 downto 13*8),   w15 => Pw(123)(15*8-1 downto 14*8),   w16 => Pw(123)(16*8-1 downto 15*8),  
w17 => Pw(123)(17*8-1 downto 16*8),   w18 => Pw(123)(18*8-1 downto 17*8),   w19 => Pw(123)(19*8-1 downto 18*8),   w20 => Pw(123)(20*8-1 downto 19*8),   
w21 => Pw(123)(21*8-1 downto 20*8),   w22 => Pw(123)(22*8-1 downto 21*8),   w23 => Pw(123)(23*8-1 downto 22*8),   w24 => Pw(123)(24*8-1 downto 23*8),  
w25 => Pw(123)(25*8-1 downto 24*8),   w26 => Pw(123)(26*8-1 downto 25*8),   w27 => Pw(123)(27*8-1 downto 26*8),   w28 => Pw(123)(28*8-1 downto 27*8),   
w29 => Pw(123)(29*8-1 downto 28*8),   w30 => Pw(123)(30*8-1 downto 29*8),   w31 => Pw(123)(31*8-1 downto 30*8),   w32 => Pw(123)(32*8-1 downto 31*8),  
w33 => Pw(123)(33*8-1 downto 32*8),   w34 => Pw(123)(34*8-1 downto 33*8),   w35 => Pw(123)(35*8-1 downto 34*8),   w36 => Pw(123)(36*8-1 downto 35*8),   
w37 => Pw(123)(37*8-1 downto 36*8),   w38 => Pw(123)(38*8-1 downto 37*8),   w39 => Pw(123)(39*8-1 downto 38*8),   w40 => Pw(123)(40*8-1 downto 39*8),  
w41 => Pw(123)(41*8-1 downto 40*8),   w42 => Pw(123)(42*8-1 downto 41*8),   w43 => Pw(123)(43*8-1 downto 42*8),   w44 => Pw(123)(44*8-1 downto 43*8),   
w45 => Pw(123)(45*8-1 downto 44*8),   w46 => Pw(123)(46*8-1 downto 45*8),   w47 => Pw(123)(47*8-1 downto 46*8),   w48 => Pw(123)(48*8-1 downto 47*8),  
w49 => Pw(123)(49*8-1 downto 48*8),   w50 => Pw(123)(50*8-1 downto 49*8),   w51 => Pw(123)(51*8-1 downto 50*8),   w52 => Pw(123)(52*8-1 downto 51*8),   
w53 => Pw(123)(53*8-1 downto 52*8),   w54 => Pw(123)(54*8-1 downto 53*8),   w55 => Pw(123)(55*8-1 downto 54*8),   w56 => Pw(123)(56*8-1 downto 55*8),  
w57 => Pw(123)(57*8-1 downto 56*8),   w58 => Pw(123)(58*8-1 downto 57*8),   w59 => Pw(123)(59*8-1 downto 58*8),   w60 => Pw(123)(60*8-1 downto 59*8),   
w61 => Pw(123)(61*8-1 downto 60*8),   w62 => Pw(123)(62*8-1 downto 61*8),   w63 => Pw(123)(63*8-1 downto 62*8),   w64 => Pw(123)(64*8-1 downto 63*8), 
w65 => Pw(123)( 65*8-1 downto  64*8), w66 => Pw(123)( 66*8-1 downto  65*8), w67 => Pw(123)( 67*8-1 downto  66*8), w68 => Pw(123)( 68*8-1 downto  67*8), 
w69 => Pw(123)( 69*8-1 downto  68*8), w70 => Pw(123)( 70*8-1 downto  69*8), w71 => Pw(123)( 71*8-1 downto  70*8), w72 => Pw(123)( 72*8-1 downto  71*8), 
w73 => Pw(123)( 73*8-1 downto  72*8), w74 => Pw(123)( 74*8-1 downto  73*8), w75 => Pw(123)( 75*8-1 downto  74*8), w76 => Pw(123)( 76*8-1 downto  75*8), 
w77 => Pw(123)( 77*8-1 downto  76*8), w78 => Pw(123)( 78*8-1 downto  77*8), w79 => Pw(123)( 79*8-1 downto  78*8), w80 => Pw(123)( 80*8-1 downto  79*8), 
w81 => Pw(123)( 81*8-1 downto  80*8), w82 => Pw(123)( 82*8-1 downto  81*8), w83 => Pw(123)( 83*8-1 downto  82*8), w84 => Pw(123)( 84*8-1 downto  83*8), 
w85 => Pw(123)( 85*8-1 downto  84*8), w86 => Pw(123)( 86*8-1 downto  85*8), w87 => Pw(123)( 87*8-1 downto  86*8), w88 => Pw(123)( 88*8-1 downto  87*8), 
w89 => Pw(123)( 89*8-1 downto  88*8), w90 => Pw(123)( 90*8-1 downto  89*8), w91 => Pw(123)( 91*8-1 downto  90*8), w92 => Pw(123)( 92*8-1 downto  91*8), 
w93 => Pw(123)( 93*8-1 downto  92*8), w94 => Pw(123)( 94*8-1 downto  93*8), w95 => Pw(123)( 95*8-1 downto  94*8), w96 => Pw(123)( 96*8-1 downto  95*8), 
w97 => Pw(123)( 97*8-1 downto  96*8), w98 => Pw(123)( 98*8-1 downto  97*8), w99 => Pw(123)( 99*8-1 downto  98*8), w100=> Pw(123)(100*8-1 downto  99*8), 
w101=> Pw(123)(101*8-1 downto 100*8), w102=> Pw(123)(102*8-1 downto 101*8), w103=> Pw(123)(103*8-1 downto 102*8), w104=> Pw(123)(104*8-1 downto 103*8), 
w105=> Pw(123)(105*8-1 downto 104*8), w106=> Pw(123)(106*8-1 downto 105*8), w107=> Pw(123)(107*8-1 downto 106*8), w108=> Pw(123)(108*8-1 downto 107*8), 
w109=> Pw(123)(109*8-1 downto 108*8), w110=> Pw(123)(110*8-1 downto 109*8), w111=> Pw(123)(111*8-1 downto 110*8), w112=> Pw(123)(112*8-1 downto 111*8), 
w113=> Pw(123)(113*8-1 downto 112*8), w114=> Pw(123)(114*8-1 downto 113*8), w115=> Pw(123)(115*8-1 downto 114*8), w116=> Pw(123)(116*8-1 downto 115*8), 
w117=> Pw(123)(117*8-1 downto 116*8), w118=> Pw(123)(118*8-1 downto 117*8), w119=> Pw(123)(119*8-1 downto 118*8), w120=> Pw(123)(120*8-1 downto 119*8), 
w121=> Pw(123)(121*8-1 downto 120*8), w122=> Pw(123)(122*8-1 downto 121*8), w123=> Pw(123)(123*8-1 downto 122*8), w124=> Pw(123)(124*8-1 downto 123*8), 
w125=> Pw(123)(125*8-1 downto 124*8), w126=> Pw(123)(126*8-1 downto 125*8), w127=> Pw(123)(127*8-1 downto 126*8), w128=> Pw(123)(128*8-1 downto 127*8), 
           d_out   => pca_d123_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_124_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(124)(     7 downto    0),   w02 => Pw(124)( 2*8-1 downto    8),   w03 => Pw(124)( 3*8-1 downto  2*8),   w04 => Pw(124)( 4*8-1 downto  3*8),   
w05 => Pw(124)( 5*8-1 downto  4*8),   w06 => Pw(124)( 6*8-1 downto  5*8),   w07 => Pw(124)( 7*8-1 downto  6*8),   w08 => Pw(124)( 8*8-1 downto  7*8),  
w09 => Pw(124)( 9*8-1 downto  8*8),   w10 => Pw(124)(10*8-1 downto  9*8),   w11 => Pw(124)(11*8-1 downto 10*8),   w12 => Pw(124)(12*8-1 downto 11*8),   
w13 => Pw(124)(13*8-1 downto 12*8),   w14 => Pw(124)(14*8-1 downto 13*8),   w15 => Pw(124)(15*8-1 downto 14*8),   w16 => Pw(124)(16*8-1 downto 15*8),  
w17 => Pw(124)(17*8-1 downto 16*8),   w18 => Pw(124)(18*8-1 downto 17*8),   w19 => Pw(124)(19*8-1 downto 18*8),   w20 => Pw(124)(20*8-1 downto 19*8),   
w21 => Pw(124)(21*8-1 downto 20*8),   w22 => Pw(124)(22*8-1 downto 21*8),   w23 => Pw(124)(23*8-1 downto 22*8),   w24 => Pw(124)(24*8-1 downto 23*8),  
w25 => Pw(124)(25*8-1 downto 24*8),   w26 => Pw(124)(26*8-1 downto 25*8),   w27 => Pw(124)(27*8-1 downto 26*8),   w28 => Pw(124)(28*8-1 downto 27*8),   
w29 => Pw(124)(29*8-1 downto 28*8),   w30 => Pw(124)(30*8-1 downto 29*8),   w31 => Pw(124)(31*8-1 downto 30*8),   w32 => Pw(124)(32*8-1 downto 31*8),  
w33 => Pw(124)(33*8-1 downto 32*8),   w34 => Pw(124)(34*8-1 downto 33*8),   w35 => Pw(124)(35*8-1 downto 34*8),   w36 => Pw(124)(36*8-1 downto 35*8),   
w37 => Pw(124)(37*8-1 downto 36*8),   w38 => Pw(124)(38*8-1 downto 37*8),   w39 => Pw(124)(39*8-1 downto 38*8),   w40 => Pw(124)(40*8-1 downto 39*8),  
w41 => Pw(124)(41*8-1 downto 40*8),   w42 => Pw(124)(42*8-1 downto 41*8),   w43 => Pw(124)(43*8-1 downto 42*8),   w44 => Pw(124)(44*8-1 downto 43*8),   
w45 => Pw(124)(45*8-1 downto 44*8),   w46 => Pw(124)(46*8-1 downto 45*8),   w47 => Pw(124)(47*8-1 downto 46*8),   w48 => Pw(124)(48*8-1 downto 47*8),  
w49 => Pw(124)(49*8-1 downto 48*8),   w50 => Pw(124)(50*8-1 downto 49*8),   w51 => Pw(124)(51*8-1 downto 50*8),   w52 => Pw(124)(52*8-1 downto 51*8),   
w53 => Pw(124)(53*8-1 downto 52*8),   w54 => Pw(124)(54*8-1 downto 53*8),   w55 => Pw(124)(55*8-1 downto 54*8),   w56 => Pw(124)(56*8-1 downto 55*8),  
w57 => Pw(124)(57*8-1 downto 56*8),   w58 => Pw(124)(58*8-1 downto 57*8),   w59 => Pw(124)(59*8-1 downto 58*8),   w60 => Pw(124)(60*8-1 downto 59*8),   
w61 => Pw(124)(61*8-1 downto 60*8),   w62 => Pw(124)(62*8-1 downto 61*8),   w63 => Pw(124)(63*8-1 downto 62*8),   w64 => Pw(124)(64*8-1 downto 63*8), 
w65 => Pw(124)( 65*8-1 downto  64*8), w66 => Pw(124)( 66*8-1 downto  65*8), w67 => Pw(124)( 67*8-1 downto  66*8), w68 => Pw(124)( 68*8-1 downto  67*8), 
w69 => Pw(124)( 69*8-1 downto  68*8), w70 => Pw(124)( 70*8-1 downto  69*8), w71 => Pw(124)( 71*8-1 downto  70*8), w72 => Pw(124)( 72*8-1 downto  71*8), 
w73 => Pw(124)( 73*8-1 downto  72*8), w74 => Pw(124)( 74*8-1 downto  73*8), w75 => Pw(124)( 75*8-1 downto  74*8), w76 => Pw(124)( 76*8-1 downto  75*8), 
w77 => Pw(124)( 77*8-1 downto  76*8), w78 => Pw(124)( 78*8-1 downto  77*8), w79 => Pw(124)( 79*8-1 downto  78*8), w80 => Pw(124)( 80*8-1 downto  79*8), 
w81 => Pw(124)( 81*8-1 downto  80*8), w82 => Pw(124)( 82*8-1 downto  81*8), w83 => Pw(124)( 83*8-1 downto  82*8), w84 => Pw(124)( 84*8-1 downto  83*8), 
w85 => Pw(124)( 85*8-1 downto  84*8), w86 => Pw(124)( 86*8-1 downto  85*8), w87 => Pw(124)( 87*8-1 downto  86*8), w88 => Pw(124)( 88*8-1 downto  87*8), 
w89 => Pw(124)( 89*8-1 downto  88*8), w90 => Pw(124)( 90*8-1 downto  89*8), w91 => Pw(124)( 91*8-1 downto  90*8), w92 => Pw(124)( 92*8-1 downto  91*8), 
w93 => Pw(124)( 93*8-1 downto  92*8), w94 => Pw(124)( 94*8-1 downto  93*8), w95 => Pw(124)( 95*8-1 downto  94*8), w96 => Pw(124)( 96*8-1 downto  95*8), 
w97 => Pw(124)( 97*8-1 downto  96*8), w98 => Pw(124)( 98*8-1 downto  97*8), w99 => Pw(124)( 99*8-1 downto  98*8), w100=> Pw(124)(100*8-1 downto  99*8), 
w101=> Pw(124)(101*8-1 downto 100*8), w102=> Pw(124)(102*8-1 downto 101*8), w103=> Pw(124)(103*8-1 downto 102*8), w104=> Pw(124)(104*8-1 downto 103*8), 
w105=> Pw(124)(105*8-1 downto 104*8), w106=> Pw(124)(106*8-1 downto 105*8), w107=> Pw(124)(107*8-1 downto 106*8), w108=> Pw(124)(108*8-1 downto 107*8), 
w109=> Pw(124)(109*8-1 downto 108*8), w110=> Pw(124)(110*8-1 downto 109*8), w111=> Pw(124)(111*8-1 downto 110*8), w112=> Pw(124)(112*8-1 downto 111*8), 
w113=> Pw(124)(113*8-1 downto 112*8), w114=> Pw(124)(114*8-1 downto 113*8), w115=> Pw(124)(115*8-1 downto 114*8), w116=> Pw(124)(116*8-1 downto 115*8), 
w117=> Pw(124)(117*8-1 downto 116*8), w118=> Pw(124)(118*8-1 downto 117*8), w119=> Pw(124)(119*8-1 downto 118*8), w120=> Pw(124)(120*8-1 downto 119*8), 
w121=> Pw(124)(121*8-1 downto 120*8), w122=> Pw(124)(122*8-1 downto 121*8), w123=> Pw(124)(123*8-1 downto 122*8), w124=> Pw(124)(124*8-1 downto 123*8), 
w125=> Pw(124)(125*8-1 downto 124*8), w126=> Pw(124)(126*8-1 downto 125*8), w127=> Pw(124)(127*8-1 downto 126*8), w128=> Pw(124)(128*8-1 downto 127*8), 
           d_out   => pca_d124_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_125_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(125)(     7 downto    0),   w02 => Pw(125)( 2*8-1 downto    8),   w03 => Pw(125)( 3*8-1 downto  2*8),   w04 => Pw(125)( 4*8-1 downto  3*8),   
w05 => Pw(125)( 5*8-1 downto  4*8),   w06 => Pw(125)( 6*8-1 downto  5*8),   w07 => Pw(125)( 7*8-1 downto  6*8),   w08 => Pw(125)( 8*8-1 downto  7*8),  
w09 => Pw(125)( 9*8-1 downto  8*8),   w10 => Pw(125)(10*8-1 downto  9*8),   w11 => Pw(125)(11*8-1 downto 10*8),   w12 => Pw(125)(12*8-1 downto 11*8),   
w13 => Pw(125)(13*8-1 downto 12*8),   w14 => Pw(125)(14*8-1 downto 13*8),   w15 => Pw(125)(15*8-1 downto 14*8),   w16 => Pw(125)(16*8-1 downto 15*8),  
w17 => Pw(125)(17*8-1 downto 16*8),   w18 => Pw(125)(18*8-1 downto 17*8),   w19 => Pw(125)(19*8-1 downto 18*8),   w20 => Pw(125)(20*8-1 downto 19*8),   
w21 => Pw(125)(21*8-1 downto 20*8),   w22 => Pw(125)(22*8-1 downto 21*8),   w23 => Pw(125)(23*8-1 downto 22*8),   w24 => Pw(125)(24*8-1 downto 23*8),  
w25 => Pw(125)(25*8-1 downto 24*8),   w26 => Pw(125)(26*8-1 downto 25*8),   w27 => Pw(125)(27*8-1 downto 26*8),   w28 => Pw(125)(28*8-1 downto 27*8),   
w29 => Pw(125)(29*8-1 downto 28*8),   w30 => Pw(125)(30*8-1 downto 29*8),   w31 => Pw(125)(31*8-1 downto 30*8),   w32 => Pw(125)(32*8-1 downto 31*8),  
w33 => Pw(125)(33*8-1 downto 32*8),   w34 => Pw(125)(34*8-1 downto 33*8),   w35 => Pw(125)(35*8-1 downto 34*8),   w36 => Pw(125)(36*8-1 downto 35*8),   
w37 => Pw(125)(37*8-1 downto 36*8),   w38 => Pw(125)(38*8-1 downto 37*8),   w39 => Pw(125)(39*8-1 downto 38*8),   w40 => Pw(125)(40*8-1 downto 39*8),  
w41 => Pw(125)(41*8-1 downto 40*8),   w42 => Pw(125)(42*8-1 downto 41*8),   w43 => Pw(125)(43*8-1 downto 42*8),   w44 => Pw(125)(44*8-1 downto 43*8),   
w45 => Pw(125)(45*8-1 downto 44*8),   w46 => Pw(125)(46*8-1 downto 45*8),   w47 => Pw(125)(47*8-1 downto 46*8),   w48 => Pw(125)(48*8-1 downto 47*8),  
w49 => Pw(125)(49*8-1 downto 48*8),   w50 => Pw(125)(50*8-1 downto 49*8),   w51 => Pw(125)(51*8-1 downto 50*8),   w52 => Pw(125)(52*8-1 downto 51*8),   
w53 => Pw(125)(53*8-1 downto 52*8),   w54 => Pw(125)(54*8-1 downto 53*8),   w55 => Pw(125)(55*8-1 downto 54*8),   w56 => Pw(125)(56*8-1 downto 55*8),  
w57 => Pw(125)(57*8-1 downto 56*8),   w58 => Pw(125)(58*8-1 downto 57*8),   w59 => Pw(125)(59*8-1 downto 58*8),   w60 => Pw(125)(60*8-1 downto 59*8),   
w61 => Pw(125)(61*8-1 downto 60*8),   w62 => Pw(125)(62*8-1 downto 61*8),   w63 => Pw(125)(63*8-1 downto 62*8),   w64 => Pw(125)(64*8-1 downto 63*8), 
w65 => Pw(125)( 65*8-1 downto  64*8), w66 => Pw(125)( 66*8-1 downto  65*8), w67 => Pw(125)( 67*8-1 downto  66*8), w68 => Pw(125)( 68*8-1 downto  67*8), 
w69 => Pw(125)( 69*8-1 downto  68*8), w70 => Pw(125)( 70*8-1 downto  69*8), w71 => Pw(125)( 71*8-1 downto  70*8), w72 => Pw(125)( 72*8-1 downto  71*8), 
w73 => Pw(125)( 73*8-1 downto  72*8), w74 => Pw(125)( 74*8-1 downto  73*8), w75 => Pw(125)( 75*8-1 downto  74*8), w76 => Pw(125)( 76*8-1 downto  75*8), 
w77 => Pw(125)( 77*8-1 downto  76*8), w78 => Pw(125)( 78*8-1 downto  77*8), w79 => Pw(125)( 79*8-1 downto  78*8), w80 => Pw(125)( 80*8-1 downto  79*8), 
w81 => Pw(125)( 81*8-1 downto  80*8), w82 => Pw(125)( 82*8-1 downto  81*8), w83 => Pw(125)( 83*8-1 downto  82*8), w84 => Pw(125)( 84*8-1 downto  83*8), 
w85 => Pw(125)( 85*8-1 downto  84*8), w86 => Pw(125)( 86*8-1 downto  85*8), w87 => Pw(125)( 87*8-1 downto  86*8), w88 => Pw(125)( 88*8-1 downto  87*8), 
w89 => Pw(125)( 89*8-1 downto  88*8), w90 => Pw(125)( 90*8-1 downto  89*8), w91 => Pw(125)( 91*8-1 downto  90*8), w92 => Pw(125)( 92*8-1 downto  91*8), 
w93 => Pw(125)( 93*8-1 downto  92*8), w94 => Pw(125)( 94*8-1 downto  93*8), w95 => Pw(125)( 95*8-1 downto  94*8), w96 => Pw(125)( 96*8-1 downto  95*8), 
w97 => Pw(125)( 97*8-1 downto  96*8), w98 => Pw(125)( 98*8-1 downto  97*8), w99 => Pw(125)( 99*8-1 downto  98*8), w100=> Pw(125)(100*8-1 downto  99*8), 
w101=> Pw(125)(101*8-1 downto 100*8), w102=> Pw(125)(102*8-1 downto 101*8), w103=> Pw(125)(103*8-1 downto 102*8), w104=> Pw(125)(104*8-1 downto 103*8), 
w105=> Pw(125)(105*8-1 downto 104*8), w106=> Pw(125)(106*8-1 downto 105*8), w107=> Pw(125)(107*8-1 downto 106*8), w108=> Pw(125)(108*8-1 downto 107*8), 
w109=> Pw(125)(109*8-1 downto 108*8), w110=> Pw(125)(110*8-1 downto 109*8), w111=> Pw(125)(111*8-1 downto 110*8), w112=> Pw(125)(112*8-1 downto 111*8), 
w113=> Pw(125)(113*8-1 downto 112*8), w114=> Pw(125)(114*8-1 downto 113*8), w115=> Pw(125)(115*8-1 downto 114*8), w116=> Pw(125)(116*8-1 downto 115*8), 
w117=> Pw(125)(117*8-1 downto 116*8), w118=> Pw(125)(118*8-1 downto 117*8), w119=> Pw(125)(119*8-1 downto 118*8), w120=> Pw(125)(120*8-1 downto 119*8), 
w121=> Pw(125)(121*8-1 downto 120*8), w122=> Pw(125)(122*8-1 downto 121*8), w123=> Pw(125)(123*8-1 downto 122*8), w124=> Pw(125)(124*8-1 downto 123*8), 
w125=> Pw(125)(125*8-1 downto 124*8), w126=> Pw(125)(126*8-1 downto 125*8), w127=> Pw(125)(127*8-1 downto 126*8), w128=> Pw(125)(128*8-1 downto 127*8), 
           d_out   => pca_d125_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_126_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(126)(     7 downto    0),   w02 => Pw(126)( 2*8-1 downto    8),   w03 => Pw(126)( 3*8-1 downto  2*8),   w04 => Pw(126)( 4*8-1 downto  3*8),   
w05 => Pw(126)( 5*8-1 downto  4*8),   w06 => Pw(126)( 6*8-1 downto  5*8),   w07 => Pw(126)( 7*8-1 downto  6*8),   w08 => Pw(126)( 8*8-1 downto  7*8),  
w09 => Pw(126)( 9*8-1 downto  8*8),   w10 => Pw(126)(10*8-1 downto  9*8),   w11 => Pw(126)(11*8-1 downto 10*8),   w12 => Pw(126)(12*8-1 downto 11*8),   
w13 => Pw(126)(13*8-1 downto 12*8),   w14 => Pw(126)(14*8-1 downto 13*8),   w15 => Pw(126)(15*8-1 downto 14*8),   w16 => Pw(126)(16*8-1 downto 15*8),  
w17 => Pw(126)(17*8-1 downto 16*8),   w18 => Pw(126)(18*8-1 downto 17*8),   w19 => Pw(126)(19*8-1 downto 18*8),   w20 => Pw(126)(20*8-1 downto 19*8),   
w21 => Pw(126)(21*8-1 downto 20*8),   w22 => Pw(126)(22*8-1 downto 21*8),   w23 => Pw(126)(23*8-1 downto 22*8),   w24 => Pw(126)(24*8-1 downto 23*8),  
w25 => Pw(126)(25*8-1 downto 24*8),   w26 => Pw(126)(26*8-1 downto 25*8),   w27 => Pw(126)(27*8-1 downto 26*8),   w28 => Pw(126)(28*8-1 downto 27*8),   
w29 => Pw(126)(29*8-1 downto 28*8),   w30 => Pw(126)(30*8-1 downto 29*8),   w31 => Pw(126)(31*8-1 downto 30*8),   w32 => Pw(126)(32*8-1 downto 31*8),  
w33 => Pw(126)(33*8-1 downto 32*8),   w34 => Pw(126)(34*8-1 downto 33*8),   w35 => Pw(126)(35*8-1 downto 34*8),   w36 => Pw(126)(36*8-1 downto 35*8),   
w37 => Pw(126)(37*8-1 downto 36*8),   w38 => Pw(126)(38*8-1 downto 37*8),   w39 => Pw(126)(39*8-1 downto 38*8),   w40 => Pw(126)(40*8-1 downto 39*8),  
w41 => Pw(126)(41*8-1 downto 40*8),   w42 => Pw(126)(42*8-1 downto 41*8),   w43 => Pw(126)(43*8-1 downto 42*8),   w44 => Pw(126)(44*8-1 downto 43*8),   
w45 => Pw(126)(45*8-1 downto 44*8),   w46 => Pw(126)(46*8-1 downto 45*8),   w47 => Pw(126)(47*8-1 downto 46*8),   w48 => Pw(126)(48*8-1 downto 47*8),  
w49 => Pw(126)(49*8-1 downto 48*8),   w50 => Pw(126)(50*8-1 downto 49*8),   w51 => Pw(126)(51*8-1 downto 50*8),   w52 => Pw(126)(52*8-1 downto 51*8),   
w53 => Pw(126)(53*8-1 downto 52*8),   w54 => Pw(126)(54*8-1 downto 53*8),   w55 => Pw(126)(55*8-1 downto 54*8),   w56 => Pw(126)(56*8-1 downto 55*8),  
w57 => Pw(126)(57*8-1 downto 56*8),   w58 => Pw(126)(58*8-1 downto 57*8),   w59 => Pw(126)(59*8-1 downto 58*8),   w60 => Pw(126)(60*8-1 downto 59*8),   
w61 => Pw(126)(61*8-1 downto 60*8),   w62 => Pw(126)(62*8-1 downto 61*8),   w63 => Pw(126)(63*8-1 downto 62*8),   w64 => Pw(126)(64*8-1 downto 63*8), 
w65 => Pw(126)( 65*8-1 downto  64*8), w66 => Pw(126)( 66*8-1 downto  65*8), w67 => Pw(126)( 67*8-1 downto  66*8), w68 => Pw(126)( 68*8-1 downto  67*8), 
w69 => Pw(126)( 69*8-1 downto  68*8), w70 => Pw(126)( 70*8-1 downto  69*8), w71 => Pw(126)( 71*8-1 downto  70*8), w72 => Pw(126)( 72*8-1 downto  71*8), 
w73 => Pw(126)( 73*8-1 downto  72*8), w74 => Pw(126)( 74*8-1 downto  73*8), w75 => Pw(126)( 75*8-1 downto  74*8), w76 => Pw(126)( 76*8-1 downto  75*8), 
w77 => Pw(126)( 77*8-1 downto  76*8), w78 => Pw(126)( 78*8-1 downto  77*8), w79 => Pw(126)( 79*8-1 downto  78*8), w80 => Pw(126)( 80*8-1 downto  79*8), 
w81 => Pw(126)( 81*8-1 downto  80*8), w82 => Pw(126)( 82*8-1 downto  81*8), w83 => Pw(126)( 83*8-1 downto  82*8), w84 => Pw(126)( 84*8-1 downto  83*8), 
w85 => Pw(126)( 85*8-1 downto  84*8), w86 => Pw(126)( 86*8-1 downto  85*8), w87 => Pw(126)( 87*8-1 downto  86*8), w88 => Pw(126)( 88*8-1 downto  87*8), 
w89 => Pw(126)( 89*8-1 downto  88*8), w90 => Pw(126)( 90*8-1 downto  89*8), w91 => Pw(126)( 91*8-1 downto  90*8), w92 => Pw(126)( 92*8-1 downto  91*8), 
w93 => Pw(126)( 93*8-1 downto  92*8), w94 => Pw(126)( 94*8-1 downto  93*8), w95 => Pw(126)( 95*8-1 downto  94*8), w96 => Pw(126)( 96*8-1 downto  95*8), 
w97 => Pw(126)( 97*8-1 downto  96*8), w98 => Pw(126)( 98*8-1 downto  97*8), w99 => Pw(126)( 99*8-1 downto  98*8), w100=> Pw(126)(100*8-1 downto  99*8), 
w101=> Pw(126)(101*8-1 downto 100*8), w102=> Pw(126)(102*8-1 downto 101*8), w103=> Pw(126)(103*8-1 downto 102*8), w104=> Pw(126)(104*8-1 downto 103*8), 
w105=> Pw(126)(105*8-1 downto 104*8), w106=> Pw(126)(106*8-1 downto 105*8), w107=> Pw(126)(107*8-1 downto 106*8), w108=> Pw(126)(108*8-1 downto 107*8), 
w109=> Pw(126)(109*8-1 downto 108*8), w110=> Pw(126)(110*8-1 downto 109*8), w111=> Pw(126)(111*8-1 downto 110*8), w112=> Pw(126)(112*8-1 downto 111*8), 
w113=> Pw(126)(113*8-1 downto 112*8), w114=> Pw(126)(114*8-1 downto 113*8), w115=> Pw(126)(115*8-1 downto 114*8), w116=> Pw(126)(116*8-1 downto 115*8), 
w117=> Pw(126)(117*8-1 downto 116*8), w118=> Pw(126)(118*8-1 downto 117*8), w119=> Pw(126)(119*8-1 downto 118*8), w120=> Pw(126)(120*8-1 downto 119*8), 
w121=> Pw(126)(121*8-1 downto 120*8), w122=> Pw(126)(122*8-1 downto 121*8), w123=> Pw(126)(123*8-1 downto 122*8), w124=> Pw(126)(124*8-1 downto 123*8), 
w125=> Pw(126)(125*8-1 downto 124*8), w126=> Pw(126)(126*8-1 downto 125*8), w127=> Pw(126)(127*8-1 downto 126*8), w128=> Pw(126)(128*8-1 downto 127*8), 
           d_out   => pca_d126_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_127_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(127)(     7 downto    0),   w02 => Pw(127)( 2*8-1 downto    8),   w03 => Pw(127)( 3*8-1 downto  2*8),   w04 => Pw(127)( 4*8-1 downto  3*8),   
w05 => Pw(127)( 5*8-1 downto  4*8),   w06 => Pw(127)( 6*8-1 downto  5*8),   w07 => Pw(127)( 7*8-1 downto  6*8),   w08 => Pw(127)( 8*8-1 downto  7*8),  
w09 => Pw(127)( 9*8-1 downto  8*8),   w10 => Pw(127)(10*8-1 downto  9*8),   w11 => Pw(127)(11*8-1 downto 10*8),   w12 => Pw(127)(12*8-1 downto 11*8),   
w13 => Pw(127)(13*8-1 downto 12*8),   w14 => Pw(127)(14*8-1 downto 13*8),   w15 => Pw(127)(15*8-1 downto 14*8),   w16 => Pw(127)(16*8-1 downto 15*8),  
w17 => Pw(127)(17*8-1 downto 16*8),   w18 => Pw(127)(18*8-1 downto 17*8),   w19 => Pw(127)(19*8-1 downto 18*8),   w20 => Pw(127)(20*8-1 downto 19*8),   
w21 => Pw(127)(21*8-1 downto 20*8),   w22 => Pw(127)(22*8-1 downto 21*8),   w23 => Pw(127)(23*8-1 downto 22*8),   w24 => Pw(127)(24*8-1 downto 23*8),  
w25 => Pw(127)(25*8-1 downto 24*8),   w26 => Pw(127)(26*8-1 downto 25*8),   w27 => Pw(127)(27*8-1 downto 26*8),   w28 => Pw(127)(28*8-1 downto 27*8),   
w29 => Pw(127)(29*8-1 downto 28*8),   w30 => Pw(127)(30*8-1 downto 29*8),   w31 => Pw(127)(31*8-1 downto 30*8),   w32 => Pw(127)(32*8-1 downto 31*8),  
w33 => Pw(127)(33*8-1 downto 32*8),   w34 => Pw(127)(34*8-1 downto 33*8),   w35 => Pw(127)(35*8-1 downto 34*8),   w36 => Pw(127)(36*8-1 downto 35*8),   
w37 => Pw(127)(37*8-1 downto 36*8),   w38 => Pw(127)(38*8-1 downto 37*8),   w39 => Pw(127)(39*8-1 downto 38*8),   w40 => Pw(127)(40*8-1 downto 39*8),  
w41 => Pw(127)(41*8-1 downto 40*8),   w42 => Pw(127)(42*8-1 downto 41*8),   w43 => Pw(127)(43*8-1 downto 42*8),   w44 => Pw(127)(44*8-1 downto 43*8),   
w45 => Pw(127)(45*8-1 downto 44*8),   w46 => Pw(127)(46*8-1 downto 45*8),   w47 => Pw(127)(47*8-1 downto 46*8),   w48 => Pw(127)(48*8-1 downto 47*8),  
w49 => Pw(127)(49*8-1 downto 48*8),   w50 => Pw(127)(50*8-1 downto 49*8),   w51 => Pw(127)(51*8-1 downto 50*8),   w52 => Pw(127)(52*8-1 downto 51*8),   
w53 => Pw(127)(53*8-1 downto 52*8),   w54 => Pw(127)(54*8-1 downto 53*8),   w55 => Pw(127)(55*8-1 downto 54*8),   w56 => Pw(127)(56*8-1 downto 55*8),  
w57 => Pw(127)(57*8-1 downto 56*8),   w58 => Pw(127)(58*8-1 downto 57*8),   w59 => Pw(127)(59*8-1 downto 58*8),   w60 => Pw(127)(60*8-1 downto 59*8),   
w61 => Pw(127)(61*8-1 downto 60*8),   w62 => Pw(127)(62*8-1 downto 61*8),   w63 => Pw(127)(63*8-1 downto 62*8),   w64 => Pw(127)(64*8-1 downto 63*8), 
w65 => Pw(127)( 65*8-1 downto  64*8), w66 => Pw(127)( 66*8-1 downto  65*8), w67 => Pw(127)( 67*8-1 downto  66*8), w68 => Pw(127)( 68*8-1 downto  67*8), 
w69 => Pw(127)( 69*8-1 downto  68*8), w70 => Pw(127)( 70*8-1 downto  69*8), w71 => Pw(127)( 71*8-1 downto  70*8), w72 => Pw(127)( 72*8-1 downto  71*8), 
w73 => Pw(127)( 73*8-1 downto  72*8), w74 => Pw(127)( 74*8-1 downto  73*8), w75 => Pw(127)( 75*8-1 downto  74*8), w76 => Pw(127)( 76*8-1 downto  75*8), 
w77 => Pw(127)( 77*8-1 downto  76*8), w78 => Pw(127)( 78*8-1 downto  77*8), w79 => Pw(127)( 79*8-1 downto  78*8), w80 => Pw(127)( 80*8-1 downto  79*8), 
w81 => Pw(127)( 81*8-1 downto  80*8), w82 => Pw(127)( 82*8-1 downto  81*8), w83 => Pw(127)( 83*8-1 downto  82*8), w84 => Pw(127)( 84*8-1 downto  83*8), 
w85 => Pw(127)( 85*8-1 downto  84*8), w86 => Pw(127)( 86*8-1 downto  85*8), w87 => Pw(127)( 87*8-1 downto  86*8), w88 => Pw(127)( 88*8-1 downto  87*8), 
w89 => Pw(127)( 89*8-1 downto  88*8), w90 => Pw(127)( 90*8-1 downto  89*8), w91 => Pw(127)( 91*8-1 downto  90*8), w92 => Pw(127)( 92*8-1 downto  91*8), 
w93 => Pw(127)( 93*8-1 downto  92*8), w94 => Pw(127)( 94*8-1 downto  93*8), w95 => Pw(127)( 95*8-1 downto  94*8), w96 => Pw(127)( 96*8-1 downto  95*8), 
w97 => Pw(127)( 97*8-1 downto  96*8), w98 => Pw(127)( 98*8-1 downto  97*8), w99 => Pw(127)( 99*8-1 downto  98*8), w100=> Pw(127)(100*8-1 downto  99*8), 
w101=> Pw(127)(101*8-1 downto 100*8), w102=> Pw(127)(102*8-1 downto 101*8), w103=> Pw(127)(103*8-1 downto 102*8), w104=> Pw(127)(104*8-1 downto 103*8), 
w105=> Pw(127)(105*8-1 downto 104*8), w106=> Pw(127)(106*8-1 downto 105*8), w107=> Pw(127)(107*8-1 downto 106*8), w108=> Pw(127)(108*8-1 downto 107*8), 
w109=> Pw(127)(109*8-1 downto 108*8), w110=> Pw(127)(110*8-1 downto 109*8), w111=> Pw(127)(111*8-1 downto 110*8), w112=> Pw(127)(112*8-1 downto 111*8), 
w113=> Pw(127)(113*8-1 downto 112*8), w114=> Pw(127)(114*8-1 downto 113*8), w115=> Pw(127)(115*8-1 downto 114*8), w116=> Pw(127)(116*8-1 downto 115*8), 
w117=> Pw(127)(117*8-1 downto 116*8), w118=> Pw(127)(118*8-1 downto 117*8), w119=> Pw(127)(119*8-1 downto 118*8), w120=> Pw(127)(120*8-1 downto 119*8), 
w121=> Pw(127)(121*8-1 downto 120*8), w122=> Pw(127)(122*8-1 downto 121*8), w123=> Pw(127)(123*8-1 downto 122*8), w124=> Pw(127)(124*8-1 downto 123*8), 
w125=> Pw(127)(125*8-1 downto 124*8), w126=> Pw(127)(126*8-1 downto 125*8), w127=> Pw(127)(127*8-1 downto 126*8), w128=> Pw(127)(128*8-1 downto 127*8), 
           d_out   => pca_d127_out   ,
           en_out  => open  ,
           sof_out => open );


  PCA128_128_inst: PCA_128 
  generic map(
           mult_sum => mult_sum_PCA,
           N        => CL_W,
           M        => PCAweightW,
           in_row   => in_row,
           in_col   => in_col
           )
  port map (
           clk       => clk    ,
           rst       => rst    ,
d01_in    => d01_out, d02_in    => d02_out, d03_in    => d03_out, d04_in    => d04_out, d05_in    => d05_out, d06_in    => d06_out, d07_in    => d07_out, d08_in    => d08_out, d09_in    => d09_out, d10_in    => d10_out, d11_in    => d11_out, d12_in    => d12_out, d13_in    => d13_out, d14_in    => d14_out, d15_in    => d15_out, d16_in    => d16_out, 
d17_in    => d17_out, d18_in    => d18_out, d19_in    => d19_out, d20_in    => d20_out, d21_in    => d21_out, d22_in    => d22_out, d23_in    => d23_out, d24_in    => d24_out, d25_in    => d25_out, d26_in    => d26_out, d27_in    => d27_out, d28_in    => d28_out, d29_in    => d29_out, d30_in    => d30_out, d31_in    => d31_out, d32_in    => d32_out, 
d33_in    => d33_out, d34_in    => d34_out, d35_in    => d35_out, d36_in    => d36_out, d37_in    => d37_out, d38_in    => d38_out, d39_in    => d39_out, d40_in    => d40_out, d41_in    => d41_out, d42_in    => d42_out, d43_in    => d43_out, d44_in    => d44_out, d45_in    => d45_out, d46_in    => d46_out, d47_in    => d47_out, d48_in    => d48_out, 
d49_in    => d49_out, d50_in    => d50_out, d51_in    => d51_out, d52_in    => d52_out, d53_in    => d53_out, d54_in    => d54_out, d55_in    => d55_out, d56_in    => d56_out,d57_in    => d57_out, d58_in    => d58_out, d59_in    => d59_out, d60_in    => d60_out, d61_in    => d61_out, d62_in    => d62_out, d63_in    => d63_out, d64_in    => d64_out, 
d65_in   => d65_out,  d66_in   => d66_out,  d67_in  => d67_out,  d68_in   => d68_out,  d69_in   => d69_out,  d70_in   => d70_out,  d71_in  => d71_out,  d72_in   => d72_out, d73_in   => d73_out,  d74_in   => d74_out,  d75_in  => d75_out,  d76_in   => d76_out,  d77_in   => d77_out,  d78_in   => d78_out,  d79_in  => d79_out,  d80_in   => d80_out, 
d81_in   => d81_out,  d82_in   => d82_out,  d83_in  => d83_out,  d84_in   => d84_out,  d85_in   => d85_out,  d86_in   => d86_out,  d87_in  => d87_out,  d88_in   => d88_out, d89_in   => d89_out,  d90_in   => d90_out,  d91_in  => d91_out,  d92_in   => d92_out,  d93_in   => d93_out,  d94_in   => d94_out,  d95_in  => d95_out,  d96_in   => d96_out, 
d97_in   => d97_out,  d98_in   => d98_out,  d99_in  => d99_out,  d100_in  => d100_out, d101_in  => d101_out, d102_in  => d102_out, d103_in => d103_out, d104_in  => d104_out,d105_in  => d105_out, d106_in  => d106_out, d107_in => d107_out, d108_in  => d108_out, d109_in  => d109_out, d110_in  => d110_out, d111_in => d111_out, d112_in  => d112_out,
d113_in  => d113_out, d114_in  => d114_out, d115_in => d115_out, d116_in  => d116_out, d117_in  => d117_out, d118_in  => d118_out, d119_in => d119_out, d120_in  => d120_out,d121_in  => d121_out, d122_in  => d122_out, d123_in => d123_out, d124_in  => d124_out, d125_in  => d125_out, d126_in  => d126_out, d127_in => d127_out, d128_in  => d128_out,
           en_in     => cl_en_out,
           sof_in    => cl_sof_out,

w01 => Pw(0)(     7 downto    0),   w02 => Pw(0)( 2*8-1 downto    8),   w03 => Pw(0)( 3*8-1 downto  2*8),   w04 => Pw(0)( 4*8-1 downto  3*8),   w05 => Pw(0)( 5*8-1 downto  4*8),   w06 => Pw(0)( 6*8-1 downto  5*8),   w07 => Pw(0)( 7*8-1 downto  6*8),   w08 => Pw(0)( 8*8-1 downto  7*8),  
w09 => Pw(0)( 9*8-1 downto  8*8),   w10 => Pw(0)(10*8-1 downto  9*8),   w11 => Pw(0)(11*8-1 downto 10*8),   w12 => Pw(0)(12*8-1 downto 11*8),   w13 => Pw(0)(13*8-1 downto 12*8),   w14 => Pw(0)(14*8-1 downto 13*8),   w15 => Pw(0)(15*8-1 downto 14*8),   w16 => Pw(0)(16*8-1 downto 15*8),  
w17 => Pw(0)(17*8-1 downto 16*8),   w18 => Pw(0)(18*8-1 downto 17*8),   w19 => Pw(0)(19*8-1 downto 18*8),   w20 => Pw(0)(20*8-1 downto 19*8),   w21 => Pw(0)(21*8-1 downto 20*8),   w22 => Pw(0)(22*8-1 downto 21*8),   w23 => Pw(0)(23*8-1 downto 22*8),   w24 => Pw(0)(24*8-1 downto 23*8),  
w25 => Pw(0)(25*8-1 downto 24*8),   w26 => Pw(0)(26*8-1 downto 25*8),   w27 => Pw(0)(27*8-1 downto 26*8),   w28 => Pw(0)(28*8-1 downto 27*8),   w29 => Pw(0)(29*8-1 downto 28*8),   w30 => Pw(0)(30*8-1 downto 29*8),   w31 => Pw(0)(31*8-1 downto 30*8),   w32 => Pw(0)(32*8-1 downto 31*8),  
w33 => Pw(0)(33*8-1 downto 32*8),   w34 => Pw(0)(34*8-1 downto 33*8),   w35 => Pw(0)(35*8-1 downto 34*8),   w36 => Pw(0)(36*8-1 downto 35*8),   w37 => Pw(0)(37*8-1 downto 36*8),   w38 => Pw(0)(38*8-1 downto 37*8),   w39 => Pw(0)(39*8-1 downto 38*8),   w40 => Pw(0)(40*8-1 downto 39*8),  
w41 => Pw(0)(41*8-1 downto 40*8),   w42 => Pw(0)(42*8-1 downto 41*8),   w43 => Pw(0)(43*8-1 downto 42*8),   w44 => Pw(0)(44*8-1 downto 43*8),   w45 => Pw(0)(45*8-1 downto 44*8),   w46 => Pw(0)(46*8-1 downto 45*8),   w47 => Pw(0)(47*8-1 downto 46*8),   w48 => Pw(0)(48*8-1 downto 47*8),  
w49 => Pw(0)(49*8-1 downto 48*8),   w50 => Pw(0)(50*8-1 downto 49*8),   w51 => Pw(0)(51*8-1 downto 50*8),   w52 => Pw(0)(52*8-1 downto 51*8),   w53 => Pw(0)(53*8-1 downto 52*8),   w54 => Pw(0)(54*8-1 downto 53*8),   w55 => Pw(0)(55*8-1 downto 54*8),   w56 => Pw(0)(56*8-1 downto 55*8),  
w57 => Pw(0)(57*8-1 downto 56*8),   w58 => Pw(0)(58*8-1 downto 57*8),   w59 => Pw(0)(59*8-1 downto 58*8),   w60 => Pw(0)(60*8-1 downto 59*8),   w61 => Pw(0)(61*8-1 downto 60*8),   w62 => Pw(0)(62*8-1 downto 61*8),   w63 => Pw(0)(63*8-1 downto 62*8),   w64 => Pw(0)(64*8-1 downto 63*8), 
w65 => Pw(0)( 65*8-1 downto  64*8), w66 => Pw(0)( 66*8-1 downto  65*8), w67 => Pw(0)( 67*8-1 downto  66*8), w68 => Pw(0)( 68*8-1 downto  67*8), w69 => Pw(0)( 69*8-1 downto  68*8), w70 => Pw(0)( 70*8-1 downto  69*8), w71 => Pw(0)( 71*8-1 downto  70*8), w72 => Pw(0)( 72*8-1 downto  71*8), 
w73 => Pw(0)( 73*8-1 downto  72*8), w74 => Pw(0)( 74*8-1 downto  73*8), w75 => Pw(0)( 75*8-1 downto  74*8), w76 => Pw(0)( 76*8-1 downto  75*8), w77 => Pw(0)( 77*8-1 downto  76*8), w78 => Pw(0)( 78*8-1 downto  77*8), w79 => Pw(0)( 79*8-1 downto  78*8), w80 => Pw(0)( 80*8-1 downto  79*8), 
w81 => Pw(0)( 81*8-1 downto  80*8), w82 => Pw(0)( 82*8-1 downto  81*8), w83 => Pw(0)( 83*8-1 downto  82*8), w84 => Pw(0)( 84*8-1 downto  83*8), w85 => Pw(0)( 85*8-1 downto  84*8), w86 => Pw(0)( 86*8-1 downto  85*8), w87 => Pw(0)( 87*8-1 downto  86*8), w88 => Pw(0)( 88*8-1 downto  87*8), 
w89 => Pw(0)( 89*8-1 downto  88*8), w90 => Pw(0)( 90*8-1 downto  89*8), w91 => Pw(0)( 91*8-1 downto  90*8), w92 => Pw(0)( 92*8-1 downto  91*8), w93 => Pw(0)( 93*8-1 downto  92*8), w94 => Pw(0)( 94*8-1 downto  93*8), w95 => Pw(0)( 95*8-1 downto  94*8), w96 => Pw(0)( 96*8-1 downto  95*8), 
w97 => Pw(0)( 97*8-1 downto  96*8), w98 => Pw(0)( 98*8-1 downto  97*8), w99 => Pw(0)( 99*8-1 downto  98*8), w100=> Pw(0)(100*8-1 downto  99*8), w101=> Pw(0)(101*8-1 downto 100*8), w102=> Pw(0)(102*8-1 downto 101*8), w103=> Pw(0)(103*8-1 downto 102*8), w104=> Pw(0)(104*8-1 downto 103*8), 
w105=> Pw(0)(105*8-1 downto 104*8), w106=> Pw(0)(106*8-1 downto 105*8), w107=> Pw(0)(107*8-1 downto 106*8), w108=> Pw(0)(108*8-1 downto 107*8), w109=> Pw(0)(109*8-1 downto 108*8), w110=> Pw(0)(110*8-1 downto 109*8), w111=> Pw(0)(111*8-1 downto 110*8), w112=> Pw(0)(112*8-1 downto 111*8), 
w113=> Pw(0)(113*8-1 downto 112*8), w114=> Pw(0)(114*8-1 downto 113*8), w115=> Pw(0)(115*8-1 downto 114*8), w116=> Pw(0)(116*8-1 downto 115*8), w117=> Pw(0)(117*8-1 downto 116*8), w118=> Pw(0)(118*8-1 downto 117*8), w119=> Pw(0)(119*8-1 downto 118*8), w120=> Pw(0)(120*8-1 downto 119*8), 
w121=> Pw(0)(121*8-1 downto 120*8), w122=> Pw(0)(122*8-1 downto 121*8), w123=> Pw(0)(123*8-1 downto 122*8), w124=> Pw(0)(124*8-1 downto 123*8), w125=> Pw(0)(125*8-1 downto 124*8), w126=> Pw(0)(126*8-1 downto 125*8), w127=> Pw(0)(127*8-1 downto 126*8), w128=> Pw(0)(128*8-1 downto 127*8), 
           d_out   => pca_d128_out   ,
           en_out  => open  ,
           sof_out => open );



end generate g_PCA_en;

g_PCA_bp: if PCA_en = FALSE generate
   pca_en_out                          <=  cl_en_out;

p_PCA_dis: process (clk)
 begin
    if  rising_edge(clk) then
pca_d01_out(pca_d01_out'left downto pca_d01_out'left - 7) <= d01_out(7 downto 0);
pca_d02_out(pca_d02_out'left downto pca_d02_out'left - 7) <= d02_out(7 downto 0);
pca_d03_out(pca_d03_out'left downto pca_d03_out'left - 7) <= d03_out(7 downto 0);
pca_d04_out(pca_d04_out'left downto pca_d04_out'left - 7) <= d04_out(7 downto 0);
pca_d05_out(pca_d05_out'left downto pca_d05_out'left - 7) <= d05_out(7 downto 0);
pca_d06_out(pca_d06_out'left downto pca_d06_out'left - 7) <= d06_out(7 downto 0);
pca_d07_out(pca_d07_out'left downto pca_d07_out'left - 7) <= d07_out(7 downto 0);
pca_d08_out(pca_d08_out'left downto pca_d08_out'left - 7) <= d08_out(7 downto 0);
pca_d09_out(pca_d09_out'left downto pca_d09_out'left - 7) <= d09_out(7 downto 0);
pca_d10_out(pca_d10_out'left downto pca_d10_out'left - 7) <= d10_out(7 downto 0);
pca_d11_out(pca_d11_out'left downto pca_d11_out'left - 7) <= d11_out(7 downto 0);
pca_d12_out(pca_d12_out'left downto pca_d12_out'left - 7) <= d12_out(7 downto 0);
pca_d13_out(pca_d13_out'left downto pca_d13_out'left - 7) <= d13_out(7 downto 0);
pca_d14_out(pca_d14_out'left downto pca_d14_out'left - 7) <= d14_out(7 downto 0);
pca_d15_out(pca_d15_out'left downto pca_d15_out'left - 7) <= d15_out(7 downto 0);
pca_d16_out(pca_d16_out'left downto pca_d16_out'left - 7) <= d16_out(7 downto 0);
pca_d17_out(pca_d17_out'left downto pca_d17_out'left - 7) <= d17_out(7 downto 0);
pca_d18_out(pca_d18_out'left downto pca_d18_out'left - 7) <= d18_out(7 downto 0);
pca_d19_out(pca_d19_out'left downto pca_d19_out'left - 7) <= d19_out(7 downto 0);
pca_d20_out(pca_d20_out'left downto pca_d20_out'left - 7) <= d20_out(7 downto 0);
pca_d21_out(pca_d21_out'left downto pca_d21_out'left - 7) <= d21_out(7 downto 0);
pca_d22_out(pca_d22_out'left downto pca_d22_out'left - 7) <= d22_out(7 downto 0);
pca_d23_out(pca_d23_out'left downto pca_d23_out'left - 7) <= d23_out(7 downto 0);
pca_d24_out(pca_d24_out'left downto pca_d24_out'left - 7) <= d24_out(7 downto 0);
pca_d25_out(pca_d25_out'left downto pca_d25_out'left - 7) <= d25_out(7 downto 0);
pca_d26_out(pca_d26_out'left downto pca_d26_out'left - 7) <= d26_out(7 downto 0);
pca_d27_out(pca_d27_out'left downto pca_d27_out'left - 7) <= d27_out(7 downto 0);
pca_d28_out(pca_d28_out'left downto pca_d28_out'left - 7) <= d28_out(7 downto 0);
pca_d29_out(pca_d29_out'left downto pca_d29_out'left - 7) <= d29_out(7 downto 0);
pca_d30_out(pca_d30_out'left downto pca_d30_out'left - 7) <= d30_out(7 downto 0);
pca_d31_out(pca_d31_out'left downto pca_d31_out'left - 7) <= d31_out(7 downto 0);
pca_d32_out(pca_d32_out'left downto pca_d32_out'left - 7) <= d32_out(7 downto 0);
pca_d33_out(pca_d33_out'left downto pca_d33_out'left - 7) <= d33_out(7 downto 0);
pca_d34_out(pca_d34_out'left downto pca_d34_out'left - 7) <= d34_out(7 downto 0);
pca_d35_out(pca_d35_out'left downto pca_d35_out'left - 7) <= d35_out(7 downto 0);
pca_d36_out(pca_d36_out'left downto pca_d36_out'left - 7) <= d36_out(7 downto 0);
pca_d37_out(pca_d37_out'left downto pca_d37_out'left - 7) <= d37_out(7 downto 0);
pca_d38_out(pca_d38_out'left downto pca_d38_out'left - 7) <= d38_out(7 downto 0);
pca_d39_out(pca_d39_out'left downto pca_d39_out'left - 7) <= d39_out(7 downto 0);
pca_d40_out(pca_d40_out'left downto pca_d40_out'left - 7) <= d40_out(7 downto 0);
pca_d41_out(pca_d41_out'left downto pca_d41_out'left - 7) <= d41_out(7 downto 0);
pca_d42_out(pca_d42_out'left downto pca_d42_out'left - 7) <= d42_out(7 downto 0);
pca_d43_out(pca_d43_out'left downto pca_d43_out'left - 7) <= d43_out(7 downto 0);
pca_d44_out(pca_d44_out'left downto pca_d44_out'left - 7) <= d44_out(7 downto 0);
pca_d45_out(pca_d45_out'left downto pca_d45_out'left - 7) <= d45_out(7 downto 0);
pca_d46_out(pca_d46_out'left downto pca_d46_out'left - 7) <= d46_out(7 downto 0);
pca_d47_out(pca_d47_out'left downto pca_d47_out'left - 7) <= d47_out(7 downto 0);
pca_d48_out(pca_d48_out'left downto pca_d48_out'left - 7) <= d48_out(7 downto 0);
pca_d49_out(pca_d49_out'left downto pca_d49_out'left - 7) <= d49_out(7 downto 0);
pca_d50_out(pca_d50_out'left downto pca_d50_out'left - 7) <= d50_out(7 downto 0);
pca_d51_out(pca_d51_out'left downto pca_d51_out'left - 7) <= d51_out(7 downto 0);
pca_d52_out(pca_d52_out'left downto pca_d52_out'left - 7) <= d52_out(7 downto 0);
pca_d53_out(pca_d53_out'left downto pca_d53_out'left - 7) <= d53_out(7 downto 0);
pca_d54_out(pca_d54_out'left downto pca_d54_out'left - 7) <= d54_out(7 downto 0);
pca_d55_out(pca_d55_out'left downto pca_d55_out'left - 7) <= d55_out(7 downto 0);
pca_d56_out(pca_d56_out'left downto pca_d56_out'left - 7) <= d56_out(7 downto 0);
pca_d57_out(pca_d57_out'left downto pca_d57_out'left - 7) <= d57_out(7 downto 0);
pca_d58_out(pca_d58_out'left downto pca_d58_out'left - 7) <= d58_out(7 downto 0);
pca_d59_out(pca_d59_out'left downto pca_d59_out'left - 7) <= d59_out(7 downto 0);
pca_d60_out(pca_d60_out'left downto pca_d60_out'left - 7) <= d60_out(7 downto 0);
pca_d61_out(pca_d61_out'left downto pca_d61_out'left - 7) <= d61_out(7 downto 0);
pca_d62_out(pca_d62_out'left downto pca_d62_out'left - 7) <= d62_out(7 downto 0);
pca_d63_out(pca_d63_out'left downto pca_d63_out'left - 7) <= d63_out(7 downto 0);
pca_d64_out(pca_d64_out'left downto pca_d64_out'left - 7) <= d64_out(7 downto 0);

pca_d65_out (pca_d65_out 'left downto pca_d65_out 'left - 7) <= d65_out (7 downto 0);
pca_d66_out (pca_d66_out 'left downto pca_d66_out 'left - 7) <= d66_out (7 downto 0);
pca_d67_out (pca_d67_out 'left downto pca_d67_out 'left - 7) <= d67_out (7 downto 0);
pca_d68_out (pca_d68_out 'left downto pca_d68_out 'left - 7) <= d68_out (7 downto 0);
pca_d69_out (pca_d69_out 'left downto pca_d69_out 'left - 7) <= d69_out (7 downto 0);
pca_d70_out (pca_d70_out 'left downto pca_d70_out 'left - 7) <= d70_out (7 downto 0);
pca_d71_out (pca_d71_out 'left downto pca_d71_out 'left - 7) <= d71_out (7 downto 0);
pca_d72_out (pca_d72_out 'left downto pca_d72_out 'left - 7) <= d72_out (7 downto 0);
pca_d73_out (pca_d73_out 'left downto pca_d73_out 'left - 7) <= d73_out (7 downto 0);
pca_d74_out (pca_d74_out 'left downto pca_d74_out 'left - 7) <= d74_out (7 downto 0);
pca_d75_out (pca_d75_out 'left downto pca_d75_out 'left - 7) <= d75_out (7 downto 0);
pca_d76_out (pca_d76_out 'left downto pca_d76_out 'left - 7) <= d76_out (7 downto 0);
pca_d77_out (pca_d77_out 'left downto pca_d77_out 'left - 7) <= d77_out (7 downto 0);
pca_d78_out (pca_d78_out 'left downto pca_d78_out 'left - 7) <= d78_out (7 downto 0);
pca_d79_out (pca_d79_out 'left downto pca_d79_out 'left - 7) <= d79_out (7 downto 0);
pca_d80_out (pca_d80_out 'left downto pca_d80_out 'left - 7) <= d80_out (7 downto 0);
pca_d81_out (pca_d81_out 'left downto pca_d81_out 'left - 7) <= d81_out (7 downto 0);
pca_d82_out (pca_d82_out 'left downto pca_d82_out 'left - 7) <= d82_out (7 downto 0);
pca_d83_out (pca_d83_out 'left downto pca_d83_out 'left - 7) <= d83_out (7 downto 0);
pca_d84_out (pca_d84_out 'left downto pca_d84_out 'left - 7) <= d84_out (7 downto 0);
pca_d85_out (pca_d85_out 'left downto pca_d85_out 'left - 7) <= d85_out (7 downto 0);
pca_d86_out (pca_d86_out 'left downto pca_d86_out 'left - 7) <= d86_out (7 downto 0);
pca_d87_out (pca_d87_out 'left downto pca_d87_out 'left - 7) <= d87_out (7 downto 0);
pca_d88_out (pca_d88_out 'left downto pca_d88_out 'left - 7) <= d88_out (7 downto 0);
pca_d89_out (pca_d89_out 'left downto pca_d89_out 'left - 7) <= d89_out (7 downto 0);
pca_d90_out (pca_d90_out 'left downto pca_d90_out 'left - 7) <= d90_out (7 downto 0);
pca_d91_out (pca_d91_out 'left downto pca_d91_out 'left - 7) <= d91_out (7 downto 0);
pca_d92_out (pca_d92_out 'left downto pca_d92_out 'left - 7) <= d92_out (7 downto 0);
pca_d93_out (pca_d93_out 'left downto pca_d93_out 'left - 7) <= d93_out (7 downto 0);
pca_d94_out (pca_d94_out 'left downto pca_d94_out 'left - 7) <= d94_out (7 downto 0);
pca_d95_out (pca_d95_out 'left downto pca_d95_out 'left - 7) <= d95_out (7 downto 0);
pca_d96_out (pca_d96_out 'left downto pca_d96_out 'left - 7) <= d96_out (7 downto 0);
pca_d97_out (pca_d97_out 'left downto pca_d97_out 'left - 7) <= d97_out (7 downto 0);
pca_d98_out (pca_d98_out 'left downto pca_d98_out 'left - 7) <= d98_out (7 downto 0);
pca_d99_out (pca_d99_out 'left downto pca_d99_out 'left - 7) <= d99_out (7 downto 0);
pca_d100_out(pca_d100_out'left downto pca_d100_out'left - 7) <= d100_out(7 downto 0);
pca_d101_out(pca_d101_out'left downto pca_d101_out'left - 7) <= d101_out(7 downto 0);
pca_d102_out(pca_d102_out'left downto pca_d102_out'left - 7) <= d102_out(7 downto 0);
pca_d103_out(pca_d103_out'left downto pca_d103_out'left - 7) <= d103_out(7 downto 0);
pca_d104_out(pca_d104_out'left downto pca_d104_out'left - 7) <= d104_out(7 downto 0);
pca_d105_out(pca_d105_out'left downto pca_d105_out'left - 7) <= d105_out(7 downto 0);
pca_d106_out(pca_d106_out'left downto pca_d106_out'left - 7) <= d106_out(7 downto 0);
pca_d107_out(pca_d107_out'left downto pca_d107_out'left - 7) <= d107_out(7 downto 0);
pca_d108_out(pca_d108_out'left downto pca_d108_out'left - 7) <= d108_out(7 downto 0);
pca_d109_out(pca_d109_out'left downto pca_d109_out'left - 7) <= d109_out(7 downto 0);
pca_d110_out(pca_d110_out'left downto pca_d110_out'left - 7) <= d110_out(7 downto 0);
pca_d111_out(pca_d111_out'left downto pca_d111_out'left - 7) <= d111_out(7 downto 0);
pca_d112_out(pca_d112_out'left downto pca_d112_out'left - 7) <= d112_out(7 downto 0);
pca_d113_out(pca_d113_out'left downto pca_d113_out'left - 7) <= d113_out(7 downto 0);
pca_d114_out(pca_d114_out'left downto pca_d114_out'left - 7) <= d114_out(7 downto 0);
pca_d115_out(pca_d115_out'left downto pca_d115_out'left - 7) <= d115_out(7 downto 0);
pca_d116_out(pca_d116_out'left downto pca_d116_out'left - 7) <= d116_out(7 downto 0);
pca_d117_out(pca_d117_out'left downto pca_d117_out'left - 7) <= d117_out(7 downto 0);
pca_d118_out(pca_d118_out'left downto pca_d118_out'left - 7) <= d118_out(7 downto 0);
pca_d119_out(pca_d119_out'left downto pca_d119_out'left - 7) <= d119_out(7 downto 0);
pca_d120_out(pca_d120_out'left downto pca_d120_out'left - 7) <= d120_out(7 downto 0);
pca_d121_out(pca_d121_out'left downto pca_d121_out'left - 7) <= d121_out(7 downto 0);
pca_d122_out(pca_d122_out'left downto pca_d122_out'left - 7) <= d122_out(7 downto 0);
pca_d123_out(pca_d123_out'left downto pca_d123_out'left - 7) <= d123_out(7 downto 0);
pca_d124_out(pca_d124_out'left downto pca_d124_out'left - 7) <= d124_out(7 downto 0);
pca_d125_out(pca_d125_out'left downto pca_d125_out'left - 7) <= d125_out(7 downto 0);
pca_d126_out(pca_d126_out'left downto pca_d126_out'left - 7) <= d126_out(7 downto 0);
pca_d127_out(pca_d127_out'left downto pca_d127_out'left - 7) <= d127_out(7 downto 0);
pca_d128_out(pca_d128_out'left downto pca_d128_out'left - 7) <= d128_out(7 downto 0);

--PCA_dis1 <= d01_out(7 downto 0)+ d02_out(7 downto 0)+ d03_out(7 downto 0)+ d04_out(7 downto 0)+ d05_out(7 downto 0)+ d06_out(7 downto 0)+ d07_out(7 downto 0)+ d08_out(7 downto 0);  
--PCA_dis2 <= d09_out(7 downto 0)+ d10_out(7 downto 0)+ d11_out(7 downto 0)+ d12_out(7 downto 0)+ d13_out(7 downto 0)+ d14_out(7 downto 0)+ d15_out(7 downto 0)+ d16_out(7 downto 0);  
--PCA_dis3 <= d17_out(7 downto 0)+ d18_out(7 downto 0)+ d19_out(7 downto 0)+ d20_out(7 downto 0)+ d21_out(7 downto 0)+ d22_out(7 downto 0)+ d23_out(7 downto 0)+ d24_out(7 downto 0);  
--PCA_dis4 <= d25_out(7 downto 0)+ d26_out(7 downto 0)+ d27_out(7 downto 0)+ d28_out(7 downto 0)+ d29_out(7 downto 0)+ d30_out(7 downto 0)+ d31_out(7 downto 0)+ d32_out(7 downto 0);  
--PCA_dis5 <= d33_out(7 downto 0)+ d34_out(7 downto 0)+ d35_out(7 downto 0)+ d36_out(7 downto 0)+ d37_out(7 downto 0)+ d38_out(7 downto 0)+ d39_out(7 downto 0)+ d40_out(7 downto 0);  
--PCA_dis6 <= d41_out(7 downto 0)+ d42_out(7 downto 0)+ d43_out(7 downto 0)+ d44_out(7 downto 0)+ d45_out(7 downto 0)+ d46_out(7 downto 0)+ d47_out(7 downto 0)+ d48_out(7 downto 0);  
--PCA_dis7 <= d49_out(7 downto 0)+ d50_out(7 downto 0)+ d51_out(7 downto 0)+ d52_out(7 downto 0)+ d53_out(7 downto 0)+ d54_out(7 downto 0)+ d55_out(7 downto 0)+ d56_out(7 downto 0); 
--PCA_dis8 <= d57_out(7 downto 0)+ d58_out(7 downto 0)+ d59_out(7 downto 0)+ d60_out(7 downto 0)+ d61_out(7 downto 0)+ d62_out(7 downto 0)+ d63_out(7 downto 0)+ d64_out(7 downto 0);  
--
-- 
--PCA_dis9  <= d65_out (7 downto 0) + d66_out (7 downto 0) + d67_out (7 downto 0) + d68_out (7 downto 0) + d69_out (7 downto 0) + d70_out (7 downto 0) + d71_out (7 downto 0) + d72_out (7 downto 0);
--PCA_dis10 <= d73_out (7 downto 0) + d74_out (7 downto 0) + d75_out (7 downto 0) + d76_out (7 downto 0) + d77_out (7 downto 0) + d78_out (7 downto 0) + d79_out (7 downto 0) + d80_out (7 downto 0);
--PCA_dis11 <= d81_out (7 downto 0) + d82_out (7 downto 0) + d83_out (7 downto 0) + d84_out (7 downto 0) + d85_out (7 downto 0) + d86_out (7 downto 0) + d87_out (7 downto 0) + d88_out (7 downto 0);
--PCA_dis12 <= d89_out (7 downto 0) + d90_out (7 downto 0) + d91_out (7 downto 0) + d92_out (7 downto 0) + d93_out (7 downto 0) + d94_out (7 downto 0) + d95_out (7 downto 0) + d96_out (7 downto 0);
--PCA_dis13 <= d97_out (7 downto 0) + d98_out (7 downto 0) + d99_out (7 downto 0) + d100_out(7 downto 0) + d101_out(7 downto 0) + d102_out(7 downto 0) + d103_out(7 downto 0) + d104_out(7 downto 0);
--PCA_dis14 <= d105_out(7 downto 0) + d106_out(7 downto 0) + d107_out(7 downto 0) + d108_out(7 downto 0) + d109_out(7 downto 0) + d110_out(7 downto 0) + d111_out(7 downto 0) + d112_out(7 downto 0);
--PCA_dis15 <= d113_out(7 downto 0) + d114_out(7 downto 0) + d115_out(7 downto 0) + d116_out(7 downto 0) + d117_out(7 downto 0) + d118_out(7 downto 0) + d119_out(7 downto 0) + d120_out(7 downto 0);
--PCA_dis16 <= d121_out(7 downto 0) + d122_out(7 downto 0) + d123_out(7 downto 0) + d124_out(7 downto 0) + d125_out(7 downto 0) + d126_out(7 downto 0) + d127_out(7 downto 0) + d128_out(7 downto 0);
--
--pca_d01_out(pca_d01_out'left downto pca_d01_out'left - 7)  <= PCA_dis1 + PCA_dis2 + PCA_dis3 + PCA_dis4 + PCA_dis5 + PCA_dis6 + PCA_dis7 + PCA_dis8 + PCA_dis9  + PCA_dis10 + PCA_dis11 + PCA_dis12 + PCA_dis13 + PCA_dis14 + PCA_dis15 + PCA_dis16;

    end if;
 end process p_PCA_dis;

end generate g_PCA_bp;

--temp connection


-- p_temp: process (clk)
-- begin
--   if  rising_edge(clk) then
--      d_tmp_1_out  <=   pca_d01_out + pca_d09_out + pca_d17_out + pca_d25_out;
--      d_tmp_2_out  <=   pca_d02_out + pca_d10_out + pca_d18_out + pca_d26_out;
--      d_tmp_3_out  <=   pca_d03_out + pca_d11_out + pca_d19_out + pca_d27_out;
--      d_tmp_4_out  <=   pca_d04_out + pca_d12_out + pca_d20_out + pca_d28_out;
--      d_tmp_5_out  <=   pca_d05_out + pca_d13_out + pca_d21_out + pca_d29_out;
--      d_tmp_6_out  <=   pca_d06_out + pca_d14_out + pca_d22_out + pca_d30_out;
--      d_tmp_7_out  <=   pca_d07_out + pca_d15_out + pca_d23_out + pca_d31_out;
--      d_tmp_8_out  <=   pca_d08_out + pca_d16_out + pca_d24_out + pca_d32_out;
--
--      d_tmp_9_out   <=   pca_d33_out + pca_d41_out + pca_d49_out + pca_d57_out;
--      d_tmp_10_out  <=   pca_d34_out + pca_d42_out + pca_d50_out + pca_d58_out;
--      d_tmp_11_out  <=   pca_d35_out + pca_d43_out + pca_d51_out + pca_d59_out;
--      d_tmp_12_out  <=   pca_d36_out + pca_d44_out + pca_d52_out + pca_d60_out;
--      d_tmp_13_out  <=   pca_d37_out + pca_d45_out + pca_d53_out + pca_d61_out;
--      d_tmp_14_out  <=   pca_d38_out + pca_d46_out + pca_d54_out + pca_d62_out;
--      d_tmp_15_out  <=   pca_d39_out + pca_d47_out + pca_d55_out + pca_d63_out;
--      d_tmp_16_out  <=   pca_d40_out + pca_d48_out + pca_d56_out + pca_d64_out;
--
--      d1_out  <=   d_tmp_1_out + d_tmp_9_out   ;
--      d2_out  <=   d_tmp_2_out + d_tmp_10_out  ;
--      d3_out  <=   d_tmp_3_out + d_tmp_11_out  ;
--      d4_out  <=   d_tmp_4_out + d_tmp_12_out  ;
--      d5_out  <=   d_tmp_5_out + d_tmp_13_out  ;
--      d6_out  <=   d_tmp_6_out + d_tmp_14_out  ;
--      d7_out  <=   d_tmp_7_out + d_tmp_15_out  ;
--      d8_out  <=   d_tmp_8_out + d_tmp_16_out  ;
--
--      
--      en_out  <= pca_en_out  ;
--      sof_out <= pca_sof_out ;
--   end if;
-- end process p_temp;

  p_huff1 : process (clk,rst)
  begin
    if rst = '1' then
       h_en        <= '0';
       h_count_en  <= '1';
       h_count_en2 <= '0';
       h_count     <= (others => '0');
    elsif rising_edge(clk) then
       if h_count_en = '1' then
          --h_num   <= h_count;
          h_count <= h_count + 1;
       end if;
       if h_count = 255 then
          h_count_en <= '0';
       end if;
       h_count_en2 <= h_count_en;
       h_en        <= h_count_en2;
    end if;
  end process p_huff1;

  p_huff2 : process (clk)
  begin
    if rising_edge(clk) then
       alpha_data  <=                                h_count  ;
       alpha_code  <=  Huff_code (conv_integer("0" & h_count));
       alpha_width <=  Huff_width(conv_integer("0" & h_count));
    end if;
  end process p_huff2;


Huffman128_inst: Huffman128 
  generic map(
           N           => 8          ,  -- input data width
           M           => Huff_wid   ,  -- max code width
           Wh          => Wh         ,
           Wb          => Wb         ,
           Huff_enc_en => Huff_enc_en,
           depth       => depth      ,
           burst       => burst
           )
  port map (
           clk      => clk  ,
           rst      => rst  , 

           init_en        => h_en       ,
           alpha_data     => alpha_data ,   
           alpha_code     => alpha_code ,    
           alpha_width    => alpha_width,

           d01_in         => pca_d01_out(pca_d01_out'left downto pca_d01_out'left - 7),
           d02_in         => pca_d02_out(pca_d02_out'left downto pca_d02_out'left - 7),
           d03_in         => pca_d03_out(pca_d03_out'left downto pca_d03_out'left - 7),
           d04_in         => pca_d04_out(pca_d04_out'left downto pca_d04_out'left - 7),
           d05_in         => pca_d05_out(pca_d05_out'left downto pca_d05_out'left - 7),
           d06_in         => pca_d06_out(pca_d06_out'left downto pca_d06_out'left - 7),
           d07_in         => pca_d07_out(pca_d07_out'left downto pca_d07_out'left - 7),
           d08_in         => pca_d08_out(pca_d08_out'left downto pca_d08_out'left - 7),
           d09_in         => pca_d09_out(pca_d09_out'left downto pca_d09_out'left - 7),
           d10_in         => pca_d10_out(pca_d10_out'left downto pca_d10_out'left - 7),
           d11_in         => pca_d11_out(pca_d11_out'left downto pca_d11_out'left - 7),
           d12_in         => pca_d12_out(pca_d12_out'left downto pca_d12_out'left - 7),
           d13_in         => pca_d13_out(pca_d13_out'left downto pca_d13_out'left - 7),
           d14_in         => pca_d14_out(pca_d14_out'left downto pca_d14_out'left - 7),
           d15_in         => pca_d15_out(pca_d15_out'left downto pca_d15_out'left - 7),
           d16_in         => pca_d16_out(pca_d16_out'left downto pca_d16_out'left - 7),
           d17_in         => pca_d17_out(pca_d17_out'left downto pca_d17_out'left - 7),
           d18_in         => pca_d18_out(pca_d18_out'left downto pca_d18_out'left - 7),
           d19_in         => pca_d19_out(pca_d19_out'left downto pca_d19_out'left - 7),
           d20_in         => pca_d20_out(pca_d20_out'left downto pca_d20_out'left - 7),
           d21_in         => pca_d21_out(pca_d21_out'left downto pca_d21_out'left - 7),
           d22_in         => pca_d22_out(pca_d22_out'left downto pca_d22_out'left - 7),
           d23_in         => pca_d23_out(pca_d23_out'left downto pca_d23_out'left - 7),
           d24_in         => pca_d24_out(pca_d24_out'left downto pca_d24_out'left - 7),
           d25_in         => pca_d25_out(pca_d25_out'left downto pca_d25_out'left - 7),
           d26_in         => pca_d26_out(pca_d26_out'left downto pca_d26_out'left - 7),
           d27_in         => pca_d27_out(pca_d27_out'left downto pca_d27_out'left - 7),
           d28_in         => pca_d28_out(pca_d28_out'left downto pca_d28_out'left - 7),
           d29_in         => pca_d29_out(pca_d29_out'left downto pca_d29_out'left - 7),
           d30_in         => pca_d30_out(pca_d30_out'left downto pca_d30_out'left - 7),
           d31_in         => pca_d31_out(pca_d31_out'left downto pca_d31_out'left - 7),
           d32_in         => pca_d32_out(pca_d32_out'left downto pca_d32_out'left - 7),
           d33_in         => pca_d33_out(pca_d33_out'left downto pca_d33_out'left - 7),
           d34_in         => pca_d34_out(pca_d34_out'left downto pca_d34_out'left - 7),
           d35_in         => pca_d35_out(pca_d35_out'left downto pca_d35_out'left - 7),
           d36_in         => pca_d36_out(pca_d36_out'left downto pca_d36_out'left - 7),
           d37_in         => pca_d37_out(pca_d37_out'left downto pca_d37_out'left - 7),
           d38_in         => pca_d38_out(pca_d38_out'left downto pca_d38_out'left - 7),
           d39_in         => pca_d39_out(pca_d39_out'left downto pca_d39_out'left - 7),
           d40_in         => pca_d40_out(pca_d40_out'left downto pca_d40_out'left - 7),
           d41_in         => pca_d41_out(pca_d41_out'left downto pca_d41_out'left - 7),
           d42_in         => pca_d42_out(pca_d42_out'left downto pca_d42_out'left - 7),
           d43_in         => pca_d43_out(pca_d43_out'left downto pca_d43_out'left - 7),
           d44_in         => pca_d44_out(pca_d44_out'left downto pca_d44_out'left - 7),
           d45_in         => pca_d45_out(pca_d45_out'left downto pca_d45_out'left - 7),
           d46_in         => pca_d46_out(pca_d46_out'left downto pca_d46_out'left - 7),
           d47_in         => pca_d47_out(pca_d47_out'left downto pca_d47_out'left - 7),
           d48_in         => pca_d48_out(pca_d48_out'left downto pca_d48_out'left - 7),
           d49_in         => pca_d49_out(pca_d49_out'left downto pca_d49_out'left - 7),
           d50_in         => pca_d50_out(pca_d50_out'left downto pca_d50_out'left - 7),
           d51_in         => pca_d51_out(pca_d51_out'left downto pca_d51_out'left - 7),
           d52_in         => pca_d52_out(pca_d52_out'left downto pca_d52_out'left - 7),
           d53_in         => pca_d53_out(pca_d53_out'left downto pca_d53_out'left - 7),
           d54_in         => pca_d54_out(pca_d54_out'left downto pca_d54_out'left - 7),
           d55_in         => pca_d55_out(pca_d55_out'left downto pca_d55_out'left - 7),
           d56_in         => pca_d56_out(pca_d56_out'left downto pca_d56_out'left - 7),
           d57_in         => pca_d57_out(pca_d57_out'left downto pca_d57_out'left - 7),
           d58_in         => pca_d58_out(pca_d58_out'left downto pca_d58_out'left - 7),
           d59_in         => pca_d59_out(pca_d59_out'left downto pca_d59_out'left - 7),
           d60_in         => pca_d60_out(pca_d60_out'left downto pca_d60_out'left - 7),
           d61_in         => pca_d61_out(pca_d61_out'left downto pca_d61_out'left - 7),
           d62_in         => pca_d62_out(pca_d62_out'left downto pca_d62_out'left - 7),
           d63_in         => pca_d63_out(pca_d63_out'left downto pca_d63_out'left - 7),
           d64_in         => pca_d64_out(pca_d64_out'left downto pca_d64_out'left - 7),

           d65_in          => pca_d65_out (pca_d65_out'left  downto pca_d65_out'left  - 7),
           d66_in          => pca_d66_out (pca_d66_out'left  downto pca_d66_out'left  - 7),
           d67_in          => pca_d67_out (pca_d67_out'left  downto pca_d67_out'left  - 7),
           d68_in          => pca_d68_out (pca_d68_out'left  downto pca_d68_out'left  - 7),
           d69_in          => pca_d69_out (pca_d69_out'left  downto pca_d69_out'left  - 7),
           d70_in          => pca_d70_out (pca_d70_out'left  downto pca_d70_out'left  - 7),
           d71_in          => pca_d71_out (pca_d71_out'left  downto pca_d71_out'left  - 7),
           d72_in          => pca_d72_out (pca_d72_out'left  downto pca_d72_out'left  - 7),
           d73_in          => pca_d73_out (pca_d73_out'left  downto pca_d73_out'left  - 7),
           d74_in          => pca_d74_out (pca_d74_out'left  downto pca_d74_out'left  - 7),
           d75_in          => pca_d75_out (pca_d75_out'left  downto pca_d75_out'left  - 7),
           d76_in          => pca_d76_out (pca_d76_out'left  downto pca_d76_out'left  - 7),
           d77_in          => pca_d77_out (pca_d77_out'left  downto pca_d77_out'left  - 7),
           d78_in          => pca_d78_out (pca_d78_out'left  downto pca_d78_out'left  - 7),
           d79_in          => pca_d79_out (pca_d79_out'left  downto pca_d79_out'left  - 7),
           d80_in          => pca_d80_out (pca_d80_out'left  downto pca_d80_out'left  - 7),
           d81_in          => pca_d81_out (pca_d81_out'left  downto pca_d81_out'left  - 7),
           d82_in          => pca_d82_out (pca_d82_out'left  downto pca_d82_out'left  - 7),
           d83_in          => pca_d83_out (pca_d83_out'left  downto pca_d83_out'left  - 7),
           d84_in          => pca_d84_out (pca_d84_out'left  downto pca_d84_out'left  - 7),
           d85_in          => pca_d85_out (pca_d85_out'left  downto pca_d85_out'left  - 7),
           d86_in          => pca_d86_out (pca_d86_out'left  downto pca_d86_out'left  - 7),
           d87_in          => pca_d87_out (pca_d87_out'left  downto pca_d87_out'left  - 7),
           d88_in          => pca_d88_out (pca_d88_out'left  downto pca_d88_out'left  - 7),
           d89_in          => pca_d89_out (pca_d89_out'left  downto pca_d89_out'left  - 7),
           d90_in          => pca_d90_out (pca_d90_out'left  downto pca_d90_out'left  - 7),
           d91_in          => pca_d91_out (pca_d91_out'left  downto pca_d91_out'left  - 7),
           d92_in          => pca_d92_out (pca_d92_out'left  downto pca_d92_out'left  - 7),
           d93_in          => pca_d93_out (pca_d93_out'left  downto pca_d93_out'left  - 7),
           d94_in          => pca_d94_out (pca_d94_out'left  downto pca_d94_out'left  - 7),
           d95_in          => pca_d95_out (pca_d95_out'left  downto pca_d95_out'left  - 7),
           d96_in          => pca_d96_out (pca_d96_out'left  downto pca_d96_out'left  - 7),
           d97_in          => pca_d97_out (pca_d97_out'left  downto pca_d97_out'left  - 7),
           d98_in          => pca_d98_out (pca_d98_out'left  downto pca_d98_out'left  - 7),
           d99_in          => pca_d99_out (pca_d99_out'left  downto pca_d99_out'left  - 7),
           d100_in         => pca_d100_out(pca_d100_out'left downto pca_d100_out'left - 7),
           d101_in         => pca_d101_out(pca_d101_out'left downto pca_d101_out'left - 7),
           d102_in         => pca_d102_out(pca_d102_out'left downto pca_d102_out'left - 7),
           d103_in         => pca_d103_out(pca_d103_out'left downto pca_d103_out'left - 7),
           d104_in         => pca_d104_out(pca_d104_out'left downto pca_d104_out'left - 7),
           d105_in         => pca_d105_out(pca_d105_out'left downto pca_d105_out'left - 7),
           d106_in         => pca_d106_out(pca_d106_out'left downto pca_d106_out'left - 7),
           d107_in         => pca_d107_out(pca_d107_out'left downto pca_d107_out'left - 7),
           d108_in         => pca_d108_out(pca_d108_out'left downto pca_d108_out'left - 7),
           d109_in         => pca_d109_out(pca_d109_out'left downto pca_d109_out'left - 7),
           d110_in         => pca_d110_out(pca_d110_out'left downto pca_d110_out'left - 7),
           d111_in         => pca_d111_out(pca_d111_out'left downto pca_d111_out'left - 7),
           d112_in         => pca_d112_out(pca_d112_out'left downto pca_d112_out'left - 7),
           d113_in         => pca_d113_out(pca_d113_out'left downto pca_d113_out'left - 7),
           d114_in         => pca_d114_out(pca_d114_out'left downto pca_d114_out'left - 7),
           d115_in         => pca_d115_out(pca_d115_out'left downto pca_d115_out'left - 7),
           d116_in         => pca_d116_out(pca_d116_out'left downto pca_d116_out'left - 7),
           d117_in         => pca_d117_out(pca_d117_out'left downto pca_d117_out'left - 7),
           d118_in         => pca_d118_out(pca_d118_out'left downto pca_d118_out'left - 7),
           d119_in         => pca_d119_out(pca_d119_out'left downto pca_d119_out'left - 7),
           d120_in         => pca_d120_out(pca_d120_out'left downto pca_d120_out'left - 7),
           d121_in         => pca_d121_out(pca_d121_out'left downto pca_d121_out'left - 7),
           d122_in         => pca_d122_out(pca_d122_out'left downto pca_d122_out'left - 7),
           d123_in         => pca_d123_out(pca_d123_out'left downto pca_d123_out'left - 7),
           d124_in         => pca_d124_out(pca_d124_out'left downto pca_d124_out'left - 7),
           d125_in         => pca_d125_out(pca_d125_out'left downto pca_d125_out'left - 7),
           d126_in         => pca_d126_out(pca_d126_out'left downto pca_d126_out'left - 7),
           d127_in         => pca_d127_out(pca_d127_out'left downto pca_d127_out'left - 7),
           d128_in         => pca_d128_out(pca_d128_out'left downto pca_d128_out'left - 7),

           en_in          => pca_en_out,        --
           sof_in         => pca_sof_out,        --                         -- start of frame
           eof_in         => '0',        --                         -- end of frame

           buf_rd        => buf_rd         ,
           buf_num       => buf_num        ,
           d_out         => huff_out       ,
           en_out        => open           ,
           eof_out       => open           );                        -- huffman codde output

    d_out  <=  huff_out;


-- PCA weights

    
--  p_pca_w : process (clk,rst)
--  begin
--    if rst = '1' then
--       pca_w_addr      <= (others => '0');
--       pca_col_count   <= (others => '0');
--       --pca_w_init      <= '1';
--    elsif rising_edge(clk) then
--       --pca_w_init      <= '0';
--       --if pca_w_init = '1' or ( cl_en_out = '1' and pca_w_addr = std_logic_vector(to_unsigned(in_col, pca_w_addr'length))) then
--       if cl_en_out = '1' and pca_col_count = std_logic_vector(to_unsigned(in_col-1, pca_w_addr'length)) then
--          pca_w_addr <= pca_w_addr + 1;
--       end if;
--
--       if cl_en_out = '1'  then
--          if pca_col_count = std_logic_vector(to_unsigned(in_col-1, pca_w_addr'length)) then
--             pca_col_count   <= (others => '0');
--          else
--             pca_col_count <= pca_col_count + 1;
--          end if;
--       end if;
--    end if;
--  end process p_pca_w;

--  p_pca_w2 : process (clk)
--  begin
--    if rising_edge(clk) then
--      pca_w_data <= PCAweight64(conv_integer("0" & pca_w_addr));
--    end if;
--  end process p_pca_w2;
--pca_w01 <= pca_w_data(   8-1 downto    0); 
--pca_w02 <= pca_w_data( 2*8-1 downto    8); 
--pca_w03 <= pca_w_data( 3*8-1 downto  2*8); 
--pca_w04 <= pca_w_data( 4*8-1 downto  3*8); 
--pca_w05 <= pca_w_data( 5*8-1 downto  4*8); 
--pca_w06 <= pca_w_data( 6*8-1 downto  5*8); 
--pca_w07 <= pca_w_data( 7*8-1 downto  6*8); 
--pca_w08 <= pca_w_data( 8*8-1 downto  7*8); 
--pca_w09 <= pca_w_data( 9*8-1 downto  8*8); 
--pca_w10 <= pca_w_data(10*8-1 downto  9*8); 
--pca_w11 <= pca_w_data(11*8-1 downto 10*8); 
--pca_w12 <= pca_w_data(12*8-1 downto 11*8); 
--pca_w13 <= pca_w_data(13*8-1 downto 12*8); 
--pca_w14 <= pca_w_data(14*8-1 downto 13*8); 
--pca_w15 <= pca_w_data(15*8-1 downto 14*8); 
--pca_w16 <= pca_w_data(16*8-1 downto 15*8); 
--pca_w17 <= pca_w_data(17*8-1 downto 16*8); 
--pca_w18 <= pca_w_data(18*8-1 downto 17*8); 
--pca_w19 <= pca_w_data(19*8-1 downto 18*8); 
--pca_w20 <= pca_w_data(20*8-1 downto 19*8); 
--pca_w21 <= pca_w_data(21*8-1 downto 20*8); 
--pca_w22 <= pca_w_data(22*8-1 downto 21*8); 
--pca_w23 <= pca_w_data(23*8-1 downto 22*8); 
--pca_w24 <= pca_w_data(24*8-1 downto 23*8); 
--pca_w25 <= pca_w_data(25*8-1 downto 24*8); 
--pca_w26 <= pca_w_data(26*8-1 downto 25*8); 
--pca_w27 <= pca_w_data(27*8-1 downto 26*8); 
--pca_w28 <= pca_w_data(28*8-1 downto 27*8); 
--pca_w29 <= pca_w_data(29*8-1 downto 28*8); 
--pca_w30 <= pca_w_data(30*8-1 downto 29*8); 
--pca_w31 <= pca_w_data(31*8-1 downto 30*8); 
--pca_w32 <= pca_w_data(32*8-1 downto 31*8); 
--pca_w33 <= pca_w_data(33*8-1 downto 32*8); 
--pca_w34 <= pca_w_data(34*8-1 downto 33*8); 
--pca_w35 <= pca_w_data(35*8-1 downto 34*8); 
--pca_w36 <= pca_w_data(36*8-1 downto 35*8); 
--pca_w37 <= pca_w_data(37*8-1 downto 36*8); 
--pca_w38 <= pca_w_data(38*8-1 downto 37*8); 
--pca_w39 <= pca_w_data(39*8-1 downto 38*8); 
--pca_w40 <= pca_w_data(40*8-1 downto 39*8); 
--pca_w41 <= pca_w_data(41*8-1 downto 40*8); 
--pca_w42 <= pca_w_data(42*8-1 downto 41*8); 
--pca_w43 <= pca_w_data(43*8-1 downto 42*8); 
--pca_w44 <= pca_w_data(44*8-1 downto 43*8); 
--pca_w45 <= pca_w_data(45*8-1 downto 44*8); 
--pca_w46 <= pca_w_data(46*8-1 downto 45*8); 
--pca_w47 <= pca_w_data(47*8-1 downto 46*8); 
--pca_w48 <= pca_w_data(48*8-1 downto 47*8); 
--pca_w49 <= pca_w_data(49*8-1 downto 48*8); 
--pca_w50 <= pca_w_data(50*8-1 downto 49*8); 
--pca_w51 <= pca_w_data(51*8-1 downto 50*8); 
--pca_w52 <= pca_w_data(52*8-1 downto 51*8); 
--pca_w53 <= pca_w_data(53*8-1 downto 52*8); 
--pca_w54 <= pca_w_data(54*8-1 downto 53*8); 
--pca_w55 <= pca_w_data(55*8-1 downto 54*8); 
--pca_w56 <= pca_w_data(56*8-1 downto 55*8); 
--pca_w57 <= pca_w_data(57*8-1 downto 56*8); 
--pca_w58 <= pca_w_data(58*8-1 downto 57*8); 
--pca_w59 <= pca_w_data(59*8-1 downto 58*8); 
--pca_w60 <= pca_w_data(60*8-1 downto 59*8); 
--pca_w61 <= pca_w_data(61*8-1 downto 60*8); 
--pca_w62 <= pca_w_data(62*8-1 downto 61*8); 
--pca_w63 <= pca_w_data(63*8-1 downto 62*8); 
--pca_w64 <= pca_w_data(64*8-1 downto 63*8); 

end a;