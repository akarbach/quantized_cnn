library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity ConvLayersNxM is
  generic (
  	       mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width      (Note, W+SR <= N+M+4)
           SR            : integer := 2; -- data shift right before output
  	       in_row        : integer := 256;
  	       in_col        : integer := 256
  	       );
  port    (
           clk     : in std_logic;
           rst     : in std_logic;
  	       d_in    : in std_logic_vector (N-1 downto 0);
  	       en_in   : in std_logic;
  	       sof_in  : in std_logic; -- start of frame

           w_d     : in std_logic_vector(M-1 downto 0); -- weight data
           w_a     : in std_logic_vector(9 downto 0);   -- weight address
           w_en    : in std_logic;                      -- weight en

           max0_out   : out std_logic_vector (W-1 downto 0);
           max1_out   : out std_logic_vector (W-1 downto 0);
           max2_out   : out std_logic_vector (W-1 downto 0);
           max3_out   : out std_logic_vector (W-1 downto 0);
           max4_out   : out std_logic_vector (W-1 downto 0);
           max5_out   : out std_logic_vector (W-1 downto 0);
           max6_out   : out std_logic_vector (W-1 downto 0);
           max7_out   : out std_logic_vector (W-1 downto 0);
           max8_out   : out std_logic_vector (W-1 downto 0);
           max9_out   : out std_logic_vector (W-1 downto 0);
           en_out  : out std_logic
           );
end ConvLayersNxM;

architecture a of ConvLayersNxM is

component ConvLayersN is
  generic (
           mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width      (Note, W+SR <= N+M+4)
           SR            : integer := 2; -- data shift right before output
           in_row        : integer := 256;
           in_col        : integer := 256
           );
  port    (
           clk     : in std_logic;
           rst     : in std_logic;
           d_in    : in std_logic_vector (N-1 downto 0);
           en_in   : in std_logic;
           sof_in  : in std_logic; -- start of frame

           w01      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w02      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w03      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w04      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w05      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w06      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w07      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w08      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w09      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w11      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w12      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w13      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w14      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w15      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w16      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w17      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w18      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w19      : in std_logic_vector(M-1 downto 0); -- weight matrix


           w21      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w22      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w23      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w24      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w25      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w26      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w27      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w28      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w29      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w31      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w32      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w33      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w34      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w35      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w36      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w37      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w38      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w39      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w41      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w42      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w43      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w44      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w45      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w46      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w47      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w48      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w49      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w51      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w52      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w53      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w54      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w55      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w56      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w57      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w58      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w59      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w61      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w62      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w63      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w64      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w65      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w66      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w67      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w68      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w69      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w71      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w72      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w73      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w74      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w75      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w76      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w77      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w78      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w79      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w81      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w82      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w83      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w84      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w85      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w86      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w87      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w88      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w89      : in std_logic_vector(M-1 downto 0); -- weight matrix

           w91      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w92      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w93      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w94      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w95      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w96      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w97      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w98      : in std_logic_vector(M-1 downto 0); -- weight matrix
           w99      : in std_logic_vector(M-1 downto 0); -- weight matrix
           d_out   : out std_logic_vector (W-1 downto 0);
           en_out  : out std_logic;
           sof_out : out std_logic);
end component;

signal           w001      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w002      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w003      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w004      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w005      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w006      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w007      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w008      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w009      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w011      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w012      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w013      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w014      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w015      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w016      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w017      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w018      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w019      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w021      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w022      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w023      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w024      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w025      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w026      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w027      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w028      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w029      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w031      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w032      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w033      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w034      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w035      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w036      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w037      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w038      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w039      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w041      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w042      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w043      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w044      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w045      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w046      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w047      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w048      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w049      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w051      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w052      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w053      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w054      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w055      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w056      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w057      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w058      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w059      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w061      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w062      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w063      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w064      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w065      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w066      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w067      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w068      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w069      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w071      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w072      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w073      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w074      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w075      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w076      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w077      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w078      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w079      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w081      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w082      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w083      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w084      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w085      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w086      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w087      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w088      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w089      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w091      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w092      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w093      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w094      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w095      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w096      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w097      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w098      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w099      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w101      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w102      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w103      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w104      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w105      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w106      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w107      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w108      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w109      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w111      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w112      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w113      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w114      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w115      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w116      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w117      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w118      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w119      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w121      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w122      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w123      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w124      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w125      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w126      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w127      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w128      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w129      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w131      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w132      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w133      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w134      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w135      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w136      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w137      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w138      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w139      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w141      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w142      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w143      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w144      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w145      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w146      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w147      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w148      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w149      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w151      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w152      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w153      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w154      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w155      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w156      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w157      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w158      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w159      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w161      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w162      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w163      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w164      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w165      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w166      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w167      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w168      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w169      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w171      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w172      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w173      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w174      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w175      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w176      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w177      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w178      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w179      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w181      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w182      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w183      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w184      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w185      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w186      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w187      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w188      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w189      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w191      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w192      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w193      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w194      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w195      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w196      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w197      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w198      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w199      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w201      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w202      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w203      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w204      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w205      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w206      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w207      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w208      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w209      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w211      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w212      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w213      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w214      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w215      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w216      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w217      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w218      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w219      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w221      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w222      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w223      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w224      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w225      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w226      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w227      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w228      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w229      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w231      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w232      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w233      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w234      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w235      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w236      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w237      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w238      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w239      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w241      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w242      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w243      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w244      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w245      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w246      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w247      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w248      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w249      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w251      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w252      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w253      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w254      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w255      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w256      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w257      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w258      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w259      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w261      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w262      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w263      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w264      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w265      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w266      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w267      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w268      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w269      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w271      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w272      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w273      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w274      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w275      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w276      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w277      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w278      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w279      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w281      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w282      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w283      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w284      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w285      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w286      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w287      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w288      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w289      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w291      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w292      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w293      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w294      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w295      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w296      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w297      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w298      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w299      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w301      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w302      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w303      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w304      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w305      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w306      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w307      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w308      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w309      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w311      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w312      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w313      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w314      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w315      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w316      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w317      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w318      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w319      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w321      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w322      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w323      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w324      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w325      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w326      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w327      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w328      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w329      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w331      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w332      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w333      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w334      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w335      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w336      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w337      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w338      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w339      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w341      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w342      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w343      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w344      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w345      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w346      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w347      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w348      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w349      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w351      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w352      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w353      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w354      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w355      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w356      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w357      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w358      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w359      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w361      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w362      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w363      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w364      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w365      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w366      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w367      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w368      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w369      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w371      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w372      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w373      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w374      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w375      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w376      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w377      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w378      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w379      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w381      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w382      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w383      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w384      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w385      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w386      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w387      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w388      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w389      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w391      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w392      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w393      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w394      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w395      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w396      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w397      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w398      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w399      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w401      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w402      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w403      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w404      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w405      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w406      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w407      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w408      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w409      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w411      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w412      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w413      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w414      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w415      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w416      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w417      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w418      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w419      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w421      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w422      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w423      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w424      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w425      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w426      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w427      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w428      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w429      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w431      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w432      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w433      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w434      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w435      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w436      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w437      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w438      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w439      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w441      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w442      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w443      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w444      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w445      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w446      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w447      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w448      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w449      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w451      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w452      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w453      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w454      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w455      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w456      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w457      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w458      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w459      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w461      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w462      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w463      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w464      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w465      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w466      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w467      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w468      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w469      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w471      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w472      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w473      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w474      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w475      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w476      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w477      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w478      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w479      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w481      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w482      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w483      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w484      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w485      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w486      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w487      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w488      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w489      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w491      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w492      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w493      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w494      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w495      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w496      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w497      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w498      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w499      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w501      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w502      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w503      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w504      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w505      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w506      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w507      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w508      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w509      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w511      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w512      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w513      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w514      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w515      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w516      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w517      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w518      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w519      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w521      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w522      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w523      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w524      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w525      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w526      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w527      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w528      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w529      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w531      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w532      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w533      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w534      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w535      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w536      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w537      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w538      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w539      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w541      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w542      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w543      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w544      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w545      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w546      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w547      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w548      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w549      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w551      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w552      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w553      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w554      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w555      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w556      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w557      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w558      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w559      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w561      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w562      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w563      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w564      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w565      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w566      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w567      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w568      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w569      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w571      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w572      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w573      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w574      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w575      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w576      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w577      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w578      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w579      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w581      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w582      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w583      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w584      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w585      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w586      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w587      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w588      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w589      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w591      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w592      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w593      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w594      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w595      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w596      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w597      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w598      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w599      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w601      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w602      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w603      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w604      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w605      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w606      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w607      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w608      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w609      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w611      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w612      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w613      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w614      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w615      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w616      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w617      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w618      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w619      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w621      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w622      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w623      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w624      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w625      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w626      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w627      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w628      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w629      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w631      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w632      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w633      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w634      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w635      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w636      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w637      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w638      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w639      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w641      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w642      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w643      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w644      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w645      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w646      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w647      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w648      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w649      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w651      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w652      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w653      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w654      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w655      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w656      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w657      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w658      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w659      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w661      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w662      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w663      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w664      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w665      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w666      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w667      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w668      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w669      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w671      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w672      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w673      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w674      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w675      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w676      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w677      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w678      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w679      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w681      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w682      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w683      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w684      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w685      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w686      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w687      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w688      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w689      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w691      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w692      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w693      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w694      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w695      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w696      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w697      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w698      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w699      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w701      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w702      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w703      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w704      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w705      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w706      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w707      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w708      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w709      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w711      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w712      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w713      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w714      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w715      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w716      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w717      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w718      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w719      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w721      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w722      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w723      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w724      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w725      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w726      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w727      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w728      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w729      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w731      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w732      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w733      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w734      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w735      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w736      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w737      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w738      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w739      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w741      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w742      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w743      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w744      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w745      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w746      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w747      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w748      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w749      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w751      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w752      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w753      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w754      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w755      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w756      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w757      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w758      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w759      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w761      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w762      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w763      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w764      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w765      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w766      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w767      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w768      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w769      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w771      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w772      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w773      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w774      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w775      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w776      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w777      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w778      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w779      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w781      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w782      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w783      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w784      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w785      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w786      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w787      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w788      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w789      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w791      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w792      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w793      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w794      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w795      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w796      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w797      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w798      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w799      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w801      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w802      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w803      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w804      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w805      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w806      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w807      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w808      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w809      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w811      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w812      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w813      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w814      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w815      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w816      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w817      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w818      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w819      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w821      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w822      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w823      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w824      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w825      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w826      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w827      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w828      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w829      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w831      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w832      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w833      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w834      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w835      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w836      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w837      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w838      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w839      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w841      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w842      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w843      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w844      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w845      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w846      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w847      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w848      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w849      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w851      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w852      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w853      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w854      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w855      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w856      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w857      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w858      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w859      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w861      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w862      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w863      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w864      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w865      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w866      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w867      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w868      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w869      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w871      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w872      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w873      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w874      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w875      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w876      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w877      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w878      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w879      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w881      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w882      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w883      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w884      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w885      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w886      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w887      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w888      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w889      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w891      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w892      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w893      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w894      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w895      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w896      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w897      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w898      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w899      : std_logic_vector(M-1 downto 0); -- weight matrix


signal           w901      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w902      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w903      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w904      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w905      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w906      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w907      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w908      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w909      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w911      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w912      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w913      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w914      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w915      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w916      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w917      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w918      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w919      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w921      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w922      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w923      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w924      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w925      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w926      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w927      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w928      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w929      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w931      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w932      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w933      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w934      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w935      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w936      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w937      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w938      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w939      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w941      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w942      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w943      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w944      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w945      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w946      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w947      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w948      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w949      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w951      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w952      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w953      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w954      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w955      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w956      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w957      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w958      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w959      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w961      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w962      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w963      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w964      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w965      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w966      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w967      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w968      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w969      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w971      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w972      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w973      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w974      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w975      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w976      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w977      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w978      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w979      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w981      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w982      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w983      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w984      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w985      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w986      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w987      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w988      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w989      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w991      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w992      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w993      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w994      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w995      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w996      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w997      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w998      : std_logic_vector(M-1 downto 0); -- weight matrix
signal           w999      : std_logic_vector(M-1 downto 0); -- weight matrix

signal     d0   : std_logic_vector (W-1 downto 0);
signal     d1   : std_logic_vector (W-1 downto 0);
signal     d2   : std_logic_vector (W-1 downto 0);
signal     d3   : std_logic_vector (W-1 downto 0);
signal     d4   : std_logic_vector (W-1 downto 0);
signal     d5   : std_logic_vector (W-1 downto 0);
signal     d6   : std_logic_vector (W-1 downto 0);
signal     d7   : std_logic_vector (W-1 downto 0);
signal     d8   : std_logic_vector (W-1 downto 0);
signal     d9   : std_logic_vector (W-1 downto 0);
signal     en0  : std_logic;
signal     en1  : std_logic;
signal     en2  : std_logic;
signal     en3  : std_logic;
signal     en4  : std_logic;
signal     en5  : std_logic;
signal     en6  : std_logic;
signal     en7  : std_logic;
signal     en8  : std_logic;
signal     en9  : std_logic;
signal     sof0 : std_logic;
signal     sof1 : std_logic;
signal     sof2 : std_logic;
signal     sof3 : std_logic;
signal     sof4 : std_logic;
signal     sof5 : std_logic;
signal     sof6 : std_logic;
signal     sof7 : std_logic;
signal     sof8 : std_logic;
signal     sof9 : std_logic;

signal w_a2  : natural range 0 to 1023 ;
signal w_d2  : std_logic_vector(M-1 downto 0);
signal w_en2 : std_logic;

begin

  weigth_encoder1 : process (clk,rst)
  begin
    if rst = '1' then
        w_en2 <= '0';
        w_a2  <= 0; 
        w_d2  <= (others => '0');
    elsif rising_edge(clk) then
      if w_en = '1' then
        w_en2 <= w_en;
        w_a2  <= conv_integer(w_a); 
        w_d2  <= w_d;
      end if;
    end if;
  end process weigth_encoder1;

  weigth_encoder2 : process (clk)
  begin
    if rising_edge(clk) then
      if w_en2 = '1' then
        if w_a2 =   1 then w001 <= w_d2; end if;
        if w_a2 =   2 then w002 <= w_d2; end if;
        if w_a2 =   3 then w003 <= w_d2; end if;
        if w_a2 =   4 then w004 <= w_d2; end if;
        if w_a2 =   5 then w005 <= w_d2; end if;
        if w_a2 =   6 then w006 <= w_d2; end if;
        if w_a2 =   7 then w007 <= w_d2; end if;
        if w_a2 =   8 then w008 <= w_d2; end if;
        if w_a2 =   9 then w009 <= w_d2; end if;
        if w_a2 =  11 then w011 <= w_d2; end if;
        if w_a2 =  12 then w012 <= w_d2; end if;
        if w_a2 =  13 then w013 <= w_d2; end if;
        if w_a2 =  14 then w014 <= w_d2; end if;
        if w_a2 =  15 then w015 <= w_d2; end if;
        if w_a2 =  16 then w016 <= w_d2; end if;
        if w_a2 =  17 then w017 <= w_d2; end if;
        if w_a2 =  18 then w018 <= w_d2; end if;
        if w_a2 =  19 then w019 <= w_d2; end if;
        if w_a2 =  21 then w021 <= w_d2; end if;
        if w_a2 =  22 then w022 <= w_d2; end if;
        if w_a2 =  23 then w023 <= w_d2; end if;
        if w_a2 =  24 then w024 <= w_d2; end if;
        if w_a2 =  25 then w025 <= w_d2; end if;
        if w_a2 =  26 then w026 <= w_d2; end if;
        if w_a2 =  27 then w027 <= w_d2; end if;
        if w_a2 =  28 then w028 <= w_d2; end if;
        if w_a2 =  29 then w029 <= w_d2; end if;
        if w_a2 =  31 then w031 <= w_d2; end if;
        if w_a2 =  32 then w032 <= w_d2; end if;
        if w_a2 =  33 then w033 <= w_d2; end if;
        if w_a2 =  34 then w034 <= w_d2; end if;
        if w_a2 =  35 then w035 <= w_d2; end if;
        if w_a2 =  36 then w036 <= w_d2; end if;
        if w_a2 =  37 then w037 <= w_d2; end if;
        if w_a2 =  38 then w038 <= w_d2; end if;
        if w_a2 =  39 then w039 <= w_d2; end if;
        if w_a2 =  41 then w041 <= w_d2; end if;
        if w_a2 =  42 then w042 <= w_d2; end if;
        if w_a2 =  43 then w043 <= w_d2; end if;
        if w_a2 =  44 then w044 <= w_d2; end if;
        if w_a2 =  45 then w045 <= w_d2; end if;
        if w_a2 =  46 then w046 <= w_d2; end if;
        if w_a2 =  47 then w047 <= w_d2; end if;
        if w_a2 =  48 then w048 <= w_d2; end if;
        if w_a2 =  49 then w049 <= w_d2; end if;
        if w_a2 =  51 then w051 <= w_d2; end if;
        if w_a2 =  52 then w052 <= w_d2; end if; 
        if w_a2 =  53 then w053 <= w_d2; end if;
        if w_a2 =  54 then w054 <= w_d2; end if;
        if w_a2 =  55 then w055 <= w_d2; end if;
        if w_a2 =  56 then w056 <= w_d2; end if;
        if w_a2 =  57 then w057 <= w_d2; end if;
        if w_a2 =  58 then w058 <= w_d2; end if;
        if w_a2 =  59 then w059 <= w_d2; end if;
        if w_a2 =  61 then w061 <= w_d2; end if;
        if w_a2 =  62 then w062 <= w_d2; end if;
        if w_a2 =  63 then w063 <= w_d2; end if;
        if w_a2 =  64 then w064 <= w_d2; end if;
        if w_a2 =  65 then w065 <= w_d2; end if;
        if w_a2 =  66 then w066 <= w_d2; end if;
        if w_a2 =  67 then w067 <= w_d2; end if;
        if w_a2 =  68 then w068 <= w_d2; end if;
        if w_a2 =  69 then w069 <= w_d2; end if;
        if w_a2 =  71 then w071 <= w_d2; end if;
        if w_a2 =  72 then w072 <= w_d2; end if;
        if w_a2 =  73 then w073 <= w_d2; end if;
        if w_a2 =  74 then w074 <= w_d2; end if;
        if w_a2 =  75 then w075 <= w_d2; end if;
        if w_a2 =  76 then w076 <= w_d2; end if;
        if w_a2 =  77 then w077 <= w_d2; end if;
        if w_a2 =  78 then w078 <= w_d2; end if;
        if w_a2 =  79 then w079 <= w_d2; end if;
        if w_a2 =  81 then w081 <= w_d2; end if;
        if w_a2 =  82 then w082 <= w_d2; end if;
        if w_a2 =  83 then w083 <= w_d2; end if;
        if w_a2 =  84 then w084 <= w_d2; end if;
        if w_a2 =  85 then w085 <= w_d2; end if;
        if w_a2 =  86 then w086 <= w_d2; end if;
        if w_a2 =  87 then w087 <= w_d2; end if;
        if w_a2 =  88 then w088 <= w_d2; end if;
        if w_a2 =  89 then w089 <= w_d2; end if;
        if w_a2 =  91 then w091 <= w_d2; end if;
        if w_a2 =  92 then w092 <= w_d2; end if;
        if w_a2 =  93 then w093 <= w_d2; end if;
        if w_a2 =  94 then w094 <= w_d2; end if;
        if w_a2 =  95 then w095 <= w_d2; end if;
        if w_a2 =  96 then w096 <= w_d2; end if;
        if w_a2 =  97 then w097 <= w_d2; end if;
        if w_a2 =  98 then w098 <= w_d2; end if;
        if w_a2 =  99 then w099 <= w_d2; end if;
        if w_a2 = 101 then w101 <= w_d2; end if;
        if w_a2 = 102 then w102 <= w_d2; end if;
        if w_a2 = 103 then w103 <= w_d2; end if;
        if w_a2 = 104 then w104 <= w_d2; end if;
        if w_a2 = 105 then w105 <= w_d2; end if;
        if w_a2 = 106 then w106 <= w_d2; end if;
        if w_a2 = 107 then w107 <= w_d2; end if;
        if w_a2 = 108 then w108 <= w_d2; end if;
        if w_a2 = 109 then w109 <= w_d2; end if;
        if w_a2 = 111 then w111 <= w_d2; end if;
        if w_a2 = 112 then w112 <= w_d2; end if;
        if w_a2 = 113 then w113 <= w_d2; end if;
        if w_a2 = 114 then w114 <= w_d2; end if;
        if w_a2 = 115 then w115 <= w_d2; end if;
        if w_a2 = 116 then w116 <= w_d2; end if;
        if w_a2 = 117 then w117 <= w_d2; end if;
        if w_a2 = 118 then w118 <= w_d2; end if;
        if w_a2 = 119 then w119 <= w_d2; end if;
        if w_a2 = 121 then w121 <= w_d2; end if;
        if w_a2 = 122 then w122 <= w_d2; end if;
        if w_a2 = 123 then w123 <= w_d2; end if;
        if w_a2 = 124 then w124 <= w_d2; end if;
        if w_a2 = 125 then w125 <= w_d2; end if;
        if w_a2 = 126 then w126 <= w_d2; end if;
        if w_a2 = 127 then w127 <= w_d2; end if;
        if w_a2 = 128 then w128 <= w_d2; end if;
        if w_a2 = 129 then w129 <= w_d2; end if;
        if w_a2 = 131 then w131 <= w_d2; end if;
        if w_a2 = 132 then w132 <= w_d2; end if;
        if w_a2 = 133 then w133 <= w_d2; end if;
        if w_a2 = 134 then w134 <= w_d2; end if;
        if w_a2 = 135 then w135 <= w_d2; end if;
        if w_a2 = 136 then w136 <= w_d2; end if;
        if w_a2 = 137 then w137 <= w_d2; end if;
        if w_a2 = 138 then w138 <= w_d2; end if;
        if w_a2 = 139 then w139 <= w_d2; end if;
        if w_a2 = 141 then w141 <= w_d2; end if;
        if w_a2 = 142 then w142 <= w_d2; end if;
        if w_a2 = 143 then w143 <= w_d2; end if;
        if w_a2 = 144 then w144 <= w_d2; end if;
        if w_a2 = 145 then w145 <= w_d2; end if;
        if w_a2 = 146 then w146 <= w_d2; end if;
        if w_a2 = 147 then w147 <= w_d2; end if;
        if w_a2 = 148 then w148 <= w_d2; end if;
        if w_a2 = 149 then w149 <= w_d2; end if;
        if w_a2 = 151 then w151 <= w_d2; end if;
        if w_a2 = 152 then w152 <= w_d2; end if;
        if w_a2 = 153 then w153 <= w_d2; end if;
        if w_a2 = 154 then w154 <= w_d2; end if;
        if w_a2 = 155 then w155 <= w_d2; end if;
        if w_a2 = 156 then w156 <= w_d2; end if;
        if w_a2 = 157 then w157 <= w_d2; end if;
        if w_a2 = 158 then w158 <= w_d2; end if;
        if w_a2 = 159 then w159 <= w_d2; end if;
        if w_a2 = 161 then w161 <= w_d2; end if;
        if w_a2 = 162 then w162 <= w_d2; end if;
        if w_a2 = 163 then w163 <= w_d2; end if;
        if w_a2 = 164 then w164 <= w_d2; end if;
        if w_a2 = 165 then w165 <= w_d2; end if;
        if w_a2 = 166 then w166 <= w_d2; end if;
        if w_a2 = 167 then w167 <= w_d2; end if;
        if w_a2 = 168 then w168 <= w_d2; end if;
        if w_a2 = 169 then w169 <= w_d2; end if;
        if w_a2 = 171 then w171 <= w_d2; end if;
        if w_a2 = 172 then w172 <= w_d2; end if;
        if w_a2 = 173 then w173 <= w_d2; end if;
        if w_a2 = 174 then w174 <= w_d2; end if;
        if w_a2 = 175 then w175 <= w_d2; end if;
        if w_a2 = 176 then w176 <= w_d2; end if;
        if w_a2 = 177 then w177 <= w_d2; end if;
        if w_a2 = 178 then w178 <= w_d2; end if;
        if w_a2 = 179 then w179 <= w_d2; end if;
        if w_a2 = 181 then w181 <= w_d2; end if;
        if w_a2 = 182 then w182 <= w_d2; end if;
        if w_a2 = 183 then w183 <= w_d2; end if;
        if w_a2 = 184 then w184 <= w_d2; end if;
        if w_a2 = 185 then w185 <= w_d2; end if;
        if w_a2 = 186 then w186 <= w_d2; end if;
        if w_a2 = 187 then w187 <= w_d2; end if;
        if w_a2 = 188 then w188 <= w_d2; end if;
        if w_a2 = 189 then w189 <= w_d2; end if;
        if w_a2 = 191 then w191 <= w_d2; end if;
        if w_a2 = 192 then w192 <= w_d2; end if;
        if w_a2 = 193 then w193 <= w_d2; end if;
        if w_a2 = 194 then w194 <= w_d2; end if;
        if w_a2 = 195 then w195 <= w_d2; end if;
        if w_a2 = 196 then w196 <= w_d2; end if;
        if w_a2 = 197 then w197 <= w_d2; end if;
        if w_a2 = 198 then w198 <= w_d2; end if;
        if w_a2 = 199 then w199 <= w_d2; end if;
        if w_a2 = 201 then w201 <= w_d2; end if;
        if w_a2 = 202 then w202 <= w_d2; end if;
        if w_a2 = 203 then w203 <= w_d2; end if;
        if w_a2 = 204 then w204 <= w_d2; end if;
        if w_a2 = 205 then w205 <= w_d2; end if;
        if w_a2 = 206 then w206 <= w_d2; end if;
        if w_a2 = 207 then w207 <= w_d2; end if;
        if w_a2 = 208 then w208 <= w_d2; end if;
        if w_a2 = 209 then w209 <= w_d2; end if;
        if w_a2 = 211 then w211 <= w_d2; end if;
        if w_a2 = 212 then w212 <= w_d2; end if;
        if w_a2 = 213 then w213 <= w_d2; end if;
        if w_a2 = 214 then w214 <= w_d2; end if;
        if w_a2 = 215 then w215 <= w_d2; end if;
        if w_a2 = 216 then w216 <= w_d2; end if;
        if w_a2 = 217 then w217 <= w_d2; end if;
        if w_a2 = 218 then w218 <= w_d2; end if;
        if w_a2 = 219 then w219 <= w_d2; end if;
        if w_a2 = 221 then w221 <= w_d2; end if;
        if w_a2 = 222 then w222 <= w_d2; end if;
        if w_a2 = 223 then w223 <= w_d2; end if;
        if w_a2 = 224 then w224 <= w_d2; end if;
        if w_a2 = 225 then w225 <= w_d2; end if;
        if w_a2 = 226 then w226 <= w_d2; end if;
        if w_a2 = 227 then w227 <= w_d2; end if;
        if w_a2 = 228 then w228 <= w_d2; end if;
        if w_a2 = 229 then w229 <= w_d2; end if;
        if w_a2 = 231 then w231 <= w_d2; end if;
        if w_a2 = 232 then w232 <= w_d2; end if;
        if w_a2 = 233 then w233 <= w_d2; end if;
        if w_a2 = 234 then w234 <= w_d2; end if;
        if w_a2 = 235 then w235 <= w_d2; end if;
        if w_a2 = 236 then w236 <= w_d2; end if;
        if w_a2 = 237 then w237 <= w_d2; end if;
        if w_a2 = 238 then w238 <= w_d2; end if;
        if w_a2 = 239 then w239 <= w_d2; end if;
        if w_a2 = 241 then w241 <= w_d2; end if;
        if w_a2 = 242 then w242 <= w_d2; end if;
        if w_a2 = 243 then w243 <= w_d2; end if;
        if w_a2 = 244 then w244 <= w_d2; end if;
        if w_a2 = 245 then w245 <= w_d2; end if;
        if w_a2 = 246 then w246 <= w_d2; end if;
        if w_a2 = 247 then w247 <= w_d2; end if;
        if w_a2 = 248 then w248 <= w_d2; end if;
        if w_a2 = 249 then w249 <= w_d2; end if;
        if w_a2 = 251 then w251 <= w_d2; end if;
        if w_a2 = 252 then w252 <= w_d2; end if;
        if w_a2 = 253 then w253 <= w_d2; end if;
        if w_a2 = 254 then w254 <= w_d2; end if;
        if w_a2 = 255 then w255 <= w_d2; end if;
        if w_a2 = 256 then w256 <= w_d2; end if;
        if w_a2 = 257 then w257 <= w_d2; end if;
        if w_a2 = 258 then w258 <= w_d2; end if;
        if w_a2 = 259 then w259 <= w_d2; end if;
        if w_a2 = 261 then w261 <= w_d2; end if;
        if w_a2 = 262 then w262 <= w_d2; end if;
        if w_a2 = 263 then w263 <= w_d2; end if;
        if w_a2 = 264 then w264 <= w_d2; end if;
        if w_a2 = 265 then w265 <= w_d2; end if;
        if w_a2 = 266 then w266 <= w_d2; end if;
        if w_a2 = 267 then w267 <= w_d2; end if;
        if w_a2 = 268 then w268 <= w_d2; end if;
        if w_a2 = 269 then w269 <= w_d2; end if;
        if w_a2 = 271 then w271 <= w_d2; end if;
        if w_a2 = 272 then w272 <= w_d2; end if;
        if w_a2 = 273 then w273 <= w_d2; end if;
        if w_a2 = 274 then w274 <= w_d2; end if;
        if w_a2 = 275 then w275 <= w_d2; end if;
        if w_a2 = 276 then w276 <= w_d2; end if;
        if w_a2 = 277 then w277 <= w_d2; end if;
        if w_a2 = 278 then w278 <= w_d2; end if;
        if w_a2 = 279 then w279 <= w_d2; end if;
        if w_a2 = 281 then w281 <= w_d2; end if;
        if w_a2 = 282 then w282 <= w_d2; end if;
        if w_a2 = 283 then w283 <= w_d2; end if;
        if w_a2 = 284 then w284 <= w_d2; end if;
        if w_a2 = 285 then w285 <= w_d2; end if;
        if w_a2 = 286 then w286 <= w_d2; end if;
        if w_a2 = 287 then w287 <= w_d2; end if;
        if w_a2 = 288 then w288 <= w_d2; end if;
        if w_a2 = 289 then w289 <= w_d2; end if;
        if w_a2 = 291 then w291 <= w_d2; end if;
        if w_a2 = 292 then w292 <= w_d2; end if;
        if w_a2 = 293 then w293 <= w_d2; end if;
        if w_a2 = 294 then w294 <= w_d2; end if;
        if w_a2 = 295 then w295 <= w_d2; end if;
        if w_a2 = 296 then w296 <= w_d2; end if;
        if w_a2 = 297 then w297 <= w_d2; end if;
        if w_a2 = 298 then w298 <= w_d2; end if;
        if w_a2 = 299 then w299 <= w_d2; end if;
        if w_a2 = 301 then w301 <= w_d2; end if;
        if w_a2 = 302 then w302 <= w_d2; end if;
        if w_a2 = 303 then w303 <= w_d2; end if;
        if w_a2 = 304 then w304 <= w_d2; end if;
        if w_a2 = 305 then w305 <= w_d2; end if;
        if w_a2 = 306 then w306 <= w_d2; end if;
        if w_a2 = 307 then w307 <= w_d2; end if;
        if w_a2 = 308 then w308 <= w_d2; end if;
        if w_a2 = 309 then w309 <= w_d2; end if;
        if w_a2 = 311 then w311 <= w_d2; end if;
        if w_a2 = 312 then w312 <= w_d2; end if;
        if w_a2 = 313 then w313 <= w_d2; end if;
        if w_a2 = 314 then w314 <= w_d2; end if;
        if w_a2 = 315 then w315 <= w_d2; end if;
        if w_a2 = 316 then w316 <= w_d2; end if;
        if w_a2 = 317 then w317 <= w_d2; end if;
        if w_a2 = 318 then w318 <= w_d2; end if;
        if w_a2 = 319 then w319 <= w_d2; end if;
        if w_a2 = 321 then w321 <= w_d2; end if;
        if w_a2 = 322 then w322 <= w_d2; end if;
        if w_a2 = 323 then w323 <= w_d2; end if;
        if w_a2 = 324 then w324 <= w_d2; end if;
        if w_a2 = 325 then w325 <= w_d2; end if;
        if w_a2 = 326 then w326 <= w_d2; end if;
        if w_a2 = 327 then w327 <= w_d2; end if;
        if w_a2 = 328 then w328 <= w_d2; end if;
        if w_a2 = 329 then w329 <= w_d2; end if;
        if w_a2 = 331 then w331 <= w_d2; end if;
        if w_a2 = 332 then w332 <= w_d2; end if;
        if w_a2 = 333 then w333 <= w_d2; end if;
        if w_a2 = 334 then w334 <= w_d2; end if;
        if w_a2 = 335 then w335 <= w_d2; end if;
        if w_a2 = 336 then w336 <= w_d2; end if;
        if w_a2 = 337 then w337 <= w_d2; end if;
        if w_a2 = 338 then w338 <= w_d2; end if;
        if w_a2 = 339 then w339 <= w_d2; end if;
        if w_a2 = 341 then w341 <= w_d2; end if;
        if w_a2 = 342 then w342 <= w_d2; end if;
        if w_a2 = 343 then w343 <= w_d2; end if;
        if w_a2 = 344 then w344 <= w_d2; end if;
        if w_a2 = 345 then w345 <= w_d2; end if;
        if w_a2 = 346 then w346 <= w_d2; end if;
        if w_a2 = 347 then w347 <= w_d2; end if;
        if w_a2 = 348 then w348 <= w_d2; end if;
        if w_a2 = 349 then w349 <= w_d2; end if;
        if w_a2 = 351 then w351 <= w_d2; end if;
        if w_a2 = 352 then w352 <= w_d2; end if;
        if w_a2 = 353 then w353 <= w_d2; end if;
        if w_a2 = 354 then w354 <= w_d2; end if;
        if w_a2 = 355 then w355 <= w_d2; end if;
        if w_a2 = 356 then w356 <= w_d2; end if;
        if w_a2 = 357 then w357 <= w_d2; end if;
        if w_a2 = 358 then w358 <= w_d2; end if;
        if w_a2 = 359 then w359 <= w_d2; end if;
        if w_a2 = 361 then w361 <= w_d2; end if;
        if w_a2 = 362 then w362 <= w_d2; end if;
        if w_a2 = 363 then w363 <= w_d2; end if;
        if w_a2 = 364 then w364 <= w_d2; end if;
        if w_a2 = 365 then w365 <= w_d2; end if;
        if w_a2 = 366 then w366 <= w_d2; end if;
        if w_a2 = 367 then w367 <= w_d2; end if;
        if w_a2 = 368 then w368 <= w_d2; end if;
        if w_a2 = 369 then w369 <= w_d2; end if;
        if w_a2 = 371 then w371 <= w_d2; end if;
        if w_a2 = 372 then w372 <= w_d2; end if;
        if w_a2 = 373 then w373 <= w_d2; end if;
        if w_a2 = 374 then w374 <= w_d2; end if;
        if w_a2 = 375 then w375 <= w_d2; end if;
        if w_a2 = 376 then w376 <= w_d2; end if;
        if w_a2 = 377 then w377 <= w_d2; end if;
        if w_a2 = 378 then w378 <= w_d2; end if;
        if w_a2 = 379 then w379 <= w_d2; end if;
        if w_a2 = 381 then w381 <= w_d2; end if;
        if w_a2 = 382 then w382 <= w_d2; end if;
        if w_a2 = 383 then w383 <= w_d2; end if;
        if w_a2 = 384 then w384 <= w_d2; end if;
        if w_a2 = 385 then w385 <= w_d2; end if;
        if w_a2 = 386 then w386 <= w_d2; end if;
        if w_a2 = 387 then w387 <= w_d2; end if;
        if w_a2 = 388 then w388 <= w_d2; end if;
        if w_a2 = 389 then w389 <= w_d2; end if;
        if w_a2 = 391 then w391 <= w_d2; end if;
        if w_a2 = 392 then w392 <= w_d2; end if;
        if w_a2 = 393 then w393 <= w_d2; end if;
        if w_a2 = 394 then w394 <= w_d2; end if;
        if w_a2 = 395 then w395 <= w_d2; end if;
        if w_a2 = 396 then w396 <= w_d2; end if;
        if w_a2 = 397 then w397 <= w_d2; end if;
        if w_a2 = 398 then w398 <= w_d2; end if;
        if w_a2 = 399 then w399 <= w_d2; end if;
        if w_a2 = 401 then w401 <= w_d2; end if;
        if w_a2 = 402 then w402 <= w_d2; end if;
        if w_a2 = 403 then w403 <= w_d2; end if;
        if w_a2 = 404 then w404 <= w_d2; end if;
        if w_a2 = 405 then w405 <= w_d2; end if;
        if w_a2 = 406 then w406 <= w_d2; end if;
        if w_a2 = 407 then w407 <= w_d2; end if;
        if w_a2 = 408 then w408 <= w_d2; end if;
        if w_a2 = 409 then w409 <= w_d2; end if;
        if w_a2 = 411 then w411 <= w_d2; end if;
        if w_a2 = 412 then w412 <= w_d2; end if;
        if w_a2 = 413 then w413 <= w_d2; end if;
        if w_a2 = 414 then w414 <= w_d2; end if;
        if w_a2 = 415 then w415 <= w_d2; end if;
        if w_a2 = 416 then w416 <= w_d2; end if;
        if w_a2 = 417 then w417 <= w_d2; end if;
        if w_a2 = 418 then w418 <= w_d2; end if;
        if w_a2 = 419 then w419 <= w_d2; end if;
        if w_a2 = 421 then w421 <= w_d2; end if;
        if w_a2 = 422 then w422 <= w_d2; end if;
        if w_a2 = 423 then w423 <= w_d2; end if;
        if w_a2 = 424 then w424 <= w_d2; end if;
        if w_a2 = 425 then w425 <= w_d2; end if;
        if w_a2 = 426 then w426 <= w_d2; end if;
        if w_a2 = 427 then w427 <= w_d2; end if;
        if w_a2 = 428 then w428 <= w_d2; end if;
        if w_a2 = 429 then w429 <= w_d2; end if;
        if w_a2 = 431 then w431 <= w_d2; end if;
        if w_a2 = 432 then w432 <= w_d2; end if;
        if w_a2 = 433 then w433 <= w_d2; end if;
        if w_a2 = 434 then w434 <= w_d2; end if;
        if w_a2 = 435 then w435 <= w_d2; end if;
        if w_a2 = 436 then w436 <= w_d2; end if;
        if w_a2 = 437 then w437 <= w_d2; end if;
        if w_a2 = 438 then w438 <= w_d2; end if;
        if w_a2 = 439 then w439 <= w_d2; end if;
        if w_a2 = 441 then w441 <= w_d2; end if;
        if w_a2 = 442 then w442 <= w_d2; end if;
        if w_a2 = 443 then w443 <= w_d2; end if;
        if w_a2 = 444 then w444 <= w_d2; end if;
        if w_a2 = 445 then w445 <= w_d2; end if;
        if w_a2 = 446 then w446 <= w_d2; end if;
        if w_a2 = 447 then w447 <= w_d2; end if;
        if w_a2 = 448 then w448 <= w_d2; end if;
        if w_a2 = 449 then w449 <= w_d2; end if;
        if w_a2 = 451 then w451 <= w_d2; end if;
        if w_a2 = 452 then w452 <= w_d2; end if;
        if w_a2 = 453 then w453 <= w_d2; end if;
        if w_a2 = 454 then w454 <= w_d2; end if;
        if w_a2 = 455 then w455 <= w_d2; end if;
        if w_a2 = 456 then w456 <= w_d2; end if;
        if w_a2 = 457 then w457 <= w_d2; end if;
        if w_a2 = 458 then w458 <= w_d2; end if;
        if w_a2 = 459 then w459 <= w_d2; end if;
        if w_a2 = 461 then w461 <= w_d2; end if;
        if w_a2 = 462 then w462 <= w_d2; end if;
        if w_a2 = 463 then w463 <= w_d2; end if;
        if w_a2 = 464 then w464 <= w_d2; end if;
        if w_a2 = 465 then w465 <= w_d2; end if;
        if w_a2 = 466 then w466 <= w_d2; end if;
        if w_a2 = 467 then w467 <= w_d2; end if;
        if w_a2 = 468 then w468 <= w_d2; end if;
        if w_a2 = 469 then w469 <= w_d2; end if;
        if w_a2 = 471 then w471 <= w_d2; end if;
        if w_a2 = 472 then w472 <= w_d2; end if;
        if w_a2 = 473 then w473 <= w_d2; end if;
        if w_a2 = 474 then w474 <= w_d2; end if;
        if w_a2 = 475 then w475 <= w_d2; end if;
        if w_a2 = 476 then w476 <= w_d2; end if;
        if w_a2 = 477 then w477 <= w_d2; end if;
        if w_a2 = 478 then w478 <= w_d2; end if;
        if w_a2 = 479 then w479 <= w_d2; end if;
        if w_a2 = 481 then w481 <= w_d2; end if;
        if w_a2 = 482 then w482 <= w_d2; end if;
        if w_a2 = 483 then w483 <= w_d2; end if;
        if w_a2 = 484 then w484 <= w_d2; end if;
        if w_a2 = 485 then w485 <= w_d2; end if;
        if w_a2 = 486 then w486 <= w_d2; end if;
        if w_a2 = 487 then w487 <= w_d2; end if;
        if w_a2 = 488 then w488 <= w_d2; end if;
        if w_a2 = 489 then w489 <= w_d2; end if;
        if w_a2 = 491 then w491 <= w_d2; end if;
        if w_a2 = 492 then w492 <= w_d2; end if;
        if w_a2 = 493 then w493 <= w_d2; end if;
        if w_a2 = 494 then w494 <= w_d2; end if;
        if w_a2 = 495 then w495 <= w_d2; end if;
        if w_a2 = 496 then w496 <= w_d2; end if;
        if w_a2 = 497 then w497 <= w_d2; end if;
        if w_a2 = 498 then w498 <= w_d2; end if;
        if w_a2 = 499 then w499 <= w_d2; end if;
        if w_a2 = 501 then w501 <= w_d2; end if;
        if w_a2 = 502 then w502 <= w_d2; end if;
        if w_a2 = 503 then w503 <= w_d2; end if;
        if w_a2 = 504 then w504 <= w_d2; end if;
        if w_a2 = 505 then w505 <= w_d2; end if;
        if w_a2 = 506 then w506 <= w_d2; end if;
        if w_a2 = 507 then w507 <= w_d2; end if;
        if w_a2 = 508 then w508 <= w_d2; end if;
        if w_a2 = 509 then w509 <= w_d2; end if;
        if w_a2 = 511 then w511 <= w_d2; end if;
        if w_a2 = 512 then w512 <= w_d2; end if;
        if w_a2 = 513 then w513 <= w_d2; end if;
        if w_a2 = 514 then w514 <= w_d2; end if;
        if w_a2 = 515 then w515 <= w_d2; end if;
        if w_a2 = 516 then w516 <= w_d2; end if;
        if w_a2 = 517 then w517 <= w_d2; end if;
        if w_a2 = 518 then w518 <= w_d2; end if;
        if w_a2 = 519 then w519 <= w_d2; end if;
        if w_a2 = 521 then w521 <= w_d2; end if;
        if w_a2 = 522 then w522 <= w_d2; end if;
        if w_a2 = 523 then w523 <= w_d2; end if;
        if w_a2 = 524 then w524 <= w_d2; end if;
        if w_a2 = 525 then w525 <= w_d2; end if;
        if w_a2 = 526 then w526 <= w_d2; end if;
        if w_a2 = 527 then w527 <= w_d2; end if;
        if w_a2 = 528 then w528 <= w_d2; end if;
        if w_a2 = 529 then w529 <= w_d2; end if;
        if w_a2 = 531 then w531 <= w_d2; end if;
        if w_a2 = 532 then w532 <= w_d2; end if;
        if w_a2 = 533 then w533 <= w_d2; end if;
        if w_a2 = 534 then w534 <= w_d2; end if;
        if w_a2 = 535 then w535 <= w_d2; end if;
        if w_a2 = 536 then w536 <= w_d2; end if;
        if w_a2 = 537 then w537 <= w_d2; end if;
        if w_a2 = 538 then w538 <= w_d2; end if;
        if w_a2 = 539 then w539 <= w_d2; end if;
        if w_a2 = 541 then w541 <= w_d2; end if;
        if w_a2 = 542 then w542 <= w_d2; end if;
        if w_a2 = 543 then w543 <= w_d2; end if;
        if w_a2 = 544 then w544 <= w_d2; end if;
        if w_a2 = 545 then w545 <= w_d2; end if;
        if w_a2 = 546 then w546 <= w_d2; end if;
        if w_a2 = 547 then w547 <= w_d2; end if;
        if w_a2 = 548 then w548 <= w_d2; end if;
        if w_a2 = 549 then w549 <= w_d2; end if;
        if w_a2 = 551 then w551 <= w_d2; end if;
        if w_a2 = 552 then w552 <= w_d2; end if;
        if w_a2 = 553 then w553 <= w_d2; end if;
        if w_a2 = 554 then w554 <= w_d2; end if;
        if w_a2 = 555 then w555 <= w_d2; end if;
        if w_a2 = 556 then w556 <= w_d2; end if;
        if w_a2 = 557 then w557 <= w_d2; end if;
        if w_a2 = 558 then w558 <= w_d2; end if;
        if w_a2 = 559 then w559 <= w_d2; end if;
        if w_a2 = 561 then w561 <= w_d2; end if;
        if w_a2 = 562 then w562 <= w_d2; end if;
        if w_a2 = 563 then w563 <= w_d2; end if;
        if w_a2 = 564 then w564 <= w_d2; end if;
        if w_a2 = 565 then w565 <= w_d2; end if;
        if w_a2 = 566 then w566 <= w_d2; end if;
        if w_a2 = 567 then w567 <= w_d2; end if;
        if w_a2 = 568 then w568 <= w_d2; end if;
        if w_a2 = 569 then w569 <= w_d2; end if;
        if w_a2 = 571 then w571 <= w_d2; end if;
        if w_a2 = 572 then w572 <= w_d2; end if;
        if w_a2 = 573 then w573 <= w_d2; end if;
        if w_a2 = 574 then w574 <= w_d2; end if;
        if w_a2 = 575 then w575 <= w_d2; end if;
        if w_a2 = 576 then w576 <= w_d2; end if;
        if w_a2 = 577 then w577 <= w_d2; end if;
        if w_a2 = 578 then w578 <= w_d2; end if;
        if w_a2 = 579 then w579 <= w_d2; end if;
        if w_a2 = 581 then w581 <= w_d2; end if;
        if w_a2 = 582 then w582 <= w_d2; end if;
        if w_a2 = 583 then w583 <= w_d2; end if;
        if w_a2 = 584 then w584 <= w_d2; end if;
        if w_a2 = 585 then w585 <= w_d2; end if;
        if w_a2 = 586 then w586 <= w_d2; end if;
        if w_a2 = 587 then w587 <= w_d2; end if;
        if w_a2 = 588 then w588 <= w_d2; end if;
        if w_a2 = 589 then w589 <= w_d2; end if;
        if w_a2 = 591 then w591 <= w_d2; end if;
        if w_a2 = 592 then w592 <= w_d2; end if;
        if w_a2 = 593 then w593 <= w_d2; end if;
        if w_a2 = 594 then w594 <= w_d2; end if;
        if w_a2 = 595 then w595 <= w_d2; end if;
        if w_a2 = 596 then w596 <= w_d2; end if;
        if w_a2 = 597 then w597 <= w_d2; end if;
        if w_a2 = 598 then w598 <= w_d2; end if;
        if w_a2 = 599 then w599 <= w_d2; end if;
        if w_a2 = 601 then w601 <= w_d2; end if;
        if w_a2 = 602 then w602 <= w_d2; end if;
        if w_a2 = 603 then w603 <= w_d2; end if;
        if w_a2 = 604 then w604 <= w_d2; end if;
        if w_a2 = 605 then w605 <= w_d2; end if;
        if w_a2 = 606 then w606 <= w_d2; end if;
        if w_a2 = 607 then w607 <= w_d2; end if;
        if w_a2 = 608 then w608 <= w_d2; end if;
        if w_a2 = 609 then w609 <= w_d2; end if;
        if w_a2 = 611 then w611 <= w_d2; end if;
        if w_a2 = 612 then w612 <= w_d2; end if;
        if w_a2 = 613 then w613 <= w_d2; end if;
        if w_a2 = 614 then w614 <= w_d2; end if;
        if w_a2 = 615 then w615 <= w_d2; end if;
        if w_a2 = 616 then w616 <= w_d2; end if;
        if w_a2 = 617 then w617 <= w_d2; end if;
        if w_a2 = 618 then w618 <= w_d2; end if;
        if w_a2 = 619 then w619 <= w_d2; end if;
        if w_a2 = 621 then w621 <= w_d2; end if;
        if w_a2 = 622 then w622 <= w_d2; end if;
        if w_a2 = 623 then w623 <= w_d2; end if;
        if w_a2 = 624 then w624 <= w_d2; end if;
        if w_a2 = 625 then w625 <= w_d2; end if;
        if w_a2 = 626 then w626 <= w_d2; end if;
        if w_a2 = 627 then w627 <= w_d2; end if;
        if w_a2 = 628 then w628 <= w_d2; end if;
        if w_a2 = 629 then w629 <= w_d2; end if;
        if w_a2 = 631 then w631 <= w_d2; end if;
        if w_a2 = 632 then w632 <= w_d2; end if;
        if w_a2 = 633 then w633 <= w_d2; end if;
        if w_a2 = 634 then w634 <= w_d2; end if;
        if w_a2 = 635 then w635 <= w_d2; end if;
        if w_a2 = 636 then w636 <= w_d2; end if;
        if w_a2 = 637 then w637 <= w_d2; end if;
        if w_a2 = 638 then w638 <= w_d2; end if;
        if w_a2 = 639 then w639 <= w_d2; end if;
        if w_a2 = 641 then w641 <= w_d2; end if;
        if w_a2 = 642 then w642 <= w_d2; end if;
        if w_a2 = 643 then w643 <= w_d2; end if;
        if w_a2 = 644 then w644 <= w_d2; end if;
        if w_a2 = 645 then w645 <= w_d2; end if;
        if w_a2 = 646 then w646 <= w_d2; end if;
        if w_a2 = 647 then w647 <= w_d2; end if;
        if w_a2 = 648 then w648 <= w_d2; end if;
        if w_a2 = 649 then w649 <= w_d2; end if;
        if w_a2 = 651 then w651 <= w_d2; end if;
        if w_a2 = 652 then w652 <= w_d2; end if;
        if w_a2 = 653 then w653 <= w_d2; end if;
        if w_a2 = 654 then w654 <= w_d2; end if;
        if w_a2 = 655 then w655 <= w_d2; end if;
        if w_a2 = 656 then w656 <= w_d2; end if;
        if w_a2 = 657 then w657 <= w_d2; end if;
        if w_a2 = 658 then w658 <= w_d2; end if;
        if w_a2 = 659 then w659 <= w_d2; end if;
        if w_a2 = 661 then w661 <= w_d2; end if;
        if w_a2 = 662 then w662 <= w_d2; end if;
        if w_a2 = 663 then w663 <= w_d2; end if;
        if w_a2 = 664 then w664 <= w_d2; end if;
        if w_a2 = 665 then w665 <= w_d2; end if;
        if w_a2 = 666 then w666 <= w_d2; end if;
        if w_a2 = 667 then w667 <= w_d2; end if;
        if w_a2 = 668 then w668 <= w_d2; end if;
        if w_a2 = 669 then w669 <= w_d2; end if;
        if w_a2 = 671 then w671 <= w_d2; end if;
        if w_a2 = 672 then w672 <= w_d2; end if;
        if w_a2 = 673 then w673 <= w_d2; end if;
        if w_a2 = 674 then w674 <= w_d2; end if;
        if w_a2 = 675 then w675 <= w_d2; end if;
        if w_a2 = 676 then w676 <= w_d2; end if;
        if w_a2 = 677 then w677 <= w_d2; end if;
        if w_a2 = 678 then w678 <= w_d2; end if;
        if w_a2 = 679 then w679 <= w_d2; end if;
        if w_a2 = 681 then w681 <= w_d2; end if;
        if w_a2 = 682 then w682 <= w_d2; end if;
        if w_a2 = 683 then w683 <= w_d2; end if;
        if w_a2 = 684 then w684 <= w_d2; end if;
        if w_a2 = 685 then w685 <= w_d2; end if;
        if w_a2 = 686 then w686 <= w_d2; end if;
        if w_a2 = 687 then w687 <= w_d2; end if;
        if w_a2 = 688 then w688 <= w_d2; end if;
        if w_a2 = 689 then w689 <= w_d2; end if;
        if w_a2 = 691 then w691 <= w_d2; end if;
        if w_a2 = 692 then w692 <= w_d2; end if;
        if w_a2 = 693 then w693 <= w_d2; end if;
        if w_a2 = 694 then w694 <= w_d2; end if;
        if w_a2 = 695 then w695 <= w_d2; end if;
        if w_a2 = 696 then w696 <= w_d2; end if;
        if w_a2 = 697 then w697 <= w_d2; end if;
        if w_a2 = 698 then w698 <= w_d2; end if;
        if w_a2 = 699 then w699 <= w_d2; end if;
        if w_a2 = 701 then w701 <= w_d2; end if;
        if w_a2 = 702 then w702 <= w_d2; end if;
        if w_a2 = 703 then w703 <= w_d2; end if;
        if w_a2 = 704 then w704 <= w_d2; end if;
        if w_a2 = 705 then w705 <= w_d2; end if;
        if w_a2 = 706 then w706 <= w_d2; end if;
        if w_a2 = 707 then w707 <= w_d2; end if;
        if w_a2 = 708 then w708 <= w_d2; end if;
        if w_a2 = 709 then w709 <= w_d2; end if;
        if w_a2 = 711 then w711 <= w_d2; end if;
        if w_a2 = 712 then w712 <= w_d2; end if;
        if w_a2 = 713 then w713 <= w_d2; end if;
        if w_a2 = 714 then w714 <= w_d2; end if;
        if w_a2 = 715 then w715 <= w_d2; end if;
        if w_a2 = 716 then w716 <= w_d2; end if;
        if w_a2 = 717 then w717 <= w_d2; end if;
        if w_a2 = 718 then w718 <= w_d2; end if;
        if w_a2 = 719 then w719 <= w_d2; end if;
        if w_a2 = 721 then w721 <= w_d2; end if;
        if w_a2 = 722 then w722 <= w_d2; end if;
        if w_a2 = 723 then w723 <= w_d2; end if;
        if w_a2 = 724 then w724 <= w_d2; end if;
        if w_a2 = 725 then w725 <= w_d2; end if;
        if w_a2 = 726 then w726 <= w_d2; end if;
        if w_a2 = 727 then w727 <= w_d2; end if;
        if w_a2 = 728 then w728 <= w_d2; end if;
        if w_a2 = 729 then w729 <= w_d2; end if;
        if w_a2 = 731 then w731 <= w_d2; end if;
        if w_a2 = 732 then w732 <= w_d2; end if;
        if w_a2 = 733 then w733 <= w_d2; end if;
        if w_a2 = 734 then w734 <= w_d2; end if;
        if w_a2 = 735 then w735 <= w_d2; end if;
        if w_a2 = 736 then w736 <= w_d2; end if;
        if w_a2 = 737 then w737 <= w_d2; end if;
        if w_a2 = 738 then w738 <= w_d2; end if;
        if w_a2 = 739 then w739 <= w_d2; end if;
        if w_a2 = 741 then w741 <= w_d2; end if;
        if w_a2 = 742 then w742 <= w_d2; end if;
        if w_a2 = 743 then w743 <= w_d2; end if;
        if w_a2 = 744 then w744 <= w_d2; end if;
        if w_a2 = 745 then w745 <= w_d2; end if;
        if w_a2 = 746 then w746 <= w_d2; end if;
        if w_a2 = 747 then w747 <= w_d2; end if;
        if w_a2 = 748 then w748 <= w_d2; end if;
        if w_a2 = 749 then w749 <= w_d2; end if;
        if w_a2 = 751 then w751 <= w_d2; end if;
        if w_a2 = 752 then w752 <= w_d2; end if;
        if w_a2 = 753 then w753 <= w_d2; end if;
        if w_a2 = 754 then w754 <= w_d2; end if;
        if w_a2 = 755 then w755 <= w_d2; end if;
        if w_a2 = 756 then w756 <= w_d2; end if;
        if w_a2 = 757 then w757 <= w_d2; end if;
        if w_a2 = 758 then w758 <= w_d2; end if;
        if w_a2 = 759 then w759 <= w_d2; end if;
        if w_a2 = 761 then w761 <= w_d2; end if;
        if w_a2 = 762 then w762 <= w_d2; end if;
        if w_a2 = 763 then w763 <= w_d2; end if;
        if w_a2 = 764 then w764 <= w_d2; end if;
        if w_a2 = 765 then w765 <= w_d2; end if;
        if w_a2 = 766 then w766 <= w_d2; end if;
        if w_a2 = 767 then w767 <= w_d2; end if;
        if w_a2 = 768 then w768 <= w_d2; end if;
        if w_a2 = 769 then w769 <= w_d2; end if;
        if w_a2 = 771 then w771 <= w_d2; end if;
        if w_a2 = 772 then w772 <= w_d2; end if;
        if w_a2 = 773 then w773 <= w_d2; end if;
        if w_a2 = 774 then w774 <= w_d2; end if;
        if w_a2 = 775 then w775 <= w_d2; end if;
        if w_a2 = 776 then w776 <= w_d2; end if;
        if w_a2 = 777 then w777 <= w_d2; end if;
        if w_a2 = 778 then w778 <= w_d2; end if;
        if w_a2 = 779 then w779 <= w_d2; end if;
        if w_a2 = 781 then w781 <= w_d2; end if;
        if w_a2 = 782 then w782 <= w_d2; end if;
        if w_a2 = 783 then w783 <= w_d2; end if;
        if w_a2 = 784 then w784 <= w_d2; end if;
        if w_a2 = 785 then w785 <= w_d2; end if;
        if w_a2 = 786 then w786 <= w_d2; end if;
        if w_a2 = 787 then w787 <= w_d2; end if;
        if w_a2 = 788 then w788 <= w_d2; end if;
        if w_a2 = 789 then w789 <= w_d2; end if;
        if w_a2 = 791 then w791 <= w_d2; end if;
        if w_a2 = 792 then w792 <= w_d2; end if;
        if w_a2 = 793 then w793 <= w_d2; end if;
        if w_a2 = 794 then w794 <= w_d2; end if;
        if w_a2 = 795 then w795 <= w_d2; end if;
        if w_a2 = 796 then w796 <= w_d2; end if;
        if w_a2 = 797 then w797 <= w_d2; end if;
        if w_a2 = 798 then w798 <= w_d2; end if;
        if w_a2 = 799 then w799 <= w_d2; end if;
        if w_a2 = 801 then w801 <= w_d2; end if;
        if w_a2 = 802 then w802 <= w_d2; end if;
        if w_a2 = 803 then w803 <= w_d2; end if;
        if w_a2 = 804 then w804 <= w_d2; end if;
        if w_a2 = 805 then w805 <= w_d2; end if;
        if w_a2 = 806 then w806 <= w_d2; end if;
        if w_a2 = 807 then w807 <= w_d2; end if;
        if w_a2 = 808 then w808 <= w_d2; end if;
        if w_a2 = 809 then w809 <= w_d2; end if;
        if w_a2 = 811 then w811 <= w_d2; end if;
        if w_a2 = 812 then w812 <= w_d2; end if;
        if w_a2 = 813 then w813 <= w_d2; end if;
        if w_a2 = 814 then w814 <= w_d2; end if;
        if w_a2 = 815 then w815 <= w_d2; end if;
        if w_a2 = 816 then w816 <= w_d2; end if;
        if w_a2 = 817 then w817 <= w_d2; end if;
        if w_a2 = 818 then w818 <= w_d2; end if;
        if w_a2 = 819 then w819 <= w_d2; end if;
        if w_a2 = 821 then w821 <= w_d2; end if;
        if w_a2 = 822 then w822 <= w_d2; end if;
        if w_a2 = 823 then w823 <= w_d2; end if;
        if w_a2 = 824 then w824 <= w_d2; end if;
        if w_a2 = 825 then w825 <= w_d2; end if;
        if w_a2 = 826 then w826 <= w_d2; end if;
        if w_a2 = 827 then w827 <= w_d2; end if;
        if w_a2 = 828 then w828 <= w_d2; end if;
        if w_a2 = 829 then w829 <= w_d2; end if;
        if w_a2 = 831 then w831 <= w_d2; end if;
        if w_a2 = 832 then w832 <= w_d2; end if;
        if w_a2 = 833 then w833 <= w_d2; end if;
        if w_a2 = 834 then w834 <= w_d2; end if;
        if w_a2 = 835 then w835 <= w_d2; end if;
        if w_a2 = 836 then w836 <= w_d2; end if;
        if w_a2 = 837 then w837 <= w_d2; end if;
        if w_a2 = 838 then w838 <= w_d2; end if;
        if w_a2 = 839 then w839 <= w_d2; end if;
        if w_a2 = 841 then w841 <= w_d2; end if;
        if w_a2 = 842 then w842 <= w_d2; end if;
        if w_a2 = 843 then w843 <= w_d2; end if;
        if w_a2 = 844 then w844 <= w_d2; end if;
        if w_a2 = 845 then w845 <= w_d2; end if;
        if w_a2 = 846 then w846 <= w_d2; end if;
        if w_a2 = 847 then w847 <= w_d2; end if;
        if w_a2 = 848 then w848 <= w_d2; end if;
        if w_a2 = 849 then w849 <= w_d2; end if;
        if w_a2 = 851 then w851 <= w_d2; end if;
        if w_a2 = 852 then w852 <= w_d2; end if;
        if w_a2 = 853 then w853 <= w_d2; end if;
        if w_a2 = 854 then w854 <= w_d2; end if;
        if w_a2 = 855 then w855 <= w_d2; end if;
        if w_a2 = 856 then w856 <= w_d2; end if;
        if w_a2 = 857 then w857 <= w_d2; end if;
        if w_a2 = 858 then w858 <= w_d2; end if;
        if w_a2 = 859 then w859 <= w_d2; end if;
        if w_a2 = 861 then w861 <= w_d2; end if;
        if w_a2 = 862 then w862 <= w_d2; end if;
        if w_a2 = 863 then w863 <= w_d2; end if;
        if w_a2 = 864 then w864 <= w_d2; end if;
        if w_a2 = 865 then w865 <= w_d2; end if;
        if w_a2 = 866 then w866 <= w_d2; end if;
        if w_a2 = 867 then w867 <= w_d2; end if;
        if w_a2 = 868 then w868 <= w_d2; end if;
        if w_a2 = 869 then w869 <= w_d2; end if;
        if w_a2 = 871 then w871 <= w_d2; end if;
        if w_a2 = 872 then w872 <= w_d2; end if;
        if w_a2 = 873 then w873 <= w_d2; end if;
        if w_a2 = 874 then w874 <= w_d2; end if;
        if w_a2 = 875 then w875 <= w_d2; end if;
        if w_a2 = 876 then w876 <= w_d2; end if;
        if w_a2 = 877 then w877 <= w_d2; end if;
        if w_a2 = 878 then w878 <= w_d2; end if;
        if w_a2 = 879 then w879 <= w_d2; end if;
        if w_a2 = 881 then w881 <= w_d2; end if;
        if w_a2 = 882 then w882 <= w_d2; end if;
        if w_a2 = 883 then w883 <= w_d2; end if;
        if w_a2 = 884 then w884 <= w_d2; end if;
        if w_a2 = 885 then w885 <= w_d2; end if;
        if w_a2 = 886 then w886 <= w_d2; end if;
        if w_a2 = 887 then w887 <= w_d2; end if;
        if w_a2 = 888 then w888 <= w_d2; end if;
        if w_a2 = 889 then w889 <= w_d2; end if;
        if w_a2 = 891 then w891 <= w_d2; end if;
        if w_a2 = 892 then w892 <= w_d2; end if;
        if w_a2 = 893 then w893 <= w_d2; end if;
        if w_a2 = 894 then w894 <= w_d2; end if;
        if w_a2 = 895 then w895 <= w_d2; end if;
        if w_a2 = 896 then w896 <= w_d2; end if;
        if w_a2 = 897 then w897 <= w_d2; end if;
        if w_a2 = 898 then w898 <= w_d2; end if;
        if w_a2 = 899 then w899 <= w_d2; end if;
        if w_a2 = 901 then w901 <= w_d2; end if;
        if w_a2 = 902 then w902 <= w_d2; end if;
        if w_a2 = 903 then w903 <= w_d2; end if;
        if w_a2 = 904 then w904 <= w_d2; end if;
        if w_a2 = 905 then w905 <= w_d2; end if;
        if w_a2 = 906 then w906 <= w_d2; end if;
        if w_a2 = 907 then w907 <= w_d2; end if;
        if w_a2 = 908 then w908 <= w_d2; end if;
        if w_a2 = 909 then w909 <= w_d2; end if;
        if w_a2 = 911 then w911 <= w_d2; end if;
        if w_a2 = 912 then w912 <= w_d2; end if;
        if w_a2 = 913 then w913 <= w_d2; end if;
        if w_a2 = 914 then w914 <= w_d2; end if;
        if w_a2 = 915 then w915 <= w_d2; end if;
        if w_a2 = 916 then w916 <= w_d2; end if;
        if w_a2 = 917 then w917 <= w_d2; end if;
        if w_a2 = 918 then w918 <= w_d2; end if;
        if w_a2 = 919 then w919 <= w_d2; end if;
        if w_a2 = 921 then w921 <= w_d2; end if;
        if w_a2 = 922 then w922 <= w_d2; end if;
        if w_a2 = 923 then w923 <= w_d2; end if;
        if w_a2 = 924 then w924 <= w_d2; end if;
        if w_a2 = 925 then w925 <= w_d2; end if;
        if w_a2 = 926 then w926 <= w_d2; end if;
        if w_a2 = 927 then w927 <= w_d2; end if;
        if w_a2 = 928 then w928 <= w_d2; end if;
        if w_a2 = 929 then w929 <= w_d2; end if;
        if w_a2 = 931 then w931 <= w_d2; end if;
        if w_a2 = 932 then w932 <= w_d2; end if;
        if w_a2 = 933 then w933 <= w_d2; end if;
        if w_a2 = 934 then w934 <= w_d2; end if;
        if w_a2 = 935 then w935 <= w_d2; end if;
        if w_a2 = 936 then w936 <= w_d2; end if;
        if w_a2 = 937 then w937 <= w_d2; end if;
        if w_a2 = 938 then w938 <= w_d2; end if;
        if w_a2 = 939 then w939 <= w_d2; end if;
        if w_a2 = 941 then w941 <= w_d2; end if;
        if w_a2 = 942 then w942 <= w_d2; end if;
        if w_a2 = 943 then w943 <= w_d2; end if;
        if w_a2 = 944 then w944 <= w_d2; end if;
        if w_a2 = 945 then w945 <= w_d2; end if;
        if w_a2 = 946 then w946 <= w_d2; end if;
        if w_a2 = 947 then w947 <= w_d2; end if;
        if w_a2 = 948 then w948 <= w_d2; end if;
        if w_a2 = 949 then w949 <= w_d2; end if;
        if w_a2 = 951 then w951 <= w_d2; end if;
        if w_a2 = 952 then w952 <= w_d2; end if;
        if w_a2 = 953 then w953 <= w_d2; end if;
        if w_a2 = 954 then w954 <= w_d2; end if;
        if w_a2 = 955 then w955 <= w_d2; end if;
        if w_a2 = 956 then w956 <= w_d2; end if;
        if w_a2 = 957 then w957 <= w_d2; end if;
        if w_a2 = 958 then w958 <= w_d2; end if;
        if w_a2 = 959 then w959 <= w_d2; end if;
        if w_a2 = 961 then w961 <= w_d2; end if;
        if w_a2 = 962 then w962 <= w_d2; end if;
        if w_a2 = 963 then w963 <= w_d2; end if;
        if w_a2 = 964 then w964 <= w_d2; end if;
        if w_a2 = 965 then w965 <= w_d2; end if;
        if w_a2 = 966 then w966 <= w_d2; end if;
        if w_a2 = 967 then w967 <= w_d2; end if;
        if w_a2 = 968 then w968 <= w_d2; end if;
        if w_a2 = 969 then w969 <= w_d2; end if;
        if w_a2 = 971 then w971 <= w_d2; end if;
        if w_a2 = 972 then w972 <= w_d2; end if;
        if w_a2 = 973 then w973 <= w_d2; end if;
        if w_a2 = 974 then w974 <= w_d2; end if;
        if w_a2 = 975 then w975 <= w_d2; end if;
        if w_a2 = 976 then w976 <= w_d2; end if;
        if w_a2 = 977 then w977 <= w_d2; end if;
        if w_a2 = 978 then w978 <= w_d2; end if;
        if w_a2 = 979 then w979 <= w_d2; end if;
        if w_a2 = 981 then w981 <= w_d2; end if;
        if w_a2 = 982 then w982 <= w_d2; end if;
        if w_a2 = 983 then w983 <= w_d2; end if;
        if w_a2 = 984 then w984 <= w_d2; end if;
        if w_a2 = 985 then w985 <= w_d2; end if;
        if w_a2 = 986 then w986 <= w_d2; end if;
        if w_a2 = 987 then w987 <= w_d2; end if;
        if w_a2 = 988 then w988 <= w_d2; end if;
        if w_a2 = 989 then w989 <= w_d2; end if;
        if w_a2 = 991 then w991 <= w_d2; end if;
        if w_a2 = 992 then w992 <= w_d2; end if;
        if w_a2 = 993 then w993 <= w_d2; end if;
        if w_a2 = 994 then w994 <= w_d2; end if;
        if w_a2 = 995 then w995 <= w_d2; end if;
        if w_a2 = 996 then w996 <= w_d2; end if;
        if w_a2 = 997 then w997 <= w_d2; end if;
        if w_a2 = 998 then w998 <= w_d2; end if;
        if w_a2 = 999 then w999 <= w_d2; end if;
      end if;
    end if;
  end process weigth_encoder2;

inst0: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w001       ,
      w02      => w002       ,
      w03      => w003       ,
      w04      => w004       ,
      w05      => w005       ,
      w06      => w006       ,
      w07      => w007       ,
      w08      => w008       ,
      w09      => w009       ,
      w11      => w011       ,
      w12      => w012       ,
      w13      => w013       ,
      w14      => w014       ,
      w15      => w015       ,
      w16      => w016       ,
      w17      => w017       ,
      w18      => w018       ,
      w19      => w019       ,
      w21      => w021       ,
      w22      => w022       ,
      w23      => w023       ,
      w24      => w024       ,
      w25      => w025       ,
      w26      => w026       ,
      w27      => w027       ,
      w28      => w028       ,
      w29      => w029       ,
      w31      => w031       ,
      w32      => w032       ,
      w33      => w033       ,
      w34      => w034       ,
      w35      => w035       ,
      w36      => w036       ,
      w37      => w037       ,
      w38      => w038       ,
      w39      => w039       ,
      w41      => w041       ,
      w42      => w042       ,
      w43      => w043       ,
      w44      => w044       ,
      w45      => w045       ,
      w46      => w046       ,
      w47      => w047       ,
      w48      => w048       ,
      w49      => w049       ,
      w51      => w051       ,
      w52      => w052       ,
      w53      => w053       ,
      w54      => w054       ,
      w55      => w055       ,
      w56      => w056       ,
      w57      => w057       ,
      w58      => w058       ,
      w59      => w059       ,
      w61      => w061       ,
      w62      => w062       ,
      w63      => w063       ,
      w64      => w064       ,
      w65      => w065       ,
      w66      => w066       ,
      w67      => w067       ,
      w68      => w068       ,
      w69      => w069       ,
      w71      => w071       ,
      w72      => w072       ,
      w73      => w073       ,
      w74      => w074       ,
      w75      => w075       ,
      w76      => w076       ,
      w77      => w077       ,
      w78      => w078       ,
      w79      => w079       ,
      w81      => w081       ,
      w82      => w082       ,
      w83      => w083       ,
      w84      => w084       ,
      w85      => w085       ,
      w86      => w086       ,
      w87      => w087       ,
      w88      => w088       ,
      w89      => w089       ,
      w91      => w091       ,
      w92      => w092       ,
      w93      => w093       ,
      w94      => w094       ,
      w95      => w095       ,
      w96      => w096       ,
      w97      => w097       ,
      w98      => w098       ,
      w99      => w099       ,
      d_out   => max0_out          ,
      en_out  => en_out         ,
      sof_out => sof0             
    );


inst1: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in       ,
      en_in   => en_in      ,
      sof_in  => sof_in     ,

      w01      => w101       ,
      w02      => w102       ,
      w03      => w103       ,
      w04      => w104       ,
      w05      => w105       ,
      w06      => w106       ,
      w07      => w107       ,
      w08      => w108       ,
      w09      => w109       ,
      w11      => w111       ,
      w12      => w112       ,
      w13      => w113       ,
      w14      => w114       ,
      w15      => w115       ,
      w16      => w116       ,
      w17      => w117       ,
      w18      => w118       ,
      w19      => w119       ,
      w21      => w121       ,
      w22      => w122       ,
      w23      => w123       ,
      w24      => w124       ,
      w25      => w125       ,
      w26      => w126       ,
      w27      => w127       ,
      w28      => w128       ,
      w29      => w129       ,
      w31      => w131       ,
      w32      => w132       ,
      w33      => w133       ,
      w34      => w134       ,
      w35      => w135       ,
      w36      => w136       ,
      w37      => w137       ,
      w38      => w138       ,
      w39      => w139       ,
      w41      => w141       ,
      w42      => w142       ,
      w43      => w143       ,
      w44      => w144       ,
      w45      => w145       ,
      w46      => w146       ,
      w47      => w147       ,
      w48      => w148       ,
      w49      => w149       ,
      w51      => w151       ,
      w52      => w152       ,
      w53      => w153       ,
      w54      => w154       ,
      w55      => w155       ,
      w56      => w156       ,
      w57      => w157       ,
      w58      => w158       ,
      w59      => w159       ,
      w61      => w161       ,
      w62      => w162       ,
      w63      => w163       ,
      w64      => w164       ,
      w65      => w165       ,
      w66      => w166       ,
      w67      => w167       ,
      w68      => w168       ,
      w69      => w169       ,
      w71      => w171       ,
      w72      => w172       ,
      w73      => w173       ,
      w74      => w174       ,
      w75      => w175       ,
      w76      => w176       ,
      w77      => w177       ,
      w78      => w178       ,
      w79      => w179       ,
      w81      => w181       ,
      w82      => w182       ,
      w83      => w183       ,
      w84      => w184       ,
      w85      => w185       ,
      w86      => w186       ,
      w87      => w187       ,
      w88      => w188       ,
      w89      => w189       ,
      w91      => w191       ,
      w92      => w192       ,
      w93      => w193       ,
      w94      => w194       ,
      w95      => w195       ,
      w96      => w196       ,
      w97      => w197       ,
      w98      => w198       ,
      w99      => w199       ,
      d_out   => max1_out    ,
      en_out  => en1   ,
      sof_out => sof1             
    );



inst2: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in       ,
      en_in   => en_in      ,
      sof_in  => sof_in     ,

      w01      => w201       ,
      w02      => w202       ,
      w03      => w203       ,
      w04      => w204       ,
      w05      => w205       ,
      w06      => w206       ,
      w07      => w207       ,
      w08      => w208       ,
      w09      => w209       ,
      w11      => w211       ,
      w12      => w212       ,
      w13      => w213       ,
      w14      => w214       ,
      w15      => w215       ,
      w16      => w216       ,
      w17      => w217       ,
      w18      => w218       ,
      w19      => w219       ,
      w21      => w221       ,
      w22      => w222       ,
      w23      => w223       ,
      w24      => w224       ,
      w25      => w225       ,
      w26      => w226       ,
      w27      => w227       ,
      w28      => w228       ,
      w29      => w229       ,
      w31      => w231       ,
      w32      => w232       ,
      w33      => w233       ,
      w34      => w234       ,
      w35      => w235       ,
      w36      => w236       ,
      w37      => w237       ,
      w38      => w238       ,
      w39      => w239       ,
      w41      => w241       ,
      w42      => w242       ,
      w43      => w243       ,
      w44      => w244       ,
      w45      => w245       ,
      w46      => w246       ,
      w47      => w247       ,
      w48      => w248       ,
      w49      => w249       ,
      w51      => w251       ,
      w52      => w252       ,
      w53      => w253       ,
      w54      => w254       ,
      w55      => w255       ,
      w56      => w256       ,
      w57      => w257       ,
      w58      => w258       ,
      w59      => w259       ,
      w61      => w261       ,
      w62      => w262       ,
      w63      => w263       ,
      w64      => w264       ,
      w65      => w265       ,
      w66      => w266       ,
      w67      => w267       ,
      w68      => w268       ,
      w69      => w269       ,
      w71      => w271       ,
      w72      => w272       ,
      w73      => w273       ,
      w74      => w274       ,
      w75      => w275       ,
      w76      => w276       ,
      w77      => w277       ,
      w78      => w278       ,
      w79      => w279       ,
      w81      => w281       ,
      w82      => w282       ,
      w83      => w283       ,
      w84      => w284       ,
      w85      => w285       ,
      w86      => w286       ,
      w87      => w287       ,
      w88      => w288       ,
      w89      => w289       ,
      w91      => w291       ,
      w92      => w292       ,
      w93      => w293       ,
      w94      => w294       ,
      w95      => w295       ,
      w96      => w296       ,
      w97      => w297       ,
      w98      => w298       ,
      w99      => w299       ,
      d_out   => max2_out    ,
      en_out  => en2   ,
      sof_out => sof2             
    );



inst3: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w301       ,
      w02      => w302       ,
      w03      => w303       ,
      w04      => w304       ,
      w05      => w305       ,
      w06      => w306       ,
      w07      => w307       ,
      w08      => w308       ,
      w09      => w309       ,
      w11      => w311       ,
      w12      => w312       ,
      w13      => w313       ,
      w14      => w314       ,
      w15      => w315       ,
      w16      => w316       ,
      w17      => w317       ,
      w18      => w318       ,
      w19      => w319       ,
      w21      => w321       ,
      w22      => w322       ,
      w23      => w323       ,
      w24      => w324       ,
      w25      => w325       ,
      w26      => w326       ,
      w27      => w327       ,
      w28      => w328       ,
      w29      => w329       ,
      w31      => w331       ,
      w32      => w332       ,
      w33      => w333       ,
      w34      => w334       ,
      w35      => w335       ,
      w36      => w336       ,
      w37      => w337       ,
      w38      => w338       ,
      w39      => w339       ,
      w41      => w341       ,
      w42      => w342       ,
      w43      => w343       ,
      w44      => w344       ,
      w45      => w345       ,
      w46      => w346       ,
      w47      => w347       ,
      w48      => w348       ,
      w49      => w349       ,
      w51      => w351       ,
      w52      => w352       ,
      w53      => w353       ,
      w54      => w354       ,
      w55      => w355       ,
      w56      => w356       ,
      w57      => w357       ,
      w58      => w358       ,
      w59      => w359       ,
      w61      => w361       ,
      w62      => w362       ,
      w63      => w363       ,
      w64      => w364       ,
      w65      => w365       ,
      w66      => w366       ,
      w67      => w367       ,
      w68      => w368       ,
      w69      => w369       ,
      w71      => w371       ,
      w72      => w372       ,
      w73      => w373       ,
      w74      => w374       ,
      w75      => w375       ,
      w76      => w376       ,
      w77      => w377       ,
      w78      => w378       ,
      w79      => w379       ,
      w81      => w381       ,
      w82      => w382       ,
      w83      => w383       ,
      w84      => w384       ,
      w85      => w385       ,
      w86      => w386       ,
      w87      => w387       ,
      w88      => w388       ,
      w89      => w389       ,
      w91      => w391       ,
      w92      => w392       ,
      w93      => w393       ,
      w94      => w394       ,
      w95      => w395       ,
      w96      => w396       ,
      w97      => w397       ,
      w98      => w398       ,
      w99      => w399       ,
      d_out   => max3_out    ,
      en_out  => en3   ,
      sof_out => sof3             
    );



inst4: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w401       ,
      w02      => w402       ,
      w03      => w403       ,
      w04      => w404       ,
      w05      => w405       ,
      w06      => w406       ,
      w07      => w407       ,
      w08      => w408       ,
      w09      => w409       ,
      w11      => w411       ,
      w12      => w412       ,
      w13      => w413       ,
      w14      => w414       ,
      w15      => w415       ,
      w16      => w416       ,
      w17      => w417       ,
      w18      => w418       ,
      w19      => w419       ,
      w21      => w421       ,
      w22      => w422       ,
      w23      => w423       ,
      w24      => w424       ,
      w25      => w425       ,
      w26      => w426       ,
      w27      => w427       ,
      w28      => w428       ,
      w29      => w429       ,
      w31      => w431       ,
      w32      => w432       ,
      w33      => w433       ,
      w34      => w434       ,
      w35      => w435       ,
      w36      => w436       ,
      w37      => w437       ,
      w38      => w438       ,
      w39      => w439       ,
      w41      => w441       ,
      w42      => w442       ,
      w43      => w443       ,
      w44      => w444       ,
      w45      => w445       ,
      w46      => w446       ,
      w47      => w447       ,
      w48      => w448       ,
      w49      => w449       ,
      w51      => w451       ,
      w52      => w452       ,
      w53      => w453       ,
      w54      => w454       ,
      w55      => w455       ,
      w56      => w456       ,
      w57      => w457       ,
      w58      => w458       ,
      w59      => w459       ,
      w61      => w461       ,
      w62      => w462       ,
      w63      => w463       ,
      w64      => w464       ,
      w65      => w465       ,
      w66      => w466       ,
      w67      => w467       ,
      w68      => w468       ,
      w69      => w469       ,
      w71      => w471       ,
      w72      => w472       ,
      w73      => w473       ,
      w74      => w474       ,
      w75      => w475       ,
      w76      => w476       ,
      w77      => w477       ,
      w78      => w478       ,
      w79      => w479       ,
      w81      => w481       ,
      w82      => w482       ,
      w83      => w483       ,
      w84      => w484       ,
      w85      => w485       ,
      w86      => w486       ,
      w87      => w487       ,
      w88      => w488       ,
      w89      => w489       ,
      w91      => w491       ,
      w92      => w492       ,
      w93      => w493       ,
      w94      => w494       ,
      w95      => w495       ,
      w96      => w496       ,
      w97      => w497       ,
      w98      => w498       ,
      w99      => w499       ,
      d_out   => max4_out    ,
      en_out  => en4   ,
      sof_out => sof4             
    );



inst5: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w501       ,
      w02      => w502       ,
      w03      => w503       ,
      w04      => w504       ,
      w05      => w505       ,
      w06      => w506       ,
      w07      => w507       ,
      w08      => w508       ,
      w09      => w509       ,
      w11      => w511       ,
      w12      => w512       ,
      w13      => w513       ,
      w14      => w514       ,
      w15      => w515       ,
      w16      => w516       ,
      w17      => w517       ,
      w18      => w518       ,
      w19      => w519       ,
      w21      => w521       ,
      w22      => w522       ,
      w23      => w523       ,
      w24      => w524       ,
      w25      => w525       ,
      w26      => w526       ,
      w27      => w527       ,
      w28      => w528       ,
      w29      => w529       ,
      w31      => w531       ,
      w32      => w532       ,
      w33      => w533       ,
      w34      => w534       ,
      w35      => w535       ,
      w36      => w536       ,
      w37      => w537       ,
      w38      => w538       ,
      w39      => w539       ,
      w41      => w541       ,
      w42      => w542       ,
      w43      => w543       ,
      w44      => w544       ,
      w45      => w545       ,
      w46      => w546       ,
      w47      => w547       ,
      w48      => w548       ,
      w49      => w549       ,
      w51      => w551       ,
      w52      => w552       ,
      w53      => w553       ,
      w54      => w554       ,
      w55      => w555       ,
      w56      => w556       ,
      w57      => w557       ,
      w58      => w558       ,
      w59      => w559       ,
      w61      => w561       ,
      w62      => w562       ,
      w63      => w563       ,
      w64      => w564       ,
      w65      => w565       ,
      w66      => w566       ,
      w67      => w567       ,
      w68      => w568       ,
      w69      => w569       ,
      w71      => w571       ,
      w72      => w572       ,
      w73      => w573       ,
      w74      => w574       ,
      w75      => w575       ,
      w76      => w576       ,
      w77      => w577       ,
      w78      => w578       ,
      w79      => w579       ,
      w81      => w581       ,
      w82      => w582       ,
      w83      => w583       ,
      w84      => w584       ,
      w85      => w585       ,
      w86      => w586       ,
      w87      => w587       ,
      w88      => w588       ,
      w89      => w589       ,
      w91      => w591       ,
      w92      => w592       ,
      w93      => w593       ,
      w94      => w594       ,
      w95      => w595       ,
      w96      => w596       ,
      w97      => w597       ,
      w98      => w598       ,
      w99      => w599       ,
      d_out   => max5_out    ,
      en_out  => en5   ,
      sof_out => sof5             
    );



inst6: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w601       ,
      w02      => w602       ,
      w03      => w603       ,
      w04      => w604       ,
      w05      => w605       ,
      w06      => w606       ,
      w07      => w607       ,
      w08      => w608       ,
      w09      => w609       ,
      w11      => w611       ,
      w12      => w612       ,
      w13      => w613       ,
      w14      => w614       ,
      w15      => w615       ,
      w16      => w616       ,
      w17      => w617       ,
      w18      => w618       ,
      w19      => w619       ,
      w21      => w621       ,
      w22      => w622       ,
      w23      => w623       ,
      w24      => w624       ,
      w25      => w625       ,
      w26      => w626       ,
      w27      => w627       ,
      w28      => w628       ,
      w29      => w629       ,
      w31      => w631       ,
      w32      => w632       ,
      w33      => w633       ,
      w34      => w634       ,
      w35      => w635       ,
      w36      => w636       ,
      w37      => w637       ,
      w38      => w638       ,
      w39      => w639       ,
      w41      => w641       ,
      w42      => w642       ,
      w43      => w643       ,
      w44      => w644       ,
      w45      => w645       ,
      w46      => w646       ,
      w47      => w647       ,
      w48      => w648       ,
      w49      => w649       ,
      w51      => w651       ,
      w52      => w652       ,
      w53      => w653       ,
      w54      => w654       ,
      w55      => w655       ,
      w56      => w656       ,
      w57      => w657       ,
      w58      => w658       ,
      w59      => w659       ,
      w61      => w661       ,
      w62      => w662       ,
      w63      => w663       ,
      w64      => w664       ,
      w65      => w665       ,
      w66      => w666       ,
      w67      => w667       ,
      w68      => w668       ,
      w69      => w669       ,
      w71      => w671       ,
      w72      => w672       ,
      w73      => w673       ,
      w74      => w674       ,
      w75      => w675       ,
      w76      => w676       ,
      w77      => w677       ,
      w78      => w678       ,
      w79      => w679       ,
      w81      => w681       ,
      w82      => w682       ,
      w83      => w683       ,
      w84      => w684       ,
      w85      => w685       ,
      w86      => w686       ,
      w87      => w687       ,
      w88      => w688       ,
      w89      => w689       ,
      w91      => w691       ,
      w92      => w692       ,
      w93      => w693       ,
      w94      => w694       ,
      w95      => w695       ,
      w96      => w696       ,
      w97      => w697       ,
      w98      => w698       ,
      w99      => w699       ,
      d_out   => max6_out    ,
      en_out  => en6   ,
      sof_out => sof6             
    );



inst7: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w701       ,
      w02      => w702       ,
      w03      => w703       ,
      w04      => w704       ,
      w05      => w705       ,
      w06      => w706       ,
      w07      => w707       ,
      w08      => w708       ,
      w09      => w709       ,
      w11      => w711       ,
      w12      => w712       ,
      w13      => w713       ,
      w14      => w714       ,
      w15      => w715       ,
      w16      => w716       ,
      w17      => w717       ,
      w18      => w718       ,
      w19      => w719       ,
      w21      => w721       ,
      w22      => w722       ,
      w23      => w723       ,
      w24      => w724       ,
      w25      => w725       ,
      w26      => w726       ,
      w27      => w727       ,
      w28      => w728       ,
      w29      => w729       ,
      w31      => w731       ,
      w32      => w732       ,
      w33      => w733       ,
      w34      => w734       ,
      w35      => w735       ,
      w36      => w736       ,
      w37      => w737       ,
      w38      => w738       ,
      w39      => w739       ,
      w41      => w741       ,
      w42      => w742       ,
      w43      => w743       ,
      w44      => w744       ,
      w45      => w745       ,
      w46      => w746       ,
      w47      => w747       ,
      w48      => w748       ,
      w49      => w749       ,
      w51      => w751       ,
      w52      => w752       ,
      w53      => w753       ,
      w54      => w754       ,
      w55      => w755       ,
      w56      => w756       ,
      w57      => w757       ,
      w58      => w758       ,
      w59      => w759       ,
      w61      => w761       ,
      w62      => w762       ,
      w63      => w763       ,
      w64      => w764       ,
      w65      => w765       ,
      w66      => w766       ,
      w67      => w767       ,
      w68      => w768       ,
      w69      => w769       ,
      w71      => w771       ,
      w72      => w772       ,
      w73      => w773       ,
      w74      => w774       ,
      w75      => w775       ,
      w76      => w776       ,
      w77      => w777       ,
      w78      => w778       ,
      w79      => w779       ,
      w81      => w781       ,
      w82      => w782       ,
      w83      => w783       ,
      w84      => w784       ,
      w85      => w785       ,
      w86      => w786       ,
      w87      => w787       ,
      w88      => w788       ,
      w89      => w789       ,
      w91      => w791       ,
      w92      => w792       ,
      w93      => w793       ,
      w94      => w794       ,
      w95      => w795       ,
      w96      => w796       ,
      w97      => w797       ,
      w98      => w798       ,
      w99      => w799       ,
      d_out   => max7_out    ,
      en_out  => en7   ,
      sof_out => sof7             
    );



inst8: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w801       ,
      w02      => w802       ,
      w03      => w803       ,
      w04      => w804       ,
      w05      => w805       ,
      w06      => w806       ,
      w07      => w807       ,
      w08      => w808       ,
      w09      => w809       ,
      w11      => w811       ,
      w12      => w812       ,
      w13      => w813       ,
      w14      => w814       ,
      w15      => w815       ,
      w16      => w816       ,
      w17      => w817       ,
      w18      => w818       ,
      w19      => w819       ,
      w21      => w821       ,
      w22      => w822       ,
      w23      => w823       ,
      w24      => w824       ,
      w25      => w825       ,
      w26      => w826       ,
      w27      => w827       ,
      w28      => w828       ,
      w29      => w829       ,
      w31      => w831       ,
      w32      => w832       ,
      w33      => w833       ,
      w34      => w834       ,
      w35      => w835       ,
      w36      => w836       ,
      w37      => w837       ,
      w38      => w838       ,
      w39      => w839       ,
      w41      => w841       ,
      w42      => w842       ,
      w43      => w843       ,
      w44      => w844       ,
      w45      => w845       ,
      w46      => w846       ,
      w47      => w847       ,
      w48      => w848       ,
      w49      => w849       ,
      w51      => w851       ,
      w52      => w852       ,
      w53      => w853       ,
      w54      => w854       ,
      w55      => w855       ,
      w56      => w856       ,
      w57      => w857       ,
      w58      => w858       ,
      w59      => w859       ,
      w61      => w861       ,
      w62      => w862       ,
      w63      => w863       ,
      w64      => w864       ,
      w65      => w865       ,
      w66      => w866       ,
      w67      => w867       ,
      w68      => w868       ,
      w69      => w869       ,
      w71      => w871       ,
      w72      => w872       ,
      w73      => w873       ,
      w74      => w874       ,
      w75      => w875       ,
      w76      => w876       ,
      w77      => w877       ,
      w78      => w878       ,
      w79      => w879       ,
      w81      => w881       ,
      w82      => w882       ,
      w83      => w883       ,
      w84      => w884       ,
      w85      => w885       ,
      w86      => w886       ,
      w87      => w887       ,
      w88      => w888       ,
      w89      => w889       ,
      w91      => w891       ,
      w92      => w892       ,
      w93      => w893       ,
      w94      => w894       ,
      w95      => w895       ,
      w96      => w896       ,
      w97      => w897       ,
      w98      => w898       ,
      w99      => w899       ,
      d_out   => max8_out    ,
      en_out  => en8  ,
      sof_out => sof8            
    );



inst9: ConvLayersN generic map (
      mult_sum => mult_sum,
      N        => N       , -- input data width
      M        => M       , -- input data width
      W        => W       ,-- output data width
      SR       => SR      ,-- output data shift right

      in_row   => in_row  ,
      in_col   => in_col
      )
port map (
      clk     => clk      ,
      rst     => rst      ,
      d_in    => d_in     ,
      en_in   => en_in    ,
      sof_in  => sof_in   ,

      w01      => w901       ,
      w02      => w902       ,
      w03      => w903       ,
      w04      => w904       ,
      w05      => w905       ,
      w06      => w906       ,
      w07      => w907       ,
      w08      => w908       ,
      w09      => w909       ,
      w11      => w911       ,
      w12      => w912       ,
      w13      => w913       ,
      w14      => w914       ,
      w15      => w915       ,
      w16      => w916       ,
      w17      => w917       ,
      w18      => w918       ,
      w19      => w919       ,
      w21      => w921       ,
      w22      => w922       ,
      w23      => w923       ,
      w24      => w924       ,
      w25      => w925       ,
      w26      => w926       ,
      w27      => w927       ,
      w28      => w928       ,
      w29      => w929       ,
      w31      => w931       ,
      w32      => w932       ,
      w33      => w933       ,
      w34      => w934       ,
      w35      => w935       ,
      w36      => w936       ,
      w37      => w937       ,
      w38      => w938       ,
      w39      => w939       ,
      w41      => w941       ,
      w42      => w942       ,
      w43      => w943       ,
      w44      => w944       ,
      w45      => w945       ,
      w46      => w946       ,
      w47      => w947       ,
      w48      => w948       ,
      w49      => w949       ,
      w51      => w951       ,
      w52      => w952       ,
      w53      => w953       ,
      w54      => w954       ,
      w55      => w955       ,
      w56      => w956       ,
      w57      => w957       ,
      w58      => w958       ,
      w59      => w959       ,
      w61      => w961       ,
      w62      => w962       ,
      w63      => w963       ,
      w64      => w964       ,
      w65      => w965       ,
      w66      => w966       ,
      w67      => w967       ,
      w68      => w968       ,
      w69      => w969       ,
      w71      => w971       ,
      w72      => w972       ,
      w73      => w973       ,
      w74      => w974       ,
      w75      => w975       ,
      w76      => w976       ,
      w77      => w977       ,
      w78      => w978       ,
      w79      => w979       ,
      w81      => w981       ,
      w82      => w982       ,
      w83      => w983       ,
      w84      => w984       ,
      w85      => w985       ,
      w86      => w986       ,
      w87      => w987       ,
      w88      => w988       ,
      w89      => w989       ,
      w91      => w991       ,
      w92      => w992       ,
      w93      => w993       ,
      w94      => w994       ,
      w95      => w995       ,
      w96      => w996       ,
      w97      => w997       ,
      w98      => w998       ,
      w99      => w999       ,
      d_out   => max9_out    ,
      en_out  => en9   ,
      sof_out => sof9             
    );


end a;