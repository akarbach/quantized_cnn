library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity multROM is
  port    (
           clk           : in  std_logic;

           ROM_addr      : in  std_logic_vector(15 downto 0);
           ROM_data      : out std_logic_vector(15 downto 0)
           );                        
end multROM;

architecture a of multROM is

    type ROM_Array is array (0 to (2**16-1)) 
  of std_logic_vector(15 downto 0);

    constant Content: ROM_Array := (
0 => conv_std_logic_vector(0, 16),
1 => conv_std_logic_vector(0, 16),
2 => conv_std_logic_vector(0, 16),
3 => conv_std_logic_vector(0, 16),
4 => conv_std_logic_vector(0, 16),
5 => conv_std_logic_vector(0, 16),
6 => conv_std_logic_vector(0, 16),
7 => conv_std_logic_vector(0, 16),
8 => conv_std_logic_vector(0, 16),
9 => conv_std_logic_vector(0, 16),
10 => conv_std_logic_vector(0, 16),
11 => conv_std_logic_vector(0, 16),
12 => conv_std_logic_vector(0, 16),
13 => conv_std_logic_vector(0, 16),
14 => conv_std_logic_vector(0, 16),
15 => conv_std_logic_vector(0, 16),
16 => conv_std_logic_vector(0, 16),
17 => conv_std_logic_vector(0, 16),
18 => conv_std_logic_vector(0, 16),
19 => conv_std_logic_vector(0, 16),
20 => conv_std_logic_vector(0, 16),
21 => conv_std_logic_vector(0, 16),
22 => conv_std_logic_vector(0, 16),
23 => conv_std_logic_vector(0, 16),
24 => conv_std_logic_vector(0, 16),
25 => conv_std_logic_vector(0, 16),
26 => conv_std_logic_vector(0, 16),
27 => conv_std_logic_vector(0, 16),
28 => conv_std_logic_vector(0, 16),
29 => conv_std_logic_vector(0, 16),
30 => conv_std_logic_vector(0, 16),
31 => conv_std_logic_vector(0, 16),
32 => conv_std_logic_vector(0, 16),
33 => conv_std_logic_vector(0, 16),
34 => conv_std_logic_vector(0, 16),
35 => conv_std_logic_vector(0, 16),
36 => conv_std_logic_vector(0, 16),
37 => conv_std_logic_vector(0, 16),
38 => conv_std_logic_vector(0, 16),
39 => conv_std_logic_vector(0, 16),
40 => conv_std_logic_vector(0, 16),
41 => conv_std_logic_vector(0, 16),
42 => conv_std_logic_vector(0, 16),
43 => conv_std_logic_vector(0, 16),
44 => conv_std_logic_vector(0, 16),
45 => conv_std_logic_vector(0, 16),
46 => conv_std_logic_vector(0, 16),
47 => conv_std_logic_vector(0, 16),
48 => conv_std_logic_vector(0, 16),
49 => conv_std_logic_vector(0, 16),
50 => conv_std_logic_vector(0, 16),
51 => conv_std_logic_vector(0, 16),
52 => conv_std_logic_vector(0, 16),
53 => conv_std_logic_vector(0, 16),
54 => conv_std_logic_vector(0, 16),
55 => conv_std_logic_vector(0, 16),
56 => conv_std_logic_vector(0, 16),
57 => conv_std_logic_vector(0, 16),
58 => conv_std_logic_vector(0, 16),
59 => conv_std_logic_vector(0, 16),
60 => conv_std_logic_vector(0, 16),
61 => conv_std_logic_vector(0, 16),
62 => conv_std_logic_vector(0, 16),
63 => conv_std_logic_vector(0, 16),
64 => conv_std_logic_vector(0, 16),
65 => conv_std_logic_vector(0, 16),
66 => conv_std_logic_vector(0, 16),
67 => conv_std_logic_vector(0, 16),
68 => conv_std_logic_vector(0, 16),
69 => conv_std_logic_vector(0, 16),
70 => conv_std_logic_vector(0, 16),
71 => conv_std_logic_vector(0, 16),
72 => conv_std_logic_vector(0, 16),
73 => conv_std_logic_vector(0, 16),
74 => conv_std_logic_vector(0, 16),
75 => conv_std_logic_vector(0, 16),
76 => conv_std_logic_vector(0, 16),
77 => conv_std_logic_vector(0, 16),
78 => conv_std_logic_vector(0, 16),
79 => conv_std_logic_vector(0, 16),
80 => conv_std_logic_vector(0, 16),
81 => conv_std_logic_vector(0, 16),
82 => conv_std_logic_vector(0, 16),
83 => conv_std_logic_vector(0, 16),
84 => conv_std_logic_vector(0, 16),
85 => conv_std_logic_vector(0, 16),
86 => conv_std_logic_vector(0, 16),
87 => conv_std_logic_vector(0, 16),
88 => conv_std_logic_vector(0, 16),
89 => conv_std_logic_vector(0, 16),
90 => conv_std_logic_vector(0, 16),
91 => conv_std_logic_vector(0, 16),
92 => conv_std_logic_vector(0, 16),
93 => conv_std_logic_vector(0, 16),
94 => conv_std_logic_vector(0, 16),
95 => conv_std_logic_vector(0, 16),
96 => conv_std_logic_vector(0, 16),
97 => conv_std_logic_vector(0, 16),
98 => conv_std_logic_vector(0, 16),
99 => conv_std_logic_vector(0, 16),
100 => conv_std_logic_vector(0, 16),
101 => conv_std_logic_vector(0, 16),
102 => conv_std_logic_vector(0, 16),
103 => conv_std_logic_vector(0, 16),
104 => conv_std_logic_vector(0, 16),
105 => conv_std_logic_vector(0, 16),
106 => conv_std_logic_vector(0, 16),
107 => conv_std_logic_vector(0, 16),
108 => conv_std_logic_vector(0, 16),
109 => conv_std_logic_vector(0, 16),
110 => conv_std_logic_vector(0, 16),
111 => conv_std_logic_vector(0, 16),
112 => conv_std_logic_vector(0, 16),
113 => conv_std_logic_vector(0, 16),
114 => conv_std_logic_vector(0, 16),
115 => conv_std_logic_vector(0, 16),
116 => conv_std_logic_vector(0, 16),
117 => conv_std_logic_vector(0, 16),
118 => conv_std_logic_vector(0, 16),
119 => conv_std_logic_vector(0, 16),
120 => conv_std_logic_vector(0, 16),
121 => conv_std_logic_vector(0, 16),
122 => conv_std_logic_vector(0, 16),
123 => conv_std_logic_vector(0, 16),
124 => conv_std_logic_vector(0, 16),
125 => conv_std_logic_vector(0, 16),
126 => conv_std_logic_vector(0, 16),
127 => conv_std_logic_vector(0, 16),
128 => conv_std_logic_vector(0, 16),
129 => conv_std_logic_vector(0, 16),
130 => conv_std_logic_vector(0, 16),
131 => conv_std_logic_vector(0, 16),
132 => conv_std_logic_vector(0, 16),
133 => conv_std_logic_vector(0, 16),
134 => conv_std_logic_vector(0, 16),
135 => conv_std_logic_vector(0, 16),
136 => conv_std_logic_vector(0, 16),
137 => conv_std_logic_vector(0, 16),
138 => conv_std_logic_vector(0, 16),
139 => conv_std_logic_vector(0, 16),
140 => conv_std_logic_vector(0, 16),
141 => conv_std_logic_vector(0, 16),
142 => conv_std_logic_vector(0, 16),
143 => conv_std_logic_vector(0, 16),
144 => conv_std_logic_vector(0, 16),
145 => conv_std_logic_vector(0, 16),
146 => conv_std_logic_vector(0, 16),
147 => conv_std_logic_vector(0, 16),
148 => conv_std_logic_vector(0, 16),
149 => conv_std_logic_vector(0, 16),
150 => conv_std_logic_vector(0, 16),
151 => conv_std_logic_vector(0, 16),
152 => conv_std_logic_vector(0, 16),
153 => conv_std_logic_vector(0, 16),
154 => conv_std_logic_vector(0, 16),
155 => conv_std_logic_vector(0, 16),
156 => conv_std_logic_vector(0, 16),
157 => conv_std_logic_vector(0, 16),
158 => conv_std_logic_vector(0, 16),
159 => conv_std_logic_vector(0, 16),
160 => conv_std_logic_vector(0, 16),
161 => conv_std_logic_vector(0, 16),
162 => conv_std_logic_vector(0, 16),
163 => conv_std_logic_vector(0, 16),
164 => conv_std_logic_vector(0, 16),
165 => conv_std_logic_vector(0, 16),
166 => conv_std_logic_vector(0, 16),
167 => conv_std_logic_vector(0, 16),
168 => conv_std_logic_vector(0, 16),
169 => conv_std_logic_vector(0, 16),
170 => conv_std_logic_vector(0, 16),
171 => conv_std_logic_vector(0, 16),
172 => conv_std_logic_vector(0, 16),
173 => conv_std_logic_vector(0, 16),
174 => conv_std_logic_vector(0, 16),
175 => conv_std_logic_vector(0, 16),
176 => conv_std_logic_vector(0, 16),
177 => conv_std_logic_vector(0, 16),
178 => conv_std_logic_vector(0, 16),
179 => conv_std_logic_vector(0, 16),
180 => conv_std_logic_vector(0, 16),
181 => conv_std_logic_vector(0, 16),
182 => conv_std_logic_vector(0, 16),
183 => conv_std_logic_vector(0, 16),
184 => conv_std_logic_vector(0, 16),
185 => conv_std_logic_vector(0, 16),
186 => conv_std_logic_vector(0, 16),
187 => conv_std_logic_vector(0, 16),
188 => conv_std_logic_vector(0, 16),
189 => conv_std_logic_vector(0, 16),
190 => conv_std_logic_vector(0, 16),
191 => conv_std_logic_vector(0, 16),
192 => conv_std_logic_vector(0, 16),
193 => conv_std_logic_vector(0, 16),
194 => conv_std_logic_vector(0, 16),
195 => conv_std_logic_vector(0, 16),
196 => conv_std_logic_vector(0, 16),
197 => conv_std_logic_vector(0, 16),
198 => conv_std_logic_vector(0, 16),
199 => conv_std_logic_vector(0, 16),
200 => conv_std_logic_vector(0, 16),
201 => conv_std_logic_vector(0, 16),
202 => conv_std_logic_vector(0, 16),
203 => conv_std_logic_vector(0, 16),
204 => conv_std_logic_vector(0, 16),
205 => conv_std_logic_vector(0, 16),
206 => conv_std_logic_vector(0, 16),
207 => conv_std_logic_vector(0, 16),
208 => conv_std_logic_vector(0, 16),
209 => conv_std_logic_vector(0, 16),
210 => conv_std_logic_vector(0, 16),
211 => conv_std_logic_vector(0, 16),
212 => conv_std_logic_vector(0, 16),
213 => conv_std_logic_vector(0, 16),
214 => conv_std_logic_vector(0, 16),
215 => conv_std_logic_vector(0, 16),
216 => conv_std_logic_vector(0, 16),
217 => conv_std_logic_vector(0, 16),
218 => conv_std_logic_vector(0, 16),
219 => conv_std_logic_vector(0, 16),
220 => conv_std_logic_vector(0, 16),
221 => conv_std_logic_vector(0, 16),
222 => conv_std_logic_vector(0, 16),
223 => conv_std_logic_vector(0, 16),
224 => conv_std_logic_vector(0, 16),
225 => conv_std_logic_vector(0, 16),
226 => conv_std_logic_vector(0, 16),
227 => conv_std_logic_vector(0, 16),
228 => conv_std_logic_vector(0, 16),
229 => conv_std_logic_vector(0, 16),
230 => conv_std_logic_vector(0, 16),
231 => conv_std_logic_vector(0, 16),
232 => conv_std_logic_vector(0, 16),
233 => conv_std_logic_vector(0, 16),
234 => conv_std_logic_vector(0, 16),
235 => conv_std_logic_vector(0, 16),
236 => conv_std_logic_vector(0, 16),
237 => conv_std_logic_vector(0, 16),
238 => conv_std_logic_vector(0, 16),
239 => conv_std_logic_vector(0, 16),
240 => conv_std_logic_vector(0, 16),
241 => conv_std_logic_vector(0, 16),
242 => conv_std_logic_vector(0, 16),
243 => conv_std_logic_vector(0, 16),
244 => conv_std_logic_vector(0, 16),
245 => conv_std_logic_vector(0, 16),
246 => conv_std_logic_vector(0, 16),
247 => conv_std_logic_vector(0, 16),
248 => conv_std_logic_vector(0, 16),
249 => conv_std_logic_vector(0, 16),
250 => conv_std_logic_vector(0, 16),
251 => conv_std_logic_vector(0, 16),
252 => conv_std_logic_vector(0, 16),
253 => conv_std_logic_vector(0, 16),
254 => conv_std_logic_vector(0, 16),
255 => conv_std_logic_vector(0, 16),
256 => conv_std_logic_vector(0, 16),
257 => conv_std_logic_vector(1, 16),
258 => conv_std_logic_vector(2, 16),
259 => conv_std_logic_vector(3, 16),
260 => conv_std_logic_vector(4, 16),
261 => conv_std_logic_vector(5, 16),
262 => conv_std_logic_vector(6, 16),
263 => conv_std_logic_vector(7, 16),
264 => conv_std_logic_vector(8, 16),
265 => conv_std_logic_vector(9, 16),
266 => conv_std_logic_vector(10, 16),
267 => conv_std_logic_vector(11, 16),
268 => conv_std_logic_vector(12, 16),
269 => conv_std_logic_vector(13, 16),
270 => conv_std_logic_vector(14, 16),
271 => conv_std_logic_vector(15, 16),
272 => conv_std_logic_vector(16, 16),
273 => conv_std_logic_vector(17, 16),
274 => conv_std_logic_vector(18, 16),
275 => conv_std_logic_vector(19, 16),
276 => conv_std_logic_vector(20, 16),
277 => conv_std_logic_vector(21, 16),
278 => conv_std_logic_vector(22, 16),
279 => conv_std_logic_vector(23, 16),
280 => conv_std_logic_vector(24, 16),
281 => conv_std_logic_vector(25, 16),
282 => conv_std_logic_vector(26, 16),
283 => conv_std_logic_vector(27, 16),
284 => conv_std_logic_vector(28, 16),
285 => conv_std_logic_vector(29, 16),
286 => conv_std_logic_vector(30, 16),
287 => conv_std_logic_vector(31, 16),
288 => conv_std_logic_vector(32, 16),
289 => conv_std_logic_vector(33, 16),
290 => conv_std_logic_vector(34, 16),
291 => conv_std_logic_vector(35, 16),
292 => conv_std_logic_vector(36, 16),
293 => conv_std_logic_vector(37, 16),
294 => conv_std_logic_vector(38, 16),
295 => conv_std_logic_vector(39, 16),
296 => conv_std_logic_vector(40, 16),
297 => conv_std_logic_vector(41, 16),
298 => conv_std_logic_vector(42, 16),
299 => conv_std_logic_vector(43, 16),
300 => conv_std_logic_vector(44, 16),
301 => conv_std_logic_vector(45, 16),
302 => conv_std_logic_vector(46, 16),
303 => conv_std_logic_vector(47, 16),
304 => conv_std_logic_vector(48, 16),
305 => conv_std_logic_vector(49, 16),
306 => conv_std_logic_vector(50, 16),
307 => conv_std_logic_vector(51, 16),
308 => conv_std_logic_vector(52, 16),
309 => conv_std_logic_vector(53, 16),
310 => conv_std_logic_vector(54, 16),
311 => conv_std_logic_vector(55, 16),
312 => conv_std_logic_vector(56, 16),
313 => conv_std_logic_vector(57, 16),
314 => conv_std_logic_vector(58, 16),
315 => conv_std_logic_vector(59, 16),
316 => conv_std_logic_vector(60, 16),
317 => conv_std_logic_vector(61, 16),
318 => conv_std_logic_vector(62, 16),
319 => conv_std_logic_vector(63, 16),
320 => conv_std_logic_vector(64, 16),
321 => conv_std_logic_vector(65, 16),
322 => conv_std_logic_vector(66, 16),
323 => conv_std_logic_vector(67, 16),
324 => conv_std_logic_vector(68, 16),
325 => conv_std_logic_vector(69, 16),
326 => conv_std_logic_vector(70, 16),
327 => conv_std_logic_vector(71, 16),
328 => conv_std_logic_vector(72, 16),
329 => conv_std_logic_vector(73, 16),
330 => conv_std_logic_vector(74, 16),
331 => conv_std_logic_vector(75, 16),
332 => conv_std_logic_vector(76, 16),
333 => conv_std_logic_vector(77, 16),
334 => conv_std_logic_vector(78, 16),
335 => conv_std_logic_vector(79, 16),
336 => conv_std_logic_vector(80, 16),
337 => conv_std_logic_vector(81, 16),
338 => conv_std_logic_vector(82, 16),
339 => conv_std_logic_vector(83, 16),
340 => conv_std_logic_vector(84, 16),
341 => conv_std_logic_vector(85, 16),
342 => conv_std_logic_vector(86, 16),
343 => conv_std_logic_vector(87, 16),
344 => conv_std_logic_vector(88, 16),
345 => conv_std_logic_vector(89, 16),
346 => conv_std_logic_vector(90, 16),
347 => conv_std_logic_vector(91, 16),
348 => conv_std_logic_vector(92, 16),
349 => conv_std_logic_vector(93, 16),
350 => conv_std_logic_vector(94, 16),
351 => conv_std_logic_vector(95, 16),
352 => conv_std_logic_vector(96, 16),
353 => conv_std_logic_vector(97, 16),
354 => conv_std_logic_vector(98, 16),
355 => conv_std_logic_vector(99, 16),
356 => conv_std_logic_vector(100, 16),
357 => conv_std_logic_vector(101, 16),
358 => conv_std_logic_vector(102, 16),
359 => conv_std_logic_vector(103, 16),
360 => conv_std_logic_vector(104, 16),
361 => conv_std_logic_vector(105, 16),
362 => conv_std_logic_vector(106, 16),
363 => conv_std_logic_vector(107, 16),
364 => conv_std_logic_vector(108, 16),
365 => conv_std_logic_vector(109, 16),
366 => conv_std_logic_vector(110, 16),
367 => conv_std_logic_vector(111, 16),
368 => conv_std_logic_vector(112, 16),
369 => conv_std_logic_vector(113, 16),
370 => conv_std_logic_vector(114, 16),
371 => conv_std_logic_vector(115, 16),
372 => conv_std_logic_vector(116, 16),
373 => conv_std_logic_vector(117, 16),
374 => conv_std_logic_vector(118, 16),
375 => conv_std_logic_vector(119, 16),
376 => conv_std_logic_vector(120, 16),
377 => conv_std_logic_vector(121, 16),
378 => conv_std_logic_vector(122, 16),
379 => conv_std_logic_vector(123, 16),
380 => conv_std_logic_vector(124, 16),
381 => conv_std_logic_vector(125, 16),
382 => conv_std_logic_vector(126, 16),
383 => conv_std_logic_vector(127, 16),
384 => conv_std_logic_vector(128, 16),
385 => conv_std_logic_vector(129, 16),
386 => conv_std_logic_vector(130, 16),
387 => conv_std_logic_vector(131, 16),
388 => conv_std_logic_vector(132, 16),
389 => conv_std_logic_vector(133, 16),
390 => conv_std_logic_vector(134, 16),
391 => conv_std_logic_vector(135, 16),
392 => conv_std_logic_vector(136, 16),
393 => conv_std_logic_vector(137, 16),
394 => conv_std_logic_vector(138, 16),
395 => conv_std_logic_vector(139, 16),
396 => conv_std_logic_vector(140, 16),
397 => conv_std_logic_vector(141, 16),
398 => conv_std_logic_vector(142, 16),
399 => conv_std_logic_vector(143, 16),
400 => conv_std_logic_vector(144, 16),
401 => conv_std_logic_vector(145, 16),
402 => conv_std_logic_vector(146, 16),
403 => conv_std_logic_vector(147, 16),
404 => conv_std_logic_vector(148, 16),
405 => conv_std_logic_vector(149, 16),
406 => conv_std_logic_vector(150, 16),
407 => conv_std_logic_vector(151, 16),
408 => conv_std_logic_vector(152, 16),
409 => conv_std_logic_vector(153, 16),
410 => conv_std_logic_vector(154, 16),
411 => conv_std_logic_vector(155, 16),
412 => conv_std_logic_vector(156, 16),
413 => conv_std_logic_vector(157, 16),
414 => conv_std_logic_vector(158, 16),
415 => conv_std_logic_vector(159, 16),
416 => conv_std_logic_vector(160, 16),
417 => conv_std_logic_vector(161, 16),
418 => conv_std_logic_vector(162, 16),
419 => conv_std_logic_vector(163, 16),
420 => conv_std_logic_vector(164, 16),
421 => conv_std_logic_vector(165, 16),
422 => conv_std_logic_vector(166, 16),
423 => conv_std_logic_vector(167, 16),
424 => conv_std_logic_vector(168, 16),
425 => conv_std_logic_vector(169, 16),
426 => conv_std_logic_vector(170, 16),
427 => conv_std_logic_vector(171, 16),
428 => conv_std_logic_vector(172, 16),
429 => conv_std_logic_vector(173, 16),
430 => conv_std_logic_vector(174, 16),
431 => conv_std_logic_vector(175, 16),
432 => conv_std_logic_vector(176, 16),
433 => conv_std_logic_vector(177, 16),
434 => conv_std_logic_vector(178, 16),
435 => conv_std_logic_vector(179, 16),
436 => conv_std_logic_vector(180, 16),
437 => conv_std_logic_vector(181, 16),
438 => conv_std_logic_vector(182, 16),
439 => conv_std_logic_vector(183, 16),
440 => conv_std_logic_vector(184, 16),
441 => conv_std_logic_vector(185, 16),
442 => conv_std_logic_vector(186, 16),
443 => conv_std_logic_vector(187, 16),
444 => conv_std_logic_vector(188, 16),
445 => conv_std_logic_vector(189, 16),
446 => conv_std_logic_vector(190, 16),
447 => conv_std_logic_vector(191, 16),
448 => conv_std_logic_vector(192, 16),
449 => conv_std_logic_vector(193, 16),
450 => conv_std_logic_vector(194, 16),
451 => conv_std_logic_vector(195, 16),
452 => conv_std_logic_vector(196, 16),
453 => conv_std_logic_vector(197, 16),
454 => conv_std_logic_vector(198, 16),
455 => conv_std_logic_vector(199, 16),
456 => conv_std_logic_vector(200, 16),
457 => conv_std_logic_vector(201, 16),
458 => conv_std_logic_vector(202, 16),
459 => conv_std_logic_vector(203, 16),
460 => conv_std_logic_vector(204, 16),
461 => conv_std_logic_vector(205, 16),
462 => conv_std_logic_vector(206, 16),
463 => conv_std_logic_vector(207, 16),
464 => conv_std_logic_vector(208, 16),
465 => conv_std_logic_vector(209, 16),
466 => conv_std_logic_vector(210, 16),
467 => conv_std_logic_vector(211, 16),
468 => conv_std_logic_vector(212, 16),
469 => conv_std_logic_vector(213, 16),
470 => conv_std_logic_vector(214, 16),
471 => conv_std_logic_vector(215, 16),
472 => conv_std_logic_vector(216, 16),
473 => conv_std_logic_vector(217, 16),
474 => conv_std_logic_vector(218, 16),
475 => conv_std_logic_vector(219, 16),
476 => conv_std_logic_vector(220, 16),
477 => conv_std_logic_vector(221, 16),
478 => conv_std_logic_vector(222, 16),
479 => conv_std_logic_vector(223, 16),
480 => conv_std_logic_vector(224, 16),
481 => conv_std_logic_vector(225, 16),
482 => conv_std_logic_vector(226, 16),
483 => conv_std_logic_vector(227, 16),
484 => conv_std_logic_vector(228, 16),
485 => conv_std_logic_vector(229, 16),
486 => conv_std_logic_vector(230, 16),
487 => conv_std_logic_vector(231, 16),
488 => conv_std_logic_vector(232, 16),
489 => conv_std_logic_vector(233, 16),
490 => conv_std_logic_vector(234, 16),
491 => conv_std_logic_vector(235, 16),
492 => conv_std_logic_vector(236, 16),
493 => conv_std_logic_vector(237, 16),
494 => conv_std_logic_vector(238, 16),
495 => conv_std_logic_vector(239, 16),
496 => conv_std_logic_vector(240, 16),
497 => conv_std_logic_vector(241, 16),
498 => conv_std_logic_vector(242, 16),
499 => conv_std_logic_vector(243, 16),
500 => conv_std_logic_vector(244, 16),
501 => conv_std_logic_vector(245, 16),
502 => conv_std_logic_vector(246, 16),
503 => conv_std_logic_vector(247, 16),
504 => conv_std_logic_vector(248, 16),
505 => conv_std_logic_vector(249, 16),
506 => conv_std_logic_vector(250, 16),
507 => conv_std_logic_vector(251, 16),
508 => conv_std_logic_vector(252, 16),
509 => conv_std_logic_vector(253, 16),
510 => conv_std_logic_vector(254, 16),
511 => conv_std_logic_vector(255, 16),
512 => conv_std_logic_vector(0, 16),
513 => conv_std_logic_vector(2, 16),
514 => conv_std_logic_vector(4, 16),
515 => conv_std_logic_vector(6, 16),
516 => conv_std_logic_vector(8, 16),
517 => conv_std_logic_vector(10, 16),
518 => conv_std_logic_vector(12, 16),
519 => conv_std_logic_vector(14, 16),
520 => conv_std_logic_vector(16, 16),
521 => conv_std_logic_vector(18, 16),
522 => conv_std_logic_vector(20, 16),
523 => conv_std_logic_vector(22, 16),
524 => conv_std_logic_vector(24, 16),
525 => conv_std_logic_vector(26, 16),
526 => conv_std_logic_vector(28, 16),
527 => conv_std_logic_vector(30, 16),
528 => conv_std_logic_vector(32, 16),
529 => conv_std_logic_vector(34, 16),
530 => conv_std_logic_vector(36, 16),
531 => conv_std_logic_vector(38, 16),
532 => conv_std_logic_vector(40, 16),
533 => conv_std_logic_vector(42, 16),
534 => conv_std_logic_vector(44, 16),
535 => conv_std_logic_vector(46, 16),
536 => conv_std_logic_vector(48, 16),
537 => conv_std_logic_vector(50, 16),
538 => conv_std_logic_vector(52, 16),
539 => conv_std_logic_vector(54, 16),
540 => conv_std_logic_vector(56, 16),
541 => conv_std_logic_vector(58, 16),
542 => conv_std_logic_vector(60, 16),
543 => conv_std_logic_vector(62, 16),
544 => conv_std_logic_vector(64, 16),
545 => conv_std_logic_vector(66, 16),
546 => conv_std_logic_vector(68, 16),
547 => conv_std_logic_vector(70, 16),
548 => conv_std_logic_vector(72, 16),
549 => conv_std_logic_vector(74, 16),
550 => conv_std_logic_vector(76, 16),
551 => conv_std_logic_vector(78, 16),
552 => conv_std_logic_vector(80, 16),
553 => conv_std_logic_vector(82, 16),
554 => conv_std_logic_vector(84, 16),
555 => conv_std_logic_vector(86, 16),
556 => conv_std_logic_vector(88, 16),
557 => conv_std_logic_vector(90, 16),
558 => conv_std_logic_vector(92, 16),
559 => conv_std_logic_vector(94, 16),
560 => conv_std_logic_vector(96, 16),
561 => conv_std_logic_vector(98, 16),
562 => conv_std_logic_vector(100, 16),
563 => conv_std_logic_vector(102, 16),
564 => conv_std_logic_vector(104, 16),
565 => conv_std_logic_vector(106, 16),
566 => conv_std_logic_vector(108, 16),
567 => conv_std_logic_vector(110, 16),
568 => conv_std_logic_vector(112, 16),
569 => conv_std_logic_vector(114, 16),
570 => conv_std_logic_vector(116, 16),
571 => conv_std_logic_vector(118, 16),
572 => conv_std_logic_vector(120, 16),
573 => conv_std_logic_vector(122, 16),
574 => conv_std_logic_vector(124, 16),
575 => conv_std_logic_vector(126, 16),
576 => conv_std_logic_vector(128, 16),
577 => conv_std_logic_vector(130, 16),
578 => conv_std_logic_vector(132, 16),
579 => conv_std_logic_vector(134, 16),
580 => conv_std_logic_vector(136, 16),
581 => conv_std_logic_vector(138, 16),
582 => conv_std_logic_vector(140, 16),
583 => conv_std_logic_vector(142, 16),
584 => conv_std_logic_vector(144, 16),
585 => conv_std_logic_vector(146, 16),
586 => conv_std_logic_vector(148, 16),
587 => conv_std_logic_vector(150, 16),
588 => conv_std_logic_vector(152, 16),
589 => conv_std_logic_vector(154, 16),
590 => conv_std_logic_vector(156, 16),
591 => conv_std_logic_vector(158, 16),
592 => conv_std_logic_vector(160, 16),
593 => conv_std_logic_vector(162, 16),
594 => conv_std_logic_vector(164, 16),
595 => conv_std_logic_vector(166, 16),
596 => conv_std_logic_vector(168, 16),
597 => conv_std_logic_vector(170, 16),
598 => conv_std_logic_vector(172, 16),
599 => conv_std_logic_vector(174, 16),
600 => conv_std_logic_vector(176, 16),
601 => conv_std_logic_vector(178, 16),
602 => conv_std_logic_vector(180, 16),
603 => conv_std_logic_vector(182, 16),
604 => conv_std_logic_vector(184, 16),
605 => conv_std_logic_vector(186, 16),
606 => conv_std_logic_vector(188, 16),
607 => conv_std_logic_vector(190, 16),
608 => conv_std_logic_vector(192, 16),
609 => conv_std_logic_vector(194, 16),
610 => conv_std_logic_vector(196, 16),
611 => conv_std_logic_vector(198, 16),
612 => conv_std_logic_vector(200, 16),
613 => conv_std_logic_vector(202, 16),
614 => conv_std_logic_vector(204, 16),
615 => conv_std_logic_vector(206, 16),
616 => conv_std_logic_vector(208, 16),
617 => conv_std_logic_vector(210, 16),
618 => conv_std_logic_vector(212, 16),
619 => conv_std_logic_vector(214, 16),
620 => conv_std_logic_vector(216, 16),
621 => conv_std_logic_vector(218, 16),
622 => conv_std_logic_vector(220, 16),
623 => conv_std_logic_vector(222, 16),
624 => conv_std_logic_vector(224, 16),
625 => conv_std_logic_vector(226, 16),
626 => conv_std_logic_vector(228, 16),
627 => conv_std_logic_vector(230, 16),
628 => conv_std_logic_vector(232, 16),
629 => conv_std_logic_vector(234, 16),
630 => conv_std_logic_vector(236, 16),
631 => conv_std_logic_vector(238, 16),
632 => conv_std_logic_vector(240, 16),
633 => conv_std_logic_vector(242, 16),
634 => conv_std_logic_vector(244, 16),
635 => conv_std_logic_vector(246, 16),
636 => conv_std_logic_vector(248, 16),
637 => conv_std_logic_vector(250, 16),
638 => conv_std_logic_vector(252, 16),
639 => conv_std_logic_vector(254, 16),
640 => conv_std_logic_vector(256, 16),
641 => conv_std_logic_vector(258, 16),
642 => conv_std_logic_vector(260, 16),
643 => conv_std_logic_vector(262, 16),
644 => conv_std_logic_vector(264, 16),
645 => conv_std_logic_vector(266, 16),
646 => conv_std_logic_vector(268, 16),
647 => conv_std_logic_vector(270, 16),
648 => conv_std_logic_vector(272, 16),
649 => conv_std_logic_vector(274, 16),
650 => conv_std_logic_vector(276, 16),
651 => conv_std_logic_vector(278, 16),
652 => conv_std_logic_vector(280, 16),
653 => conv_std_logic_vector(282, 16),
654 => conv_std_logic_vector(284, 16),
655 => conv_std_logic_vector(286, 16),
656 => conv_std_logic_vector(288, 16),
657 => conv_std_logic_vector(290, 16),
658 => conv_std_logic_vector(292, 16),
659 => conv_std_logic_vector(294, 16),
660 => conv_std_logic_vector(296, 16),
661 => conv_std_logic_vector(298, 16),
662 => conv_std_logic_vector(300, 16),
663 => conv_std_logic_vector(302, 16),
664 => conv_std_logic_vector(304, 16),
665 => conv_std_logic_vector(306, 16),
666 => conv_std_logic_vector(308, 16),
667 => conv_std_logic_vector(310, 16),
668 => conv_std_logic_vector(312, 16),
669 => conv_std_logic_vector(314, 16),
670 => conv_std_logic_vector(316, 16),
671 => conv_std_logic_vector(318, 16),
672 => conv_std_logic_vector(320, 16),
673 => conv_std_logic_vector(322, 16),
674 => conv_std_logic_vector(324, 16),
675 => conv_std_logic_vector(326, 16),
676 => conv_std_logic_vector(328, 16),
677 => conv_std_logic_vector(330, 16),
678 => conv_std_logic_vector(332, 16),
679 => conv_std_logic_vector(334, 16),
680 => conv_std_logic_vector(336, 16),
681 => conv_std_logic_vector(338, 16),
682 => conv_std_logic_vector(340, 16),
683 => conv_std_logic_vector(342, 16),
684 => conv_std_logic_vector(344, 16),
685 => conv_std_logic_vector(346, 16),
686 => conv_std_logic_vector(348, 16),
687 => conv_std_logic_vector(350, 16),
688 => conv_std_logic_vector(352, 16),
689 => conv_std_logic_vector(354, 16),
690 => conv_std_logic_vector(356, 16),
691 => conv_std_logic_vector(358, 16),
692 => conv_std_logic_vector(360, 16),
693 => conv_std_logic_vector(362, 16),
694 => conv_std_logic_vector(364, 16),
695 => conv_std_logic_vector(366, 16),
696 => conv_std_logic_vector(368, 16),
697 => conv_std_logic_vector(370, 16),
698 => conv_std_logic_vector(372, 16),
699 => conv_std_logic_vector(374, 16),
700 => conv_std_logic_vector(376, 16),
701 => conv_std_logic_vector(378, 16),
702 => conv_std_logic_vector(380, 16),
703 => conv_std_logic_vector(382, 16),
704 => conv_std_logic_vector(384, 16),
705 => conv_std_logic_vector(386, 16),
706 => conv_std_logic_vector(388, 16),
707 => conv_std_logic_vector(390, 16),
708 => conv_std_logic_vector(392, 16),
709 => conv_std_logic_vector(394, 16),
710 => conv_std_logic_vector(396, 16),
711 => conv_std_logic_vector(398, 16),
712 => conv_std_logic_vector(400, 16),
713 => conv_std_logic_vector(402, 16),
714 => conv_std_logic_vector(404, 16),
715 => conv_std_logic_vector(406, 16),
716 => conv_std_logic_vector(408, 16),
717 => conv_std_logic_vector(410, 16),
718 => conv_std_logic_vector(412, 16),
719 => conv_std_logic_vector(414, 16),
720 => conv_std_logic_vector(416, 16),
721 => conv_std_logic_vector(418, 16),
722 => conv_std_logic_vector(420, 16),
723 => conv_std_logic_vector(422, 16),
724 => conv_std_logic_vector(424, 16),
725 => conv_std_logic_vector(426, 16),
726 => conv_std_logic_vector(428, 16),
727 => conv_std_logic_vector(430, 16),
728 => conv_std_logic_vector(432, 16),
729 => conv_std_logic_vector(434, 16),
730 => conv_std_logic_vector(436, 16),
731 => conv_std_logic_vector(438, 16),
732 => conv_std_logic_vector(440, 16),
733 => conv_std_logic_vector(442, 16),
734 => conv_std_logic_vector(444, 16),
735 => conv_std_logic_vector(446, 16),
736 => conv_std_logic_vector(448, 16),
737 => conv_std_logic_vector(450, 16),
738 => conv_std_logic_vector(452, 16),
739 => conv_std_logic_vector(454, 16),
740 => conv_std_logic_vector(456, 16),
741 => conv_std_logic_vector(458, 16),
742 => conv_std_logic_vector(460, 16),
743 => conv_std_logic_vector(462, 16),
744 => conv_std_logic_vector(464, 16),
745 => conv_std_logic_vector(466, 16),
746 => conv_std_logic_vector(468, 16),
747 => conv_std_logic_vector(470, 16),
748 => conv_std_logic_vector(472, 16),
749 => conv_std_logic_vector(474, 16),
750 => conv_std_logic_vector(476, 16),
751 => conv_std_logic_vector(478, 16),
752 => conv_std_logic_vector(480, 16),
753 => conv_std_logic_vector(482, 16),
754 => conv_std_logic_vector(484, 16),
755 => conv_std_logic_vector(486, 16),
756 => conv_std_logic_vector(488, 16),
757 => conv_std_logic_vector(490, 16),
758 => conv_std_logic_vector(492, 16),
759 => conv_std_logic_vector(494, 16),
760 => conv_std_logic_vector(496, 16),
761 => conv_std_logic_vector(498, 16),
762 => conv_std_logic_vector(500, 16),
763 => conv_std_logic_vector(502, 16),
764 => conv_std_logic_vector(504, 16),
765 => conv_std_logic_vector(506, 16),
766 => conv_std_logic_vector(508, 16),
767 => conv_std_logic_vector(510, 16),
768 => conv_std_logic_vector(0, 16),
769 => conv_std_logic_vector(3, 16),
770 => conv_std_logic_vector(6, 16),
771 => conv_std_logic_vector(9, 16),
772 => conv_std_logic_vector(12, 16),
773 => conv_std_logic_vector(15, 16),
774 => conv_std_logic_vector(18, 16),
775 => conv_std_logic_vector(21, 16),
776 => conv_std_logic_vector(24, 16),
777 => conv_std_logic_vector(27, 16),
778 => conv_std_logic_vector(30, 16),
779 => conv_std_logic_vector(33, 16),
780 => conv_std_logic_vector(36, 16),
781 => conv_std_logic_vector(39, 16),
782 => conv_std_logic_vector(42, 16),
783 => conv_std_logic_vector(45, 16),
784 => conv_std_logic_vector(48, 16),
785 => conv_std_logic_vector(51, 16),
786 => conv_std_logic_vector(54, 16),
787 => conv_std_logic_vector(57, 16),
788 => conv_std_logic_vector(60, 16),
789 => conv_std_logic_vector(63, 16),
790 => conv_std_logic_vector(66, 16),
791 => conv_std_logic_vector(69, 16),
792 => conv_std_logic_vector(72, 16),
793 => conv_std_logic_vector(75, 16),
794 => conv_std_logic_vector(78, 16),
795 => conv_std_logic_vector(81, 16),
796 => conv_std_logic_vector(84, 16),
797 => conv_std_logic_vector(87, 16),
798 => conv_std_logic_vector(90, 16),
799 => conv_std_logic_vector(93, 16),
800 => conv_std_logic_vector(96, 16),
801 => conv_std_logic_vector(99, 16),
802 => conv_std_logic_vector(102, 16),
803 => conv_std_logic_vector(105, 16),
804 => conv_std_logic_vector(108, 16),
805 => conv_std_logic_vector(111, 16),
806 => conv_std_logic_vector(114, 16),
807 => conv_std_logic_vector(117, 16),
808 => conv_std_logic_vector(120, 16),
809 => conv_std_logic_vector(123, 16),
810 => conv_std_logic_vector(126, 16),
811 => conv_std_logic_vector(129, 16),
812 => conv_std_logic_vector(132, 16),
813 => conv_std_logic_vector(135, 16),
814 => conv_std_logic_vector(138, 16),
815 => conv_std_logic_vector(141, 16),
816 => conv_std_logic_vector(144, 16),
817 => conv_std_logic_vector(147, 16),
818 => conv_std_logic_vector(150, 16),
819 => conv_std_logic_vector(153, 16),
820 => conv_std_logic_vector(156, 16),
821 => conv_std_logic_vector(159, 16),
822 => conv_std_logic_vector(162, 16),
823 => conv_std_logic_vector(165, 16),
824 => conv_std_logic_vector(168, 16),
825 => conv_std_logic_vector(171, 16),
826 => conv_std_logic_vector(174, 16),
827 => conv_std_logic_vector(177, 16),
828 => conv_std_logic_vector(180, 16),
829 => conv_std_logic_vector(183, 16),
830 => conv_std_logic_vector(186, 16),
831 => conv_std_logic_vector(189, 16),
832 => conv_std_logic_vector(192, 16),
833 => conv_std_logic_vector(195, 16),
834 => conv_std_logic_vector(198, 16),
835 => conv_std_logic_vector(201, 16),
836 => conv_std_logic_vector(204, 16),
837 => conv_std_logic_vector(207, 16),
838 => conv_std_logic_vector(210, 16),
839 => conv_std_logic_vector(213, 16),
840 => conv_std_logic_vector(216, 16),
841 => conv_std_logic_vector(219, 16),
842 => conv_std_logic_vector(222, 16),
843 => conv_std_logic_vector(225, 16),
844 => conv_std_logic_vector(228, 16),
845 => conv_std_logic_vector(231, 16),
846 => conv_std_logic_vector(234, 16),
847 => conv_std_logic_vector(237, 16),
848 => conv_std_logic_vector(240, 16),
849 => conv_std_logic_vector(243, 16),
850 => conv_std_logic_vector(246, 16),
851 => conv_std_logic_vector(249, 16),
852 => conv_std_logic_vector(252, 16),
853 => conv_std_logic_vector(255, 16),
854 => conv_std_logic_vector(258, 16),
855 => conv_std_logic_vector(261, 16),
856 => conv_std_logic_vector(264, 16),
857 => conv_std_logic_vector(267, 16),
858 => conv_std_logic_vector(270, 16),
859 => conv_std_logic_vector(273, 16),
860 => conv_std_logic_vector(276, 16),
861 => conv_std_logic_vector(279, 16),
862 => conv_std_logic_vector(282, 16),
863 => conv_std_logic_vector(285, 16),
864 => conv_std_logic_vector(288, 16),
865 => conv_std_logic_vector(291, 16),
866 => conv_std_logic_vector(294, 16),
867 => conv_std_logic_vector(297, 16),
868 => conv_std_logic_vector(300, 16),
869 => conv_std_logic_vector(303, 16),
870 => conv_std_logic_vector(306, 16),
871 => conv_std_logic_vector(309, 16),
872 => conv_std_logic_vector(312, 16),
873 => conv_std_logic_vector(315, 16),
874 => conv_std_logic_vector(318, 16),
875 => conv_std_logic_vector(321, 16),
876 => conv_std_logic_vector(324, 16),
877 => conv_std_logic_vector(327, 16),
878 => conv_std_logic_vector(330, 16),
879 => conv_std_logic_vector(333, 16),
880 => conv_std_logic_vector(336, 16),
881 => conv_std_logic_vector(339, 16),
882 => conv_std_logic_vector(342, 16),
883 => conv_std_logic_vector(345, 16),
884 => conv_std_logic_vector(348, 16),
885 => conv_std_logic_vector(351, 16),
886 => conv_std_logic_vector(354, 16),
887 => conv_std_logic_vector(357, 16),
888 => conv_std_logic_vector(360, 16),
889 => conv_std_logic_vector(363, 16),
890 => conv_std_logic_vector(366, 16),
891 => conv_std_logic_vector(369, 16),
892 => conv_std_logic_vector(372, 16),
893 => conv_std_logic_vector(375, 16),
894 => conv_std_logic_vector(378, 16),
895 => conv_std_logic_vector(381, 16),
896 => conv_std_logic_vector(384, 16),
897 => conv_std_logic_vector(387, 16),
898 => conv_std_logic_vector(390, 16),
899 => conv_std_logic_vector(393, 16),
900 => conv_std_logic_vector(396, 16),
901 => conv_std_logic_vector(399, 16),
902 => conv_std_logic_vector(402, 16),
903 => conv_std_logic_vector(405, 16),
904 => conv_std_logic_vector(408, 16),
905 => conv_std_logic_vector(411, 16),
906 => conv_std_logic_vector(414, 16),
907 => conv_std_logic_vector(417, 16),
908 => conv_std_logic_vector(420, 16),
909 => conv_std_logic_vector(423, 16),
910 => conv_std_logic_vector(426, 16),
911 => conv_std_logic_vector(429, 16),
912 => conv_std_logic_vector(432, 16),
913 => conv_std_logic_vector(435, 16),
914 => conv_std_logic_vector(438, 16),
915 => conv_std_logic_vector(441, 16),
916 => conv_std_logic_vector(444, 16),
917 => conv_std_logic_vector(447, 16),
918 => conv_std_logic_vector(450, 16),
919 => conv_std_logic_vector(453, 16),
920 => conv_std_logic_vector(456, 16),
921 => conv_std_logic_vector(459, 16),
922 => conv_std_logic_vector(462, 16),
923 => conv_std_logic_vector(465, 16),
924 => conv_std_logic_vector(468, 16),
925 => conv_std_logic_vector(471, 16),
926 => conv_std_logic_vector(474, 16),
927 => conv_std_logic_vector(477, 16),
928 => conv_std_logic_vector(480, 16),
929 => conv_std_logic_vector(483, 16),
930 => conv_std_logic_vector(486, 16),
931 => conv_std_logic_vector(489, 16),
932 => conv_std_logic_vector(492, 16),
933 => conv_std_logic_vector(495, 16),
934 => conv_std_logic_vector(498, 16),
935 => conv_std_logic_vector(501, 16),
936 => conv_std_logic_vector(504, 16),
937 => conv_std_logic_vector(507, 16),
938 => conv_std_logic_vector(510, 16),
939 => conv_std_logic_vector(513, 16),
940 => conv_std_logic_vector(516, 16),
941 => conv_std_logic_vector(519, 16),
942 => conv_std_logic_vector(522, 16),
943 => conv_std_logic_vector(525, 16),
944 => conv_std_logic_vector(528, 16),
945 => conv_std_logic_vector(531, 16),
946 => conv_std_logic_vector(534, 16),
947 => conv_std_logic_vector(537, 16),
948 => conv_std_logic_vector(540, 16),
949 => conv_std_logic_vector(543, 16),
950 => conv_std_logic_vector(546, 16),
951 => conv_std_logic_vector(549, 16),
952 => conv_std_logic_vector(552, 16),
953 => conv_std_logic_vector(555, 16),
954 => conv_std_logic_vector(558, 16),
955 => conv_std_logic_vector(561, 16),
956 => conv_std_logic_vector(564, 16),
957 => conv_std_logic_vector(567, 16),
958 => conv_std_logic_vector(570, 16),
959 => conv_std_logic_vector(573, 16),
960 => conv_std_logic_vector(576, 16),
961 => conv_std_logic_vector(579, 16),
962 => conv_std_logic_vector(582, 16),
963 => conv_std_logic_vector(585, 16),
964 => conv_std_logic_vector(588, 16),
965 => conv_std_logic_vector(591, 16),
966 => conv_std_logic_vector(594, 16),
967 => conv_std_logic_vector(597, 16),
968 => conv_std_logic_vector(600, 16),
969 => conv_std_logic_vector(603, 16),
970 => conv_std_logic_vector(606, 16),
971 => conv_std_logic_vector(609, 16),
972 => conv_std_logic_vector(612, 16),
973 => conv_std_logic_vector(615, 16),
974 => conv_std_logic_vector(618, 16),
975 => conv_std_logic_vector(621, 16),
976 => conv_std_logic_vector(624, 16),
977 => conv_std_logic_vector(627, 16),
978 => conv_std_logic_vector(630, 16),
979 => conv_std_logic_vector(633, 16),
980 => conv_std_logic_vector(636, 16),
981 => conv_std_logic_vector(639, 16),
982 => conv_std_logic_vector(642, 16),
983 => conv_std_logic_vector(645, 16),
984 => conv_std_logic_vector(648, 16),
985 => conv_std_logic_vector(651, 16),
986 => conv_std_logic_vector(654, 16),
987 => conv_std_logic_vector(657, 16),
988 => conv_std_logic_vector(660, 16),
989 => conv_std_logic_vector(663, 16),
990 => conv_std_logic_vector(666, 16),
991 => conv_std_logic_vector(669, 16),
992 => conv_std_logic_vector(672, 16),
993 => conv_std_logic_vector(675, 16),
994 => conv_std_logic_vector(678, 16),
995 => conv_std_logic_vector(681, 16),
996 => conv_std_logic_vector(684, 16),
997 => conv_std_logic_vector(687, 16),
998 => conv_std_logic_vector(690, 16),
999 => conv_std_logic_vector(693, 16),
1000 => conv_std_logic_vector(696, 16),
1001 => conv_std_logic_vector(699, 16),
1002 => conv_std_logic_vector(702, 16),
1003 => conv_std_logic_vector(705, 16),
1004 => conv_std_logic_vector(708, 16),
1005 => conv_std_logic_vector(711, 16),
1006 => conv_std_logic_vector(714, 16),
1007 => conv_std_logic_vector(717, 16),
1008 => conv_std_logic_vector(720, 16),
1009 => conv_std_logic_vector(723, 16),
1010 => conv_std_logic_vector(726, 16),
1011 => conv_std_logic_vector(729, 16),
1012 => conv_std_logic_vector(732, 16),
1013 => conv_std_logic_vector(735, 16),
1014 => conv_std_logic_vector(738, 16),
1015 => conv_std_logic_vector(741, 16),
1016 => conv_std_logic_vector(744, 16),
1017 => conv_std_logic_vector(747, 16),
1018 => conv_std_logic_vector(750, 16),
1019 => conv_std_logic_vector(753, 16),
1020 => conv_std_logic_vector(756, 16),
1021 => conv_std_logic_vector(759, 16),
1022 => conv_std_logic_vector(762, 16),
1023 => conv_std_logic_vector(765, 16),
1024 => conv_std_logic_vector(0, 16),
1025 => conv_std_logic_vector(4, 16),
1026 => conv_std_logic_vector(8, 16),
1027 => conv_std_logic_vector(12, 16),
1028 => conv_std_logic_vector(16, 16),
1029 => conv_std_logic_vector(20, 16),
1030 => conv_std_logic_vector(24, 16),
1031 => conv_std_logic_vector(28, 16),
1032 => conv_std_logic_vector(32, 16),
1033 => conv_std_logic_vector(36, 16),
1034 => conv_std_logic_vector(40, 16),
1035 => conv_std_logic_vector(44, 16),
1036 => conv_std_logic_vector(48, 16),
1037 => conv_std_logic_vector(52, 16),
1038 => conv_std_logic_vector(56, 16),
1039 => conv_std_logic_vector(60, 16),
1040 => conv_std_logic_vector(64, 16),
1041 => conv_std_logic_vector(68, 16),
1042 => conv_std_logic_vector(72, 16),
1043 => conv_std_logic_vector(76, 16),
1044 => conv_std_logic_vector(80, 16),
1045 => conv_std_logic_vector(84, 16),
1046 => conv_std_logic_vector(88, 16),
1047 => conv_std_logic_vector(92, 16),
1048 => conv_std_logic_vector(96, 16),
1049 => conv_std_logic_vector(100, 16),
1050 => conv_std_logic_vector(104, 16),
1051 => conv_std_logic_vector(108, 16),
1052 => conv_std_logic_vector(112, 16),
1053 => conv_std_logic_vector(116, 16),
1054 => conv_std_logic_vector(120, 16),
1055 => conv_std_logic_vector(124, 16),
1056 => conv_std_logic_vector(128, 16),
1057 => conv_std_logic_vector(132, 16),
1058 => conv_std_logic_vector(136, 16),
1059 => conv_std_logic_vector(140, 16),
1060 => conv_std_logic_vector(144, 16),
1061 => conv_std_logic_vector(148, 16),
1062 => conv_std_logic_vector(152, 16),
1063 => conv_std_logic_vector(156, 16),
1064 => conv_std_logic_vector(160, 16),
1065 => conv_std_logic_vector(164, 16),
1066 => conv_std_logic_vector(168, 16),
1067 => conv_std_logic_vector(172, 16),
1068 => conv_std_logic_vector(176, 16),
1069 => conv_std_logic_vector(180, 16),
1070 => conv_std_logic_vector(184, 16),
1071 => conv_std_logic_vector(188, 16),
1072 => conv_std_logic_vector(192, 16),
1073 => conv_std_logic_vector(196, 16),
1074 => conv_std_logic_vector(200, 16),
1075 => conv_std_logic_vector(204, 16),
1076 => conv_std_logic_vector(208, 16),
1077 => conv_std_logic_vector(212, 16),
1078 => conv_std_logic_vector(216, 16),
1079 => conv_std_logic_vector(220, 16),
1080 => conv_std_logic_vector(224, 16),
1081 => conv_std_logic_vector(228, 16),
1082 => conv_std_logic_vector(232, 16),
1083 => conv_std_logic_vector(236, 16),
1084 => conv_std_logic_vector(240, 16),
1085 => conv_std_logic_vector(244, 16),
1086 => conv_std_logic_vector(248, 16),
1087 => conv_std_logic_vector(252, 16),
1088 => conv_std_logic_vector(256, 16),
1089 => conv_std_logic_vector(260, 16),
1090 => conv_std_logic_vector(264, 16),
1091 => conv_std_logic_vector(268, 16),
1092 => conv_std_logic_vector(272, 16),
1093 => conv_std_logic_vector(276, 16),
1094 => conv_std_logic_vector(280, 16),
1095 => conv_std_logic_vector(284, 16),
1096 => conv_std_logic_vector(288, 16),
1097 => conv_std_logic_vector(292, 16),
1098 => conv_std_logic_vector(296, 16),
1099 => conv_std_logic_vector(300, 16),
1100 => conv_std_logic_vector(304, 16),
1101 => conv_std_logic_vector(308, 16),
1102 => conv_std_logic_vector(312, 16),
1103 => conv_std_logic_vector(316, 16),
1104 => conv_std_logic_vector(320, 16),
1105 => conv_std_logic_vector(324, 16),
1106 => conv_std_logic_vector(328, 16),
1107 => conv_std_logic_vector(332, 16),
1108 => conv_std_logic_vector(336, 16),
1109 => conv_std_logic_vector(340, 16),
1110 => conv_std_logic_vector(344, 16),
1111 => conv_std_logic_vector(348, 16),
1112 => conv_std_logic_vector(352, 16),
1113 => conv_std_logic_vector(356, 16),
1114 => conv_std_logic_vector(360, 16),
1115 => conv_std_logic_vector(364, 16),
1116 => conv_std_logic_vector(368, 16),
1117 => conv_std_logic_vector(372, 16),
1118 => conv_std_logic_vector(376, 16),
1119 => conv_std_logic_vector(380, 16),
1120 => conv_std_logic_vector(384, 16),
1121 => conv_std_logic_vector(388, 16),
1122 => conv_std_logic_vector(392, 16),
1123 => conv_std_logic_vector(396, 16),
1124 => conv_std_logic_vector(400, 16),
1125 => conv_std_logic_vector(404, 16),
1126 => conv_std_logic_vector(408, 16),
1127 => conv_std_logic_vector(412, 16),
1128 => conv_std_logic_vector(416, 16),
1129 => conv_std_logic_vector(420, 16),
1130 => conv_std_logic_vector(424, 16),
1131 => conv_std_logic_vector(428, 16),
1132 => conv_std_logic_vector(432, 16),
1133 => conv_std_logic_vector(436, 16),
1134 => conv_std_logic_vector(440, 16),
1135 => conv_std_logic_vector(444, 16),
1136 => conv_std_logic_vector(448, 16),
1137 => conv_std_logic_vector(452, 16),
1138 => conv_std_logic_vector(456, 16),
1139 => conv_std_logic_vector(460, 16),
1140 => conv_std_logic_vector(464, 16),
1141 => conv_std_logic_vector(468, 16),
1142 => conv_std_logic_vector(472, 16),
1143 => conv_std_logic_vector(476, 16),
1144 => conv_std_logic_vector(480, 16),
1145 => conv_std_logic_vector(484, 16),
1146 => conv_std_logic_vector(488, 16),
1147 => conv_std_logic_vector(492, 16),
1148 => conv_std_logic_vector(496, 16),
1149 => conv_std_logic_vector(500, 16),
1150 => conv_std_logic_vector(504, 16),
1151 => conv_std_logic_vector(508, 16),
1152 => conv_std_logic_vector(512, 16),
1153 => conv_std_logic_vector(516, 16),
1154 => conv_std_logic_vector(520, 16),
1155 => conv_std_logic_vector(524, 16),
1156 => conv_std_logic_vector(528, 16),
1157 => conv_std_logic_vector(532, 16),
1158 => conv_std_logic_vector(536, 16),
1159 => conv_std_logic_vector(540, 16),
1160 => conv_std_logic_vector(544, 16),
1161 => conv_std_logic_vector(548, 16),
1162 => conv_std_logic_vector(552, 16),
1163 => conv_std_logic_vector(556, 16),
1164 => conv_std_logic_vector(560, 16),
1165 => conv_std_logic_vector(564, 16),
1166 => conv_std_logic_vector(568, 16),
1167 => conv_std_logic_vector(572, 16),
1168 => conv_std_logic_vector(576, 16),
1169 => conv_std_logic_vector(580, 16),
1170 => conv_std_logic_vector(584, 16),
1171 => conv_std_logic_vector(588, 16),
1172 => conv_std_logic_vector(592, 16),
1173 => conv_std_logic_vector(596, 16),
1174 => conv_std_logic_vector(600, 16),
1175 => conv_std_logic_vector(604, 16),
1176 => conv_std_logic_vector(608, 16),
1177 => conv_std_logic_vector(612, 16),
1178 => conv_std_logic_vector(616, 16),
1179 => conv_std_logic_vector(620, 16),
1180 => conv_std_logic_vector(624, 16),
1181 => conv_std_logic_vector(628, 16),
1182 => conv_std_logic_vector(632, 16),
1183 => conv_std_logic_vector(636, 16),
1184 => conv_std_logic_vector(640, 16),
1185 => conv_std_logic_vector(644, 16),
1186 => conv_std_logic_vector(648, 16),
1187 => conv_std_logic_vector(652, 16),
1188 => conv_std_logic_vector(656, 16),
1189 => conv_std_logic_vector(660, 16),
1190 => conv_std_logic_vector(664, 16),
1191 => conv_std_logic_vector(668, 16),
1192 => conv_std_logic_vector(672, 16),
1193 => conv_std_logic_vector(676, 16),
1194 => conv_std_logic_vector(680, 16),
1195 => conv_std_logic_vector(684, 16),
1196 => conv_std_logic_vector(688, 16),
1197 => conv_std_logic_vector(692, 16),
1198 => conv_std_logic_vector(696, 16),
1199 => conv_std_logic_vector(700, 16),
1200 => conv_std_logic_vector(704, 16),
1201 => conv_std_logic_vector(708, 16),
1202 => conv_std_logic_vector(712, 16),
1203 => conv_std_logic_vector(716, 16),
1204 => conv_std_logic_vector(720, 16),
1205 => conv_std_logic_vector(724, 16),
1206 => conv_std_logic_vector(728, 16),
1207 => conv_std_logic_vector(732, 16),
1208 => conv_std_logic_vector(736, 16),
1209 => conv_std_logic_vector(740, 16),
1210 => conv_std_logic_vector(744, 16),
1211 => conv_std_logic_vector(748, 16),
1212 => conv_std_logic_vector(752, 16),
1213 => conv_std_logic_vector(756, 16),
1214 => conv_std_logic_vector(760, 16),
1215 => conv_std_logic_vector(764, 16),
1216 => conv_std_logic_vector(768, 16),
1217 => conv_std_logic_vector(772, 16),
1218 => conv_std_logic_vector(776, 16),
1219 => conv_std_logic_vector(780, 16),
1220 => conv_std_logic_vector(784, 16),
1221 => conv_std_logic_vector(788, 16),
1222 => conv_std_logic_vector(792, 16),
1223 => conv_std_logic_vector(796, 16),
1224 => conv_std_logic_vector(800, 16),
1225 => conv_std_logic_vector(804, 16),
1226 => conv_std_logic_vector(808, 16),
1227 => conv_std_logic_vector(812, 16),
1228 => conv_std_logic_vector(816, 16),
1229 => conv_std_logic_vector(820, 16),
1230 => conv_std_logic_vector(824, 16),
1231 => conv_std_logic_vector(828, 16),
1232 => conv_std_logic_vector(832, 16),
1233 => conv_std_logic_vector(836, 16),
1234 => conv_std_logic_vector(840, 16),
1235 => conv_std_logic_vector(844, 16),
1236 => conv_std_logic_vector(848, 16),
1237 => conv_std_logic_vector(852, 16),
1238 => conv_std_logic_vector(856, 16),
1239 => conv_std_logic_vector(860, 16),
1240 => conv_std_logic_vector(864, 16),
1241 => conv_std_logic_vector(868, 16),
1242 => conv_std_logic_vector(872, 16),
1243 => conv_std_logic_vector(876, 16),
1244 => conv_std_logic_vector(880, 16),
1245 => conv_std_logic_vector(884, 16),
1246 => conv_std_logic_vector(888, 16),
1247 => conv_std_logic_vector(892, 16),
1248 => conv_std_logic_vector(896, 16),
1249 => conv_std_logic_vector(900, 16),
1250 => conv_std_logic_vector(904, 16),
1251 => conv_std_logic_vector(908, 16),
1252 => conv_std_logic_vector(912, 16),
1253 => conv_std_logic_vector(916, 16),
1254 => conv_std_logic_vector(920, 16),
1255 => conv_std_logic_vector(924, 16),
1256 => conv_std_logic_vector(928, 16),
1257 => conv_std_logic_vector(932, 16),
1258 => conv_std_logic_vector(936, 16),
1259 => conv_std_logic_vector(940, 16),
1260 => conv_std_logic_vector(944, 16),
1261 => conv_std_logic_vector(948, 16),
1262 => conv_std_logic_vector(952, 16),
1263 => conv_std_logic_vector(956, 16),
1264 => conv_std_logic_vector(960, 16),
1265 => conv_std_logic_vector(964, 16),
1266 => conv_std_logic_vector(968, 16),
1267 => conv_std_logic_vector(972, 16),
1268 => conv_std_logic_vector(976, 16),
1269 => conv_std_logic_vector(980, 16),
1270 => conv_std_logic_vector(984, 16),
1271 => conv_std_logic_vector(988, 16),
1272 => conv_std_logic_vector(992, 16),
1273 => conv_std_logic_vector(996, 16),
1274 => conv_std_logic_vector(1000, 16),
1275 => conv_std_logic_vector(1004, 16),
1276 => conv_std_logic_vector(1008, 16),
1277 => conv_std_logic_vector(1012, 16),
1278 => conv_std_logic_vector(1016, 16),
1279 => conv_std_logic_vector(1020, 16),
1280 => conv_std_logic_vector(0, 16),
1281 => conv_std_logic_vector(5, 16),
1282 => conv_std_logic_vector(10, 16),
1283 => conv_std_logic_vector(15, 16),
1284 => conv_std_logic_vector(20, 16),
1285 => conv_std_logic_vector(25, 16),
1286 => conv_std_logic_vector(30, 16),
1287 => conv_std_logic_vector(35, 16),
1288 => conv_std_logic_vector(40, 16),
1289 => conv_std_logic_vector(45, 16),
1290 => conv_std_logic_vector(50, 16),
1291 => conv_std_logic_vector(55, 16),
1292 => conv_std_logic_vector(60, 16),
1293 => conv_std_logic_vector(65, 16),
1294 => conv_std_logic_vector(70, 16),
1295 => conv_std_logic_vector(75, 16),
1296 => conv_std_logic_vector(80, 16),
1297 => conv_std_logic_vector(85, 16),
1298 => conv_std_logic_vector(90, 16),
1299 => conv_std_logic_vector(95, 16),
1300 => conv_std_logic_vector(100, 16),
1301 => conv_std_logic_vector(105, 16),
1302 => conv_std_logic_vector(110, 16),
1303 => conv_std_logic_vector(115, 16),
1304 => conv_std_logic_vector(120, 16),
1305 => conv_std_logic_vector(125, 16),
1306 => conv_std_logic_vector(130, 16),
1307 => conv_std_logic_vector(135, 16),
1308 => conv_std_logic_vector(140, 16),
1309 => conv_std_logic_vector(145, 16),
1310 => conv_std_logic_vector(150, 16),
1311 => conv_std_logic_vector(155, 16),
1312 => conv_std_logic_vector(160, 16),
1313 => conv_std_logic_vector(165, 16),
1314 => conv_std_logic_vector(170, 16),
1315 => conv_std_logic_vector(175, 16),
1316 => conv_std_logic_vector(180, 16),
1317 => conv_std_logic_vector(185, 16),
1318 => conv_std_logic_vector(190, 16),
1319 => conv_std_logic_vector(195, 16),
1320 => conv_std_logic_vector(200, 16),
1321 => conv_std_logic_vector(205, 16),
1322 => conv_std_logic_vector(210, 16),
1323 => conv_std_logic_vector(215, 16),
1324 => conv_std_logic_vector(220, 16),
1325 => conv_std_logic_vector(225, 16),
1326 => conv_std_logic_vector(230, 16),
1327 => conv_std_logic_vector(235, 16),
1328 => conv_std_logic_vector(240, 16),
1329 => conv_std_logic_vector(245, 16),
1330 => conv_std_logic_vector(250, 16),
1331 => conv_std_logic_vector(255, 16),
1332 => conv_std_logic_vector(260, 16),
1333 => conv_std_logic_vector(265, 16),
1334 => conv_std_logic_vector(270, 16),
1335 => conv_std_logic_vector(275, 16),
1336 => conv_std_logic_vector(280, 16),
1337 => conv_std_logic_vector(285, 16),
1338 => conv_std_logic_vector(290, 16),
1339 => conv_std_logic_vector(295, 16),
1340 => conv_std_logic_vector(300, 16),
1341 => conv_std_logic_vector(305, 16),
1342 => conv_std_logic_vector(310, 16),
1343 => conv_std_logic_vector(315, 16),
1344 => conv_std_logic_vector(320, 16),
1345 => conv_std_logic_vector(325, 16),
1346 => conv_std_logic_vector(330, 16),
1347 => conv_std_logic_vector(335, 16),
1348 => conv_std_logic_vector(340, 16),
1349 => conv_std_logic_vector(345, 16),
1350 => conv_std_logic_vector(350, 16),
1351 => conv_std_logic_vector(355, 16),
1352 => conv_std_logic_vector(360, 16),
1353 => conv_std_logic_vector(365, 16),
1354 => conv_std_logic_vector(370, 16),
1355 => conv_std_logic_vector(375, 16),
1356 => conv_std_logic_vector(380, 16),
1357 => conv_std_logic_vector(385, 16),
1358 => conv_std_logic_vector(390, 16),
1359 => conv_std_logic_vector(395, 16),
1360 => conv_std_logic_vector(400, 16),
1361 => conv_std_logic_vector(405, 16),
1362 => conv_std_logic_vector(410, 16),
1363 => conv_std_logic_vector(415, 16),
1364 => conv_std_logic_vector(420, 16),
1365 => conv_std_logic_vector(425, 16),
1366 => conv_std_logic_vector(430, 16),
1367 => conv_std_logic_vector(435, 16),
1368 => conv_std_logic_vector(440, 16),
1369 => conv_std_logic_vector(445, 16),
1370 => conv_std_logic_vector(450, 16),
1371 => conv_std_logic_vector(455, 16),
1372 => conv_std_logic_vector(460, 16),
1373 => conv_std_logic_vector(465, 16),
1374 => conv_std_logic_vector(470, 16),
1375 => conv_std_logic_vector(475, 16),
1376 => conv_std_logic_vector(480, 16),
1377 => conv_std_logic_vector(485, 16),
1378 => conv_std_logic_vector(490, 16),
1379 => conv_std_logic_vector(495, 16),
1380 => conv_std_logic_vector(500, 16),
1381 => conv_std_logic_vector(505, 16),
1382 => conv_std_logic_vector(510, 16),
1383 => conv_std_logic_vector(515, 16),
1384 => conv_std_logic_vector(520, 16),
1385 => conv_std_logic_vector(525, 16),
1386 => conv_std_logic_vector(530, 16),
1387 => conv_std_logic_vector(535, 16),
1388 => conv_std_logic_vector(540, 16),
1389 => conv_std_logic_vector(545, 16),
1390 => conv_std_logic_vector(550, 16),
1391 => conv_std_logic_vector(555, 16),
1392 => conv_std_logic_vector(560, 16),
1393 => conv_std_logic_vector(565, 16),
1394 => conv_std_logic_vector(570, 16),
1395 => conv_std_logic_vector(575, 16),
1396 => conv_std_logic_vector(580, 16),
1397 => conv_std_logic_vector(585, 16),
1398 => conv_std_logic_vector(590, 16),
1399 => conv_std_logic_vector(595, 16),
1400 => conv_std_logic_vector(600, 16),
1401 => conv_std_logic_vector(605, 16),
1402 => conv_std_logic_vector(610, 16),
1403 => conv_std_logic_vector(615, 16),
1404 => conv_std_logic_vector(620, 16),
1405 => conv_std_logic_vector(625, 16),
1406 => conv_std_logic_vector(630, 16),
1407 => conv_std_logic_vector(635, 16),
1408 => conv_std_logic_vector(640, 16),
1409 => conv_std_logic_vector(645, 16),
1410 => conv_std_logic_vector(650, 16),
1411 => conv_std_logic_vector(655, 16),
1412 => conv_std_logic_vector(660, 16),
1413 => conv_std_logic_vector(665, 16),
1414 => conv_std_logic_vector(670, 16),
1415 => conv_std_logic_vector(675, 16),
1416 => conv_std_logic_vector(680, 16),
1417 => conv_std_logic_vector(685, 16),
1418 => conv_std_logic_vector(690, 16),
1419 => conv_std_logic_vector(695, 16),
1420 => conv_std_logic_vector(700, 16),
1421 => conv_std_logic_vector(705, 16),
1422 => conv_std_logic_vector(710, 16),
1423 => conv_std_logic_vector(715, 16),
1424 => conv_std_logic_vector(720, 16),
1425 => conv_std_logic_vector(725, 16),
1426 => conv_std_logic_vector(730, 16),
1427 => conv_std_logic_vector(735, 16),
1428 => conv_std_logic_vector(740, 16),
1429 => conv_std_logic_vector(745, 16),
1430 => conv_std_logic_vector(750, 16),
1431 => conv_std_logic_vector(755, 16),
1432 => conv_std_logic_vector(760, 16),
1433 => conv_std_logic_vector(765, 16),
1434 => conv_std_logic_vector(770, 16),
1435 => conv_std_logic_vector(775, 16),
1436 => conv_std_logic_vector(780, 16),
1437 => conv_std_logic_vector(785, 16),
1438 => conv_std_logic_vector(790, 16),
1439 => conv_std_logic_vector(795, 16),
1440 => conv_std_logic_vector(800, 16),
1441 => conv_std_logic_vector(805, 16),
1442 => conv_std_logic_vector(810, 16),
1443 => conv_std_logic_vector(815, 16),
1444 => conv_std_logic_vector(820, 16),
1445 => conv_std_logic_vector(825, 16),
1446 => conv_std_logic_vector(830, 16),
1447 => conv_std_logic_vector(835, 16),
1448 => conv_std_logic_vector(840, 16),
1449 => conv_std_logic_vector(845, 16),
1450 => conv_std_logic_vector(850, 16),
1451 => conv_std_logic_vector(855, 16),
1452 => conv_std_logic_vector(860, 16),
1453 => conv_std_logic_vector(865, 16),
1454 => conv_std_logic_vector(870, 16),
1455 => conv_std_logic_vector(875, 16),
1456 => conv_std_logic_vector(880, 16),
1457 => conv_std_logic_vector(885, 16),
1458 => conv_std_logic_vector(890, 16),
1459 => conv_std_logic_vector(895, 16),
1460 => conv_std_logic_vector(900, 16),
1461 => conv_std_logic_vector(905, 16),
1462 => conv_std_logic_vector(910, 16),
1463 => conv_std_logic_vector(915, 16),
1464 => conv_std_logic_vector(920, 16),
1465 => conv_std_logic_vector(925, 16),
1466 => conv_std_logic_vector(930, 16),
1467 => conv_std_logic_vector(935, 16),
1468 => conv_std_logic_vector(940, 16),
1469 => conv_std_logic_vector(945, 16),
1470 => conv_std_logic_vector(950, 16),
1471 => conv_std_logic_vector(955, 16),
1472 => conv_std_logic_vector(960, 16),
1473 => conv_std_logic_vector(965, 16),
1474 => conv_std_logic_vector(970, 16),
1475 => conv_std_logic_vector(975, 16),
1476 => conv_std_logic_vector(980, 16),
1477 => conv_std_logic_vector(985, 16),
1478 => conv_std_logic_vector(990, 16),
1479 => conv_std_logic_vector(995, 16),
1480 => conv_std_logic_vector(1000, 16),
1481 => conv_std_logic_vector(1005, 16),
1482 => conv_std_logic_vector(1010, 16),
1483 => conv_std_logic_vector(1015, 16),
1484 => conv_std_logic_vector(1020, 16),
1485 => conv_std_logic_vector(1025, 16),
1486 => conv_std_logic_vector(1030, 16),
1487 => conv_std_logic_vector(1035, 16),
1488 => conv_std_logic_vector(1040, 16),
1489 => conv_std_logic_vector(1045, 16),
1490 => conv_std_logic_vector(1050, 16),
1491 => conv_std_logic_vector(1055, 16),
1492 => conv_std_logic_vector(1060, 16),
1493 => conv_std_logic_vector(1065, 16),
1494 => conv_std_logic_vector(1070, 16),
1495 => conv_std_logic_vector(1075, 16),
1496 => conv_std_logic_vector(1080, 16),
1497 => conv_std_logic_vector(1085, 16),
1498 => conv_std_logic_vector(1090, 16),
1499 => conv_std_logic_vector(1095, 16),
1500 => conv_std_logic_vector(1100, 16),
1501 => conv_std_logic_vector(1105, 16),
1502 => conv_std_logic_vector(1110, 16),
1503 => conv_std_logic_vector(1115, 16),
1504 => conv_std_logic_vector(1120, 16),
1505 => conv_std_logic_vector(1125, 16),
1506 => conv_std_logic_vector(1130, 16),
1507 => conv_std_logic_vector(1135, 16),
1508 => conv_std_logic_vector(1140, 16),
1509 => conv_std_logic_vector(1145, 16),
1510 => conv_std_logic_vector(1150, 16),
1511 => conv_std_logic_vector(1155, 16),
1512 => conv_std_logic_vector(1160, 16),
1513 => conv_std_logic_vector(1165, 16),
1514 => conv_std_logic_vector(1170, 16),
1515 => conv_std_logic_vector(1175, 16),
1516 => conv_std_logic_vector(1180, 16),
1517 => conv_std_logic_vector(1185, 16),
1518 => conv_std_logic_vector(1190, 16),
1519 => conv_std_logic_vector(1195, 16),
1520 => conv_std_logic_vector(1200, 16),
1521 => conv_std_logic_vector(1205, 16),
1522 => conv_std_logic_vector(1210, 16),
1523 => conv_std_logic_vector(1215, 16),
1524 => conv_std_logic_vector(1220, 16),
1525 => conv_std_logic_vector(1225, 16),
1526 => conv_std_logic_vector(1230, 16),
1527 => conv_std_logic_vector(1235, 16),
1528 => conv_std_logic_vector(1240, 16),
1529 => conv_std_logic_vector(1245, 16),
1530 => conv_std_logic_vector(1250, 16),
1531 => conv_std_logic_vector(1255, 16),
1532 => conv_std_logic_vector(1260, 16),
1533 => conv_std_logic_vector(1265, 16),
1534 => conv_std_logic_vector(1270, 16),
1535 => conv_std_logic_vector(1275, 16),
1536 => conv_std_logic_vector(0, 16),
1537 => conv_std_logic_vector(6, 16),
1538 => conv_std_logic_vector(12, 16),
1539 => conv_std_logic_vector(18, 16),
1540 => conv_std_logic_vector(24, 16),
1541 => conv_std_logic_vector(30, 16),
1542 => conv_std_logic_vector(36, 16),
1543 => conv_std_logic_vector(42, 16),
1544 => conv_std_logic_vector(48, 16),
1545 => conv_std_logic_vector(54, 16),
1546 => conv_std_logic_vector(60, 16),
1547 => conv_std_logic_vector(66, 16),
1548 => conv_std_logic_vector(72, 16),
1549 => conv_std_logic_vector(78, 16),
1550 => conv_std_logic_vector(84, 16),
1551 => conv_std_logic_vector(90, 16),
1552 => conv_std_logic_vector(96, 16),
1553 => conv_std_logic_vector(102, 16),
1554 => conv_std_logic_vector(108, 16),
1555 => conv_std_logic_vector(114, 16),
1556 => conv_std_logic_vector(120, 16),
1557 => conv_std_logic_vector(126, 16),
1558 => conv_std_logic_vector(132, 16),
1559 => conv_std_logic_vector(138, 16),
1560 => conv_std_logic_vector(144, 16),
1561 => conv_std_logic_vector(150, 16),
1562 => conv_std_logic_vector(156, 16),
1563 => conv_std_logic_vector(162, 16),
1564 => conv_std_logic_vector(168, 16),
1565 => conv_std_logic_vector(174, 16),
1566 => conv_std_logic_vector(180, 16),
1567 => conv_std_logic_vector(186, 16),
1568 => conv_std_logic_vector(192, 16),
1569 => conv_std_logic_vector(198, 16),
1570 => conv_std_logic_vector(204, 16),
1571 => conv_std_logic_vector(210, 16),
1572 => conv_std_logic_vector(216, 16),
1573 => conv_std_logic_vector(222, 16),
1574 => conv_std_logic_vector(228, 16),
1575 => conv_std_logic_vector(234, 16),
1576 => conv_std_logic_vector(240, 16),
1577 => conv_std_logic_vector(246, 16),
1578 => conv_std_logic_vector(252, 16),
1579 => conv_std_logic_vector(258, 16),
1580 => conv_std_logic_vector(264, 16),
1581 => conv_std_logic_vector(270, 16),
1582 => conv_std_logic_vector(276, 16),
1583 => conv_std_logic_vector(282, 16),
1584 => conv_std_logic_vector(288, 16),
1585 => conv_std_logic_vector(294, 16),
1586 => conv_std_logic_vector(300, 16),
1587 => conv_std_logic_vector(306, 16),
1588 => conv_std_logic_vector(312, 16),
1589 => conv_std_logic_vector(318, 16),
1590 => conv_std_logic_vector(324, 16),
1591 => conv_std_logic_vector(330, 16),
1592 => conv_std_logic_vector(336, 16),
1593 => conv_std_logic_vector(342, 16),
1594 => conv_std_logic_vector(348, 16),
1595 => conv_std_logic_vector(354, 16),
1596 => conv_std_logic_vector(360, 16),
1597 => conv_std_logic_vector(366, 16),
1598 => conv_std_logic_vector(372, 16),
1599 => conv_std_logic_vector(378, 16),
1600 => conv_std_logic_vector(384, 16),
1601 => conv_std_logic_vector(390, 16),
1602 => conv_std_logic_vector(396, 16),
1603 => conv_std_logic_vector(402, 16),
1604 => conv_std_logic_vector(408, 16),
1605 => conv_std_logic_vector(414, 16),
1606 => conv_std_logic_vector(420, 16),
1607 => conv_std_logic_vector(426, 16),
1608 => conv_std_logic_vector(432, 16),
1609 => conv_std_logic_vector(438, 16),
1610 => conv_std_logic_vector(444, 16),
1611 => conv_std_logic_vector(450, 16),
1612 => conv_std_logic_vector(456, 16),
1613 => conv_std_logic_vector(462, 16),
1614 => conv_std_logic_vector(468, 16),
1615 => conv_std_logic_vector(474, 16),
1616 => conv_std_logic_vector(480, 16),
1617 => conv_std_logic_vector(486, 16),
1618 => conv_std_logic_vector(492, 16),
1619 => conv_std_logic_vector(498, 16),
1620 => conv_std_logic_vector(504, 16),
1621 => conv_std_logic_vector(510, 16),
1622 => conv_std_logic_vector(516, 16),
1623 => conv_std_logic_vector(522, 16),
1624 => conv_std_logic_vector(528, 16),
1625 => conv_std_logic_vector(534, 16),
1626 => conv_std_logic_vector(540, 16),
1627 => conv_std_logic_vector(546, 16),
1628 => conv_std_logic_vector(552, 16),
1629 => conv_std_logic_vector(558, 16),
1630 => conv_std_logic_vector(564, 16),
1631 => conv_std_logic_vector(570, 16),
1632 => conv_std_logic_vector(576, 16),
1633 => conv_std_logic_vector(582, 16),
1634 => conv_std_logic_vector(588, 16),
1635 => conv_std_logic_vector(594, 16),
1636 => conv_std_logic_vector(600, 16),
1637 => conv_std_logic_vector(606, 16),
1638 => conv_std_logic_vector(612, 16),
1639 => conv_std_logic_vector(618, 16),
1640 => conv_std_logic_vector(624, 16),
1641 => conv_std_logic_vector(630, 16),
1642 => conv_std_logic_vector(636, 16),
1643 => conv_std_logic_vector(642, 16),
1644 => conv_std_logic_vector(648, 16),
1645 => conv_std_logic_vector(654, 16),
1646 => conv_std_logic_vector(660, 16),
1647 => conv_std_logic_vector(666, 16),
1648 => conv_std_logic_vector(672, 16),
1649 => conv_std_logic_vector(678, 16),
1650 => conv_std_logic_vector(684, 16),
1651 => conv_std_logic_vector(690, 16),
1652 => conv_std_logic_vector(696, 16),
1653 => conv_std_logic_vector(702, 16),
1654 => conv_std_logic_vector(708, 16),
1655 => conv_std_logic_vector(714, 16),
1656 => conv_std_logic_vector(720, 16),
1657 => conv_std_logic_vector(726, 16),
1658 => conv_std_logic_vector(732, 16),
1659 => conv_std_logic_vector(738, 16),
1660 => conv_std_logic_vector(744, 16),
1661 => conv_std_logic_vector(750, 16),
1662 => conv_std_logic_vector(756, 16),
1663 => conv_std_logic_vector(762, 16),
1664 => conv_std_logic_vector(768, 16),
1665 => conv_std_logic_vector(774, 16),
1666 => conv_std_logic_vector(780, 16),
1667 => conv_std_logic_vector(786, 16),
1668 => conv_std_logic_vector(792, 16),
1669 => conv_std_logic_vector(798, 16),
1670 => conv_std_logic_vector(804, 16),
1671 => conv_std_logic_vector(810, 16),
1672 => conv_std_logic_vector(816, 16),
1673 => conv_std_logic_vector(822, 16),
1674 => conv_std_logic_vector(828, 16),
1675 => conv_std_logic_vector(834, 16),
1676 => conv_std_logic_vector(840, 16),
1677 => conv_std_logic_vector(846, 16),
1678 => conv_std_logic_vector(852, 16),
1679 => conv_std_logic_vector(858, 16),
1680 => conv_std_logic_vector(864, 16),
1681 => conv_std_logic_vector(870, 16),
1682 => conv_std_logic_vector(876, 16),
1683 => conv_std_logic_vector(882, 16),
1684 => conv_std_logic_vector(888, 16),
1685 => conv_std_logic_vector(894, 16),
1686 => conv_std_logic_vector(900, 16),
1687 => conv_std_logic_vector(906, 16),
1688 => conv_std_logic_vector(912, 16),
1689 => conv_std_logic_vector(918, 16),
1690 => conv_std_logic_vector(924, 16),
1691 => conv_std_logic_vector(930, 16),
1692 => conv_std_logic_vector(936, 16),
1693 => conv_std_logic_vector(942, 16),
1694 => conv_std_logic_vector(948, 16),
1695 => conv_std_logic_vector(954, 16),
1696 => conv_std_logic_vector(960, 16),
1697 => conv_std_logic_vector(966, 16),
1698 => conv_std_logic_vector(972, 16),
1699 => conv_std_logic_vector(978, 16),
1700 => conv_std_logic_vector(984, 16),
1701 => conv_std_logic_vector(990, 16),
1702 => conv_std_logic_vector(996, 16),
1703 => conv_std_logic_vector(1002, 16),
1704 => conv_std_logic_vector(1008, 16),
1705 => conv_std_logic_vector(1014, 16),
1706 => conv_std_logic_vector(1020, 16),
1707 => conv_std_logic_vector(1026, 16),
1708 => conv_std_logic_vector(1032, 16),
1709 => conv_std_logic_vector(1038, 16),
1710 => conv_std_logic_vector(1044, 16),
1711 => conv_std_logic_vector(1050, 16),
1712 => conv_std_logic_vector(1056, 16),
1713 => conv_std_logic_vector(1062, 16),
1714 => conv_std_logic_vector(1068, 16),
1715 => conv_std_logic_vector(1074, 16),
1716 => conv_std_logic_vector(1080, 16),
1717 => conv_std_logic_vector(1086, 16),
1718 => conv_std_logic_vector(1092, 16),
1719 => conv_std_logic_vector(1098, 16),
1720 => conv_std_logic_vector(1104, 16),
1721 => conv_std_logic_vector(1110, 16),
1722 => conv_std_logic_vector(1116, 16),
1723 => conv_std_logic_vector(1122, 16),
1724 => conv_std_logic_vector(1128, 16),
1725 => conv_std_logic_vector(1134, 16),
1726 => conv_std_logic_vector(1140, 16),
1727 => conv_std_logic_vector(1146, 16),
1728 => conv_std_logic_vector(1152, 16),
1729 => conv_std_logic_vector(1158, 16),
1730 => conv_std_logic_vector(1164, 16),
1731 => conv_std_logic_vector(1170, 16),
1732 => conv_std_logic_vector(1176, 16),
1733 => conv_std_logic_vector(1182, 16),
1734 => conv_std_logic_vector(1188, 16),
1735 => conv_std_logic_vector(1194, 16),
1736 => conv_std_logic_vector(1200, 16),
1737 => conv_std_logic_vector(1206, 16),
1738 => conv_std_logic_vector(1212, 16),
1739 => conv_std_logic_vector(1218, 16),
1740 => conv_std_logic_vector(1224, 16),
1741 => conv_std_logic_vector(1230, 16),
1742 => conv_std_logic_vector(1236, 16),
1743 => conv_std_logic_vector(1242, 16),
1744 => conv_std_logic_vector(1248, 16),
1745 => conv_std_logic_vector(1254, 16),
1746 => conv_std_logic_vector(1260, 16),
1747 => conv_std_logic_vector(1266, 16),
1748 => conv_std_logic_vector(1272, 16),
1749 => conv_std_logic_vector(1278, 16),
1750 => conv_std_logic_vector(1284, 16),
1751 => conv_std_logic_vector(1290, 16),
1752 => conv_std_logic_vector(1296, 16),
1753 => conv_std_logic_vector(1302, 16),
1754 => conv_std_logic_vector(1308, 16),
1755 => conv_std_logic_vector(1314, 16),
1756 => conv_std_logic_vector(1320, 16),
1757 => conv_std_logic_vector(1326, 16),
1758 => conv_std_logic_vector(1332, 16),
1759 => conv_std_logic_vector(1338, 16),
1760 => conv_std_logic_vector(1344, 16),
1761 => conv_std_logic_vector(1350, 16),
1762 => conv_std_logic_vector(1356, 16),
1763 => conv_std_logic_vector(1362, 16),
1764 => conv_std_logic_vector(1368, 16),
1765 => conv_std_logic_vector(1374, 16),
1766 => conv_std_logic_vector(1380, 16),
1767 => conv_std_logic_vector(1386, 16),
1768 => conv_std_logic_vector(1392, 16),
1769 => conv_std_logic_vector(1398, 16),
1770 => conv_std_logic_vector(1404, 16),
1771 => conv_std_logic_vector(1410, 16),
1772 => conv_std_logic_vector(1416, 16),
1773 => conv_std_logic_vector(1422, 16),
1774 => conv_std_logic_vector(1428, 16),
1775 => conv_std_logic_vector(1434, 16),
1776 => conv_std_logic_vector(1440, 16),
1777 => conv_std_logic_vector(1446, 16),
1778 => conv_std_logic_vector(1452, 16),
1779 => conv_std_logic_vector(1458, 16),
1780 => conv_std_logic_vector(1464, 16),
1781 => conv_std_logic_vector(1470, 16),
1782 => conv_std_logic_vector(1476, 16),
1783 => conv_std_logic_vector(1482, 16),
1784 => conv_std_logic_vector(1488, 16),
1785 => conv_std_logic_vector(1494, 16),
1786 => conv_std_logic_vector(1500, 16),
1787 => conv_std_logic_vector(1506, 16),
1788 => conv_std_logic_vector(1512, 16),
1789 => conv_std_logic_vector(1518, 16),
1790 => conv_std_logic_vector(1524, 16),
1791 => conv_std_logic_vector(1530, 16),
1792 => conv_std_logic_vector(0, 16),
1793 => conv_std_logic_vector(7, 16),
1794 => conv_std_logic_vector(14, 16),
1795 => conv_std_logic_vector(21, 16),
1796 => conv_std_logic_vector(28, 16),
1797 => conv_std_logic_vector(35, 16),
1798 => conv_std_logic_vector(42, 16),
1799 => conv_std_logic_vector(49, 16),
1800 => conv_std_logic_vector(56, 16),
1801 => conv_std_logic_vector(63, 16),
1802 => conv_std_logic_vector(70, 16),
1803 => conv_std_logic_vector(77, 16),
1804 => conv_std_logic_vector(84, 16),
1805 => conv_std_logic_vector(91, 16),
1806 => conv_std_logic_vector(98, 16),
1807 => conv_std_logic_vector(105, 16),
1808 => conv_std_logic_vector(112, 16),
1809 => conv_std_logic_vector(119, 16),
1810 => conv_std_logic_vector(126, 16),
1811 => conv_std_logic_vector(133, 16),
1812 => conv_std_logic_vector(140, 16),
1813 => conv_std_logic_vector(147, 16),
1814 => conv_std_logic_vector(154, 16),
1815 => conv_std_logic_vector(161, 16),
1816 => conv_std_logic_vector(168, 16),
1817 => conv_std_logic_vector(175, 16),
1818 => conv_std_logic_vector(182, 16),
1819 => conv_std_logic_vector(189, 16),
1820 => conv_std_logic_vector(196, 16),
1821 => conv_std_logic_vector(203, 16),
1822 => conv_std_logic_vector(210, 16),
1823 => conv_std_logic_vector(217, 16),
1824 => conv_std_logic_vector(224, 16),
1825 => conv_std_logic_vector(231, 16),
1826 => conv_std_logic_vector(238, 16),
1827 => conv_std_logic_vector(245, 16),
1828 => conv_std_logic_vector(252, 16),
1829 => conv_std_logic_vector(259, 16),
1830 => conv_std_logic_vector(266, 16),
1831 => conv_std_logic_vector(273, 16),
1832 => conv_std_logic_vector(280, 16),
1833 => conv_std_logic_vector(287, 16),
1834 => conv_std_logic_vector(294, 16),
1835 => conv_std_logic_vector(301, 16),
1836 => conv_std_logic_vector(308, 16),
1837 => conv_std_logic_vector(315, 16),
1838 => conv_std_logic_vector(322, 16),
1839 => conv_std_logic_vector(329, 16),
1840 => conv_std_logic_vector(336, 16),
1841 => conv_std_logic_vector(343, 16),
1842 => conv_std_logic_vector(350, 16),
1843 => conv_std_logic_vector(357, 16),
1844 => conv_std_logic_vector(364, 16),
1845 => conv_std_logic_vector(371, 16),
1846 => conv_std_logic_vector(378, 16),
1847 => conv_std_logic_vector(385, 16),
1848 => conv_std_logic_vector(392, 16),
1849 => conv_std_logic_vector(399, 16),
1850 => conv_std_logic_vector(406, 16),
1851 => conv_std_logic_vector(413, 16),
1852 => conv_std_logic_vector(420, 16),
1853 => conv_std_logic_vector(427, 16),
1854 => conv_std_logic_vector(434, 16),
1855 => conv_std_logic_vector(441, 16),
1856 => conv_std_logic_vector(448, 16),
1857 => conv_std_logic_vector(455, 16),
1858 => conv_std_logic_vector(462, 16),
1859 => conv_std_logic_vector(469, 16),
1860 => conv_std_logic_vector(476, 16),
1861 => conv_std_logic_vector(483, 16),
1862 => conv_std_logic_vector(490, 16),
1863 => conv_std_logic_vector(497, 16),
1864 => conv_std_logic_vector(504, 16),
1865 => conv_std_logic_vector(511, 16),
1866 => conv_std_logic_vector(518, 16),
1867 => conv_std_logic_vector(525, 16),
1868 => conv_std_logic_vector(532, 16),
1869 => conv_std_logic_vector(539, 16),
1870 => conv_std_logic_vector(546, 16),
1871 => conv_std_logic_vector(553, 16),
1872 => conv_std_logic_vector(560, 16),
1873 => conv_std_logic_vector(567, 16),
1874 => conv_std_logic_vector(574, 16),
1875 => conv_std_logic_vector(581, 16),
1876 => conv_std_logic_vector(588, 16),
1877 => conv_std_logic_vector(595, 16),
1878 => conv_std_logic_vector(602, 16),
1879 => conv_std_logic_vector(609, 16),
1880 => conv_std_logic_vector(616, 16),
1881 => conv_std_logic_vector(623, 16),
1882 => conv_std_logic_vector(630, 16),
1883 => conv_std_logic_vector(637, 16),
1884 => conv_std_logic_vector(644, 16),
1885 => conv_std_logic_vector(651, 16),
1886 => conv_std_logic_vector(658, 16),
1887 => conv_std_logic_vector(665, 16),
1888 => conv_std_logic_vector(672, 16),
1889 => conv_std_logic_vector(679, 16),
1890 => conv_std_logic_vector(686, 16),
1891 => conv_std_logic_vector(693, 16),
1892 => conv_std_logic_vector(700, 16),
1893 => conv_std_logic_vector(707, 16),
1894 => conv_std_logic_vector(714, 16),
1895 => conv_std_logic_vector(721, 16),
1896 => conv_std_logic_vector(728, 16),
1897 => conv_std_logic_vector(735, 16),
1898 => conv_std_logic_vector(742, 16),
1899 => conv_std_logic_vector(749, 16),
1900 => conv_std_logic_vector(756, 16),
1901 => conv_std_logic_vector(763, 16),
1902 => conv_std_logic_vector(770, 16),
1903 => conv_std_logic_vector(777, 16),
1904 => conv_std_logic_vector(784, 16),
1905 => conv_std_logic_vector(791, 16),
1906 => conv_std_logic_vector(798, 16),
1907 => conv_std_logic_vector(805, 16),
1908 => conv_std_logic_vector(812, 16),
1909 => conv_std_logic_vector(819, 16),
1910 => conv_std_logic_vector(826, 16),
1911 => conv_std_logic_vector(833, 16),
1912 => conv_std_logic_vector(840, 16),
1913 => conv_std_logic_vector(847, 16),
1914 => conv_std_logic_vector(854, 16),
1915 => conv_std_logic_vector(861, 16),
1916 => conv_std_logic_vector(868, 16),
1917 => conv_std_logic_vector(875, 16),
1918 => conv_std_logic_vector(882, 16),
1919 => conv_std_logic_vector(889, 16),
1920 => conv_std_logic_vector(896, 16),
1921 => conv_std_logic_vector(903, 16),
1922 => conv_std_logic_vector(910, 16),
1923 => conv_std_logic_vector(917, 16),
1924 => conv_std_logic_vector(924, 16),
1925 => conv_std_logic_vector(931, 16),
1926 => conv_std_logic_vector(938, 16),
1927 => conv_std_logic_vector(945, 16),
1928 => conv_std_logic_vector(952, 16),
1929 => conv_std_logic_vector(959, 16),
1930 => conv_std_logic_vector(966, 16),
1931 => conv_std_logic_vector(973, 16),
1932 => conv_std_logic_vector(980, 16),
1933 => conv_std_logic_vector(987, 16),
1934 => conv_std_logic_vector(994, 16),
1935 => conv_std_logic_vector(1001, 16),
1936 => conv_std_logic_vector(1008, 16),
1937 => conv_std_logic_vector(1015, 16),
1938 => conv_std_logic_vector(1022, 16),
1939 => conv_std_logic_vector(1029, 16),
1940 => conv_std_logic_vector(1036, 16),
1941 => conv_std_logic_vector(1043, 16),
1942 => conv_std_logic_vector(1050, 16),
1943 => conv_std_logic_vector(1057, 16),
1944 => conv_std_logic_vector(1064, 16),
1945 => conv_std_logic_vector(1071, 16),
1946 => conv_std_logic_vector(1078, 16),
1947 => conv_std_logic_vector(1085, 16),
1948 => conv_std_logic_vector(1092, 16),
1949 => conv_std_logic_vector(1099, 16),
1950 => conv_std_logic_vector(1106, 16),
1951 => conv_std_logic_vector(1113, 16),
1952 => conv_std_logic_vector(1120, 16),
1953 => conv_std_logic_vector(1127, 16),
1954 => conv_std_logic_vector(1134, 16),
1955 => conv_std_logic_vector(1141, 16),
1956 => conv_std_logic_vector(1148, 16),
1957 => conv_std_logic_vector(1155, 16),
1958 => conv_std_logic_vector(1162, 16),
1959 => conv_std_logic_vector(1169, 16),
1960 => conv_std_logic_vector(1176, 16),
1961 => conv_std_logic_vector(1183, 16),
1962 => conv_std_logic_vector(1190, 16),
1963 => conv_std_logic_vector(1197, 16),
1964 => conv_std_logic_vector(1204, 16),
1965 => conv_std_logic_vector(1211, 16),
1966 => conv_std_logic_vector(1218, 16),
1967 => conv_std_logic_vector(1225, 16),
1968 => conv_std_logic_vector(1232, 16),
1969 => conv_std_logic_vector(1239, 16),
1970 => conv_std_logic_vector(1246, 16),
1971 => conv_std_logic_vector(1253, 16),
1972 => conv_std_logic_vector(1260, 16),
1973 => conv_std_logic_vector(1267, 16),
1974 => conv_std_logic_vector(1274, 16),
1975 => conv_std_logic_vector(1281, 16),
1976 => conv_std_logic_vector(1288, 16),
1977 => conv_std_logic_vector(1295, 16),
1978 => conv_std_logic_vector(1302, 16),
1979 => conv_std_logic_vector(1309, 16),
1980 => conv_std_logic_vector(1316, 16),
1981 => conv_std_logic_vector(1323, 16),
1982 => conv_std_logic_vector(1330, 16),
1983 => conv_std_logic_vector(1337, 16),
1984 => conv_std_logic_vector(1344, 16),
1985 => conv_std_logic_vector(1351, 16),
1986 => conv_std_logic_vector(1358, 16),
1987 => conv_std_logic_vector(1365, 16),
1988 => conv_std_logic_vector(1372, 16),
1989 => conv_std_logic_vector(1379, 16),
1990 => conv_std_logic_vector(1386, 16),
1991 => conv_std_logic_vector(1393, 16),
1992 => conv_std_logic_vector(1400, 16),
1993 => conv_std_logic_vector(1407, 16),
1994 => conv_std_logic_vector(1414, 16),
1995 => conv_std_logic_vector(1421, 16),
1996 => conv_std_logic_vector(1428, 16),
1997 => conv_std_logic_vector(1435, 16),
1998 => conv_std_logic_vector(1442, 16),
1999 => conv_std_logic_vector(1449, 16),
2000 => conv_std_logic_vector(1456, 16),
2001 => conv_std_logic_vector(1463, 16),
2002 => conv_std_logic_vector(1470, 16),
2003 => conv_std_logic_vector(1477, 16),
2004 => conv_std_logic_vector(1484, 16),
2005 => conv_std_logic_vector(1491, 16),
2006 => conv_std_logic_vector(1498, 16),
2007 => conv_std_logic_vector(1505, 16),
2008 => conv_std_logic_vector(1512, 16),
2009 => conv_std_logic_vector(1519, 16),
2010 => conv_std_logic_vector(1526, 16),
2011 => conv_std_logic_vector(1533, 16),
2012 => conv_std_logic_vector(1540, 16),
2013 => conv_std_logic_vector(1547, 16),
2014 => conv_std_logic_vector(1554, 16),
2015 => conv_std_logic_vector(1561, 16),
2016 => conv_std_logic_vector(1568, 16),
2017 => conv_std_logic_vector(1575, 16),
2018 => conv_std_logic_vector(1582, 16),
2019 => conv_std_logic_vector(1589, 16),
2020 => conv_std_logic_vector(1596, 16),
2021 => conv_std_logic_vector(1603, 16),
2022 => conv_std_logic_vector(1610, 16),
2023 => conv_std_logic_vector(1617, 16),
2024 => conv_std_logic_vector(1624, 16),
2025 => conv_std_logic_vector(1631, 16),
2026 => conv_std_logic_vector(1638, 16),
2027 => conv_std_logic_vector(1645, 16),
2028 => conv_std_logic_vector(1652, 16),
2029 => conv_std_logic_vector(1659, 16),
2030 => conv_std_logic_vector(1666, 16),
2031 => conv_std_logic_vector(1673, 16),
2032 => conv_std_logic_vector(1680, 16),
2033 => conv_std_logic_vector(1687, 16),
2034 => conv_std_logic_vector(1694, 16),
2035 => conv_std_logic_vector(1701, 16),
2036 => conv_std_logic_vector(1708, 16),
2037 => conv_std_logic_vector(1715, 16),
2038 => conv_std_logic_vector(1722, 16),
2039 => conv_std_logic_vector(1729, 16),
2040 => conv_std_logic_vector(1736, 16),
2041 => conv_std_logic_vector(1743, 16),
2042 => conv_std_logic_vector(1750, 16),
2043 => conv_std_logic_vector(1757, 16),
2044 => conv_std_logic_vector(1764, 16),
2045 => conv_std_logic_vector(1771, 16),
2046 => conv_std_logic_vector(1778, 16),
2047 => conv_std_logic_vector(1785, 16),
2048 => conv_std_logic_vector(0, 16),
2049 => conv_std_logic_vector(8, 16),
2050 => conv_std_logic_vector(16, 16),
2051 => conv_std_logic_vector(24, 16),
2052 => conv_std_logic_vector(32, 16),
2053 => conv_std_logic_vector(40, 16),
2054 => conv_std_logic_vector(48, 16),
2055 => conv_std_logic_vector(56, 16),
2056 => conv_std_logic_vector(64, 16),
2057 => conv_std_logic_vector(72, 16),
2058 => conv_std_logic_vector(80, 16),
2059 => conv_std_logic_vector(88, 16),
2060 => conv_std_logic_vector(96, 16),
2061 => conv_std_logic_vector(104, 16),
2062 => conv_std_logic_vector(112, 16),
2063 => conv_std_logic_vector(120, 16),
2064 => conv_std_logic_vector(128, 16),
2065 => conv_std_logic_vector(136, 16),
2066 => conv_std_logic_vector(144, 16),
2067 => conv_std_logic_vector(152, 16),
2068 => conv_std_logic_vector(160, 16),
2069 => conv_std_logic_vector(168, 16),
2070 => conv_std_logic_vector(176, 16),
2071 => conv_std_logic_vector(184, 16),
2072 => conv_std_logic_vector(192, 16),
2073 => conv_std_logic_vector(200, 16),
2074 => conv_std_logic_vector(208, 16),
2075 => conv_std_logic_vector(216, 16),
2076 => conv_std_logic_vector(224, 16),
2077 => conv_std_logic_vector(232, 16),
2078 => conv_std_logic_vector(240, 16),
2079 => conv_std_logic_vector(248, 16),
2080 => conv_std_logic_vector(256, 16),
2081 => conv_std_logic_vector(264, 16),
2082 => conv_std_logic_vector(272, 16),
2083 => conv_std_logic_vector(280, 16),
2084 => conv_std_logic_vector(288, 16),
2085 => conv_std_logic_vector(296, 16),
2086 => conv_std_logic_vector(304, 16),
2087 => conv_std_logic_vector(312, 16),
2088 => conv_std_logic_vector(320, 16),
2089 => conv_std_logic_vector(328, 16),
2090 => conv_std_logic_vector(336, 16),
2091 => conv_std_logic_vector(344, 16),
2092 => conv_std_logic_vector(352, 16),
2093 => conv_std_logic_vector(360, 16),
2094 => conv_std_logic_vector(368, 16),
2095 => conv_std_logic_vector(376, 16),
2096 => conv_std_logic_vector(384, 16),
2097 => conv_std_logic_vector(392, 16),
2098 => conv_std_logic_vector(400, 16),
2099 => conv_std_logic_vector(408, 16),
2100 => conv_std_logic_vector(416, 16),
2101 => conv_std_logic_vector(424, 16),
2102 => conv_std_logic_vector(432, 16),
2103 => conv_std_logic_vector(440, 16),
2104 => conv_std_logic_vector(448, 16),
2105 => conv_std_logic_vector(456, 16),
2106 => conv_std_logic_vector(464, 16),
2107 => conv_std_logic_vector(472, 16),
2108 => conv_std_logic_vector(480, 16),
2109 => conv_std_logic_vector(488, 16),
2110 => conv_std_logic_vector(496, 16),
2111 => conv_std_logic_vector(504, 16),
2112 => conv_std_logic_vector(512, 16),
2113 => conv_std_logic_vector(520, 16),
2114 => conv_std_logic_vector(528, 16),
2115 => conv_std_logic_vector(536, 16),
2116 => conv_std_logic_vector(544, 16),
2117 => conv_std_logic_vector(552, 16),
2118 => conv_std_logic_vector(560, 16),
2119 => conv_std_logic_vector(568, 16),
2120 => conv_std_logic_vector(576, 16),
2121 => conv_std_logic_vector(584, 16),
2122 => conv_std_logic_vector(592, 16),
2123 => conv_std_logic_vector(600, 16),
2124 => conv_std_logic_vector(608, 16),
2125 => conv_std_logic_vector(616, 16),
2126 => conv_std_logic_vector(624, 16),
2127 => conv_std_logic_vector(632, 16),
2128 => conv_std_logic_vector(640, 16),
2129 => conv_std_logic_vector(648, 16),
2130 => conv_std_logic_vector(656, 16),
2131 => conv_std_logic_vector(664, 16),
2132 => conv_std_logic_vector(672, 16),
2133 => conv_std_logic_vector(680, 16),
2134 => conv_std_logic_vector(688, 16),
2135 => conv_std_logic_vector(696, 16),
2136 => conv_std_logic_vector(704, 16),
2137 => conv_std_logic_vector(712, 16),
2138 => conv_std_logic_vector(720, 16),
2139 => conv_std_logic_vector(728, 16),
2140 => conv_std_logic_vector(736, 16),
2141 => conv_std_logic_vector(744, 16),
2142 => conv_std_logic_vector(752, 16),
2143 => conv_std_logic_vector(760, 16),
2144 => conv_std_logic_vector(768, 16),
2145 => conv_std_logic_vector(776, 16),
2146 => conv_std_logic_vector(784, 16),
2147 => conv_std_logic_vector(792, 16),
2148 => conv_std_logic_vector(800, 16),
2149 => conv_std_logic_vector(808, 16),
2150 => conv_std_logic_vector(816, 16),
2151 => conv_std_logic_vector(824, 16),
2152 => conv_std_logic_vector(832, 16),
2153 => conv_std_logic_vector(840, 16),
2154 => conv_std_logic_vector(848, 16),
2155 => conv_std_logic_vector(856, 16),
2156 => conv_std_logic_vector(864, 16),
2157 => conv_std_logic_vector(872, 16),
2158 => conv_std_logic_vector(880, 16),
2159 => conv_std_logic_vector(888, 16),
2160 => conv_std_logic_vector(896, 16),
2161 => conv_std_logic_vector(904, 16),
2162 => conv_std_logic_vector(912, 16),
2163 => conv_std_logic_vector(920, 16),
2164 => conv_std_logic_vector(928, 16),
2165 => conv_std_logic_vector(936, 16),
2166 => conv_std_logic_vector(944, 16),
2167 => conv_std_logic_vector(952, 16),
2168 => conv_std_logic_vector(960, 16),
2169 => conv_std_logic_vector(968, 16),
2170 => conv_std_logic_vector(976, 16),
2171 => conv_std_logic_vector(984, 16),
2172 => conv_std_logic_vector(992, 16),
2173 => conv_std_logic_vector(1000, 16),
2174 => conv_std_logic_vector(1008, 16),
2175 => conv_std_logic_vector(1016, 16),
2176 => conv_std_logic_vector(1024, 16),
2177 => conv_std_logic_vector(1032, 16),
2178 => conv_std_logic_vector(1040, 16),
2179 => conv_std_logic_vector(1048, 16),
2180 => conv_std_logic_vector(1056, 16),
2181 => conv_std_logic_vector(1064, 16),
2182 => conv_std_logic_vector(1072, 16),
2183 => conv_std_logic_vector(1080, 16),
2184 => conv_std_logic_vector(1088, 16),
2185 => conv_std_logic_vector(1096, 16),
2186 => conv_std_logic_vector(1104, 16),
2187 => conv_std_logic_vector(1112, 16),
2188 => conv_std_logic_vector(1120, 16),
2189 => conv_std_logic_vector(1128, 16),
2190 => conv_std_logic_vector(1136, 16),
2191 => conv_std_logic_vector(1144, 16),
2192 => conv_std_logic_vector(1152, 16),
2193 => conv_std_logic_vector(1160, 16),
2194 => conv_std_logic_vector(1168, 16),
2195 => conv_std_logic_vector(1176, 16),
2196 => conv_std_logic_vector(1184, 16),
2197 => conv_std_logic_vector(1192, 16),
2198 => conv_std_logic_vector(1200, 16),
2199 => conv_std_logic_vector(1208, 16),
2200 => conv_std_logic_vector(1216, 16),
2201 => conv_std_logic_vector(1224, 16),
2202 => conv_std_logic_vector(1232, 16),
2203 => conv_std_logic_vector(1240, 16),
2204 => conv_std_logic_vector(1248, 16),
2205 => conv_std_logic_vector(1256, 16),
2206 => conv_std_logic_vector(1264, 16),
2207 => conv_std_logic_vector(1272, 16),
2208 => conv_std_logic_vector(1280, 16),
2209 => conv_std_logic_vector(1288, 16),
2210 => conv_std_logic_vector(1296, 16),
2211 => conv_std_logic_vector(1304, 16),
2212 => conv_std_logic_vector(1312, 16),
2213 => conv_std_logic_vector(1320, 16),
2214 => conv_std_logic_vector(1328, 16),
2215 => conv_std_logic_vector(1336, 16),
2216 => conv_std_logic_vector(1344, 16),
2217 => conv_std_logic_vector(1352, 16),
2218 => conv_std_logic_vector(1360, 16),
2219 => conv_std_logic_vector(1368, 16),
2220 => conv_std_logic_vector(1376, 16),
2221 => conv_std_logic_vector(1384, 16),
2222 => conv_std_logic_vector(1392, 16),
2223 => conv_std_logic_vector(1400, 16),
2224 => conv_std_logic_vector(1408, 16),
2225 => conv_std_logic_vector(1416, 16),
2226 => conv_std_logic_vector(1424, 16),
2227 => conv_std_logic_vector(1432, 16),
2228 => conv_std_logic_vector(1440, 16),
2229 => conv_std_logic_vector(1448, 16),
2230 => conv_std_logic_vector(1456, 16),
2231 => conv_std_logic_vector(1464, 16),
2232 => conv_std_logic_vector(1472, 16),
2233 => conv_std_logic_vector(1480, 16),
2234 => conv_std_logic_vector(1488, 16),
2235 => conv_std_logic_vector(1496, 16),
2236 => conv_std_logic_vector(1504, 16),
2237 => conv_std_logic_vector(1512, 16),
2238 => conv_std_logic_vector(1520, 16),
2239 => conv_std_logic_vector(1528, 16),
2240 => conv_std_logic_vector(1536, 16),
2241 => conv_std_logic_vector(1544, 16),
2242 => conv_std_logic_vector(1552, 16),
2243 => conv_std_logic_vector(1560, 16),
2244 => conv_std_logic_vector(1568, 16),
2245 => conv_std_logic_vector(1576, 16),
2246 => conv_std_logic_vector(1584, 16),
2247 => conv_std_logic_vector(1592, 16),
2248 => conv_std_logic_vector(1600, 16),
2249 => conv_std_logic_vector(1608, 16),
2250 => conv_std_logic_vector(1616, 16),
2251 => conv_std_logic_vector(1624, 16),
2252 => conv_std_logic_vector(1632, 16),
2253 => conv_std_logic_vector(1640, 16),
2254 => conv_std_logic_vector(1648, 16),
2255 => conv_std_logic_vector(1656, 16),
2256 => conv_std_logic_vector(1664, 16),
2257 => conv_std_logic_vector(1672, 16),
2258 => conv_std_logic_vector(1680, 16),
2259 => conv_std_logic_vector(1688, 16),
2260 => conv_std_logic_vector(1696, 16),
2261 => conv_std_logic_vector(1704, 16),
2262 => conv_std_logic_vector(1712, 16),
2263 => conv_std_logic_vector(1720, 16),
2264 => conv_std_logic_vector(1728, 16),
2265 => conv_std_logic_vector(1736, 16),
2266 => conv_std_logic_vector(1744, 16),
2267 => conv_std_logic_vector(1752, 16),
2268 => conv_std_logic_vector(1760, 16),
2269 => conv_std_logic_vector(1768, 16),
2270 => conv_std_logic_vector(1776, 16),
2271 => conv_std_logic_vector(1784, 16),
2272 => conv_std_logic_vector(1792, 16),
2273 => conv_std_logic_vector(1800, 16),
2274 => conv_std_logic_vector(1808, 16),
2275 => conv_std_logic_vector(1816, 16),
2276 => conv_std_logic_vector(1824, 16),
2277 => conv_std_logic_vector(1832, 16),
2278 => conv_std_logic_vector(1840, 16),
2279 => conv_std_logic_vector(1848, 16),
2280 => conv_std_logic_vector(1856, 16),
2281 => conv_std_logic_vector(1864, 16),
2282 => conv_std_logic_vector(1872, 16),
2283 => conv_std_logic_vector(1880, 16),
2284 => conv_std_logic_vector(1888, 16),
2285 => conv_std_logic_vector(1896, 16),
2286 => conv_std_logic_vector(1904, 16),
2287 => conv_std_logic_vector(1912, 16),
2288 => conv_std_logic_vector(1920, 16),
2289 => conv_std_logic_vector(1928, 16),
2290 => conv_std_logic_vector(1936, 16),
2291 => conv_std_logic_vector(1944, 16),
2292 => conv_std_logic_vector(1952, 16),
2293 => conv_std_logic_vector(1960, 16),
2294 => conv_std_logic_vector(1968, 16),
2295 => conv_std_logic_vector(1976, 16),
2296 => conv_std_logic_vector(1984, 16),
2297 => conv_std_logic_vector(1992, 16),
2298 => conv_std_logic_vector(2000, 16),
2299 => conv_std_logic_vector(2008, 16),
2300 => conv_std_logic_vector(2016, 16),
2301 => conv_std_logic_vector(2024, 16),
2302 => conv_std_logic_vector(2032, 16),
2303 => conv_std_logic_vector(2040, 16),
2304 => conv_std_logic_vector(0, 16),
2305 => conv_std_logic_vector(9, 16),
2306 => conv_std_logic_vector(18, 16),
2307 => conv_std_logic_vector(27, 16),
2308 => conv_std_logic_vector(36, 16),
2309 => conv_std_logic_vector(45, 16),
2310 => conv_std_logic_vector(54, 16),
2311 => conv_std_logic_vector(63, 16),
2312 => conv_std_logic_vector(72, 16),
2313 => conv_std_logic_vector(81, 16),
2314 => conv_std_logic_vector(90, 16),
2315 => conv_std_logic_vector(99, 16),
2316 => conv_std_logic_vector(108, 16),
2317 => conv_std_logic_vector(117, 16),
2318 => conv_std_logic_vector(126, 16),
2319 => conv_std_logic_vector(135, 16),
2320 => conv_std_logic_vector(144, 16),
2321 => conv_std_logic_vector(153, 16),
2322 => conv_std_logic_vector(162, 16),
2323 => conv_std_logic_vector(171, 16),
2324 => conv_std_logic_vector(180, 16),
2325 => conv_std_logic_vector(189, 16),
2326 => conv_std_logic_vector(198, 16),
2327 => conv_std_logic_vector(207, 16),
2328 => conv_std_logic_vector(216, 16),
2329 => conv_std_logic_vector(225, 16),
2330 => conv_std_logic_vector(234, 16),
2331 => conv_std_logic_vector(243, 16),
2332 => conv_std_logic_vector(252, 16),
2333 => conv_std_logic_vector(261, 16),
2334 => conv_std_logic_vector(270, 16),
2335 => conv_std_logic_vector(279, 16),
2336 => conv_std_logic_vector(288, 16),
2337 => conv_std_logic_vector(297, 16),
2338 => conv_std_logic_vector(306, 16),
2339 => conv_std_logic_vector(315, 16),
2340 => conv_std_logic_vector(324, 16),
2341 => conv_std_logic_vector(333, 16),
2342 => conv_std_logic_vector(342, 16),
2343 => conv_std_logic_vector(351, 16),
2344 => conv_std_logic_vector(360, 16),
2345 => conv_std_logic_vector(369, 16),
2346 => conv_std_logic_vector(378, 16),
2347 => conv_std_logic_vector(387, 16),
2348 => conv_std_logic_vector(396, 16),
2349 => conv_std_logic_vector(405, 16),
2350 => conv_std_logic_vector(414, 16),
2351 => conv_std_logic_vector(423, 16),
2352 => conv_std_logic_vector(432, 16),
2353 => conv_std_logic_vector(441, 16),
2354 => conv_std_logic_vector(450, 16),
2355 => conv_std_logic_vector(459, 16),
2356 => conv_std_logic_vector(468, 16),
2357 => conv_std_logic_vector(477, 16),
2358 => conv_std_logic_vector(486, 16),
2359 => conv_std_logic_vector(495, 16),
2360 => conv_std_logic_vector(504, 16),
2361 => conv_std_logic_vector(513, 16),
2362 => conv_std_logic_vector(522, 16),
2363 => conv_std_logic_vector(531, 16),
2364 => conv_std_logic_vector(540, 16),
2365 => conv_std_logic_vector(549, 16),
2366 => conv_std_logic_vector(558, 16),
2367 => conv_std_logic_vector(567, 16),
2368 => conv_std_logic_vector(576, 16),
2369 => conv_std_logic_vector(585, 16),
2370 => conv_std_logic_vector(594, 16),
2371 => conv_std_logic_vector(603, 16),
2372 => conv_std_logic_vector(612, 16),
2373 => conv_std_logic_vector(621, 16),
2374 => conv_std_logic_vector(630, 16),
2375 => conv_std_logic_vector(639, 16),
2376 => conv_std_logic_vector(648, 16),
2377 => conv_std_logic_vector(657, 16),
2378 => conv_std_logic_vector(666, 16),
2379 => conv_std_logic_vector(675, 16),
2380 => conv_std_logic_vector(684, 16),
2381 => conv_std_logic_vector(693, 16),
2382 => conv_std_logic_vector(702, 16),
2383 => conv_std_logic_vector(711, 16),
2384 => conv_std_logic_vector(720, 16),
2385 => conv_std_logic_vector(729, 16),
2386 => conv_std_logic_vector(738, 16),
2387 => conv_std_logic_vector(747, 16),
2388 => conv_std_logic_vector(756, 16),
2389 => conv_std_logic_vector(765, 16),
2390 => conv_std_logic_vector(774, 16),
2391 => conv_std_logic_vector(783, 16),
2392 => conv_std_logic_vector(792, 16),
2393 => conv_std_logic_vector(801, 16),
2394 => conv_std_logic_vector(810, 16),
2395 => conv_std_logic_vector(819, 16),
2396 => conv_std_logic_vector(828, 16),
2397 => conv_std_logic_vector(837, 16),
2398 => conv_std_logic_vector(846, 16),
2399 => conv_std_logic_vector(855, 16),
2400 => conv_std_logic_vector(864, 16),
2401 => conv_std_logic_vector(873, 16),
2402 => conv_std_logic_vector(882, 16),
2403 => conv_std_logic_vector(891, 16),
2404 => conv_std_logic_vector(900, 16),
2405 => conv_std_logic_vector(909, 16),
2406 => conv_std_logic_vector(918, 16),
2407 => conv_std_logic_vector(927, 16),
2408 => conv_std_logic_vector(936, 16),
2409 => conv_std_logic_vector(945, 16),
2410 => conv_std_logic_vector(954, 16),
2411 => conv_std_logic_vector(963, 16),
2412 => conv_std_logic_vector(972, 16),
2413 => conv_std_logic_vector(981, 16),
2414 => conv_std_logic_vector(990, 16),
2415 => conv_std_logic_vector(999, 16),
2416 => conv_std_logic_vector(1008, 16),
2417 => conv_std_logic_vector(1017, 16),
2418 => conv_std_logic_vector(1026, 16),
2419 => conv_std_logic_vector(1035, 16),
2420 => conv_std_logic_vector(1044, 16),
2421 => conv_std_logic_vector(1053, 16),
2422 => conv_std_logic_vector(1062, 16),
2423 => conv_std_logic_vector(1071, 16),
2424 => conv_std_logic_vector(1080, 16),
2425 => conv_std_logic_vector(1089, 16),
2426 => conv_std_logic_vector(1098, 16),
2427 => conv_std_logic_vector(1107, 16),
2428 => conv_std_logic_vector(1116, 16),
2429 => conv_std_logic_vector(1125, 16),
2430 => conv_std_logic_vector(1134, 16),
2431 => conv_std_logic_vector(1143, 16),
2432 => conv_std_logic_vector(1152, 16),
2433 => conv_std_logic_vector(1161, 16),
2434 => conv_std_logic_vector(1170, 16),
2435 => conv_std_logic_vector(1179, 16),
2436 => conv_std_logic_vector(1188, 16),
2437 => conv_std_logic_vector(1197, 16),
2438 => conv_std_logic_vector(1206, 16),
2439 => conv_std_logic_vector(1215, 16),
2440 => conv_std_logic_vector(1224, 16),
2441 => conv_std_logic_vector(1233, 16),
2442 => conv_std_logic_vector(1242, 16),
2443 => conv_std_logic_vector(1251, 16),
2444 => conv_std_logic_vector(1260, 16),
2445 => conv_std_logic_vector(1269, 16),
2446 => conv_std_logic_vector(1278, 16),
2447 => conv_std_logic_vector(1287, 16),
2448 => conv_std_logic_vector(1296, 16),
2449 => conv_std_logic_vector(1305, 16),
2450 => conv_std_logic_vector(1314, 16),
2451 => conv_std_logic_vector(1323, 16),
2452 => conv_std_logic_vector(1332, 16),
2453 => conv_std_logic_vector(1341, 16),
2454 => conv_std_logic_vector(1350, 16),
2455 => conv_std_logic_vector(1359, 16),
2456 => conv_std_logic_vector(1368, 16),
2457 => conv_std_logic_vector(1377, 16),
2458 => conv_std_logic_vector(1386, 16),
2459 => conv_std_logic_vector(1395, 16),
2460 => conv_std_logic_vector(1404, 16),
2461 => conv_std_logic_vector(1413, 16),
2462 => conv_std_logic_vector(1422, 16),
2463 => conv_std_logic_vector(1431, 16),
2464 => conv_std_logic_vector(1440, 16),
2465 => conv_std_logic_vector(1449, 16),
2466 => conv_std_logic_vector(1458, 16),
2467 => conv_std_logic_vector(1467, 16),
2468 => conv_std_logic_vector(1476, 16),
2469 => conv_std_logic_vector(1485, 16),
2470 => conv_std_logic_vector(1494, 16),
2471 => conv_std_logic_vector(1503, 16),
2472 => conv_std_logic_vector(1512, 16),
2473 => conv_std_logic_vector(1521, 16),
2474 => conv_std_logic_vector(1530, 16),
2475 => conv_std_logic_vector(1539, 16),
2476 => conv_std_logic_vector(1548, 16),
2477 => conv_std_logic_vector(1557, 16),
2478 => conv_std_logic_vector(1566, 16),
2479 => conv_std_logic_vector(1575, 16),
2480 => conv_std_logic_vector(1584, 16),
2481 => conv_std_logic_vector(1593, 16),
2482 => conv_std_logic_vector(1602, 16),
2483 => conv_std_logic_vector(1611, 16),
2484 => conv_std_logic_vector(1620, 16),
2485 => conv_std_logic_vector(1629, 16),
2486 => conv_std_logic_vector(1638, 16),
2487 => conv_std_logic_vector(1647, 16),
2488 => conv_std_logic_vector(1656, 16),
2489 => conv_std_logic_vector(1665, 16),
2490 => conv_std_logic_vector(1674, 16),
2491 => conv_std_logic_vector(1683, 16),
2492 => conv_std_logic_vector(1692, 16),
2493 => conv_std_logic_vector(1701, 16),
2494 => conv_std_logic_vector(1710, 16),
2495 => conv_std_logic_vector(1719, 16),
2496 => conv_std_logic_vector(1728, 16),
2497 => conv_std_logic_vector(1737, 16),
2498 => conv_std_logic_vector(1746, 16),
2499 => conv_std_logic_vector(1755, 16),
2500 => conv_std_logic_vector(1764, 16),
2501 => conv_std_logic_vector(1773, 16),
2502 => conv_std_logic_vector(1782, 16),
2503 => conv_std_logic_vector(1791, 16),
2504 => conv_std_logic_vector(1800, 16),
2505 => conv_std_logic_vector(1809, 16),
2506 => conv_std_logic_vector(1818, 16),
2507 => conv_std_logic_vector(1827, 16),
2508 => conv_std_logic_vector(1836, 16),
2509 => conv_std_logic_vector(1845, 16),
2510 => conv_std_logic_vector(1854, 16),
2511 => conv_std_logic_vector(1863, 16),
2512 => conv_std_logic_vector(1872, 16),
2513 => conv_std_logic_vector(1881, 16),
2514 => conv_std_logic_vector(1890, 16),
2515 => conv_std_logic_vector(1899, 16),
2516 => conv_std_logic_vector(1908, 16),
2517 => conv_std_logic_vector(1917, 16),
2518 => conv_std_logic_vector(1926, 16),
2519 => conv_std_logic_vector(1935, 16),
2520 => conv_std_logic_vector(1944, 16),
2521 => conv_std_logic_vector(1953, 16),
2522 => conv_std_logic_vector(1962, 16),
2523 => conv_std_logic_vector(1971, 16),
2524 => conv_std_logic_vector(1980, 16),
2525 => conv_std_logic_vector(1989, 16),
2526 => conv_std_logic_vector(1998, 16),
2527 => conv_std_logic_vector(2007, 16),
2528 => conv_std_logic_vector(2016, 16),
2529 => conv_std_logic_vector(2025, 16),
2530 => conv_std_logic_vector(2034, 16),
2531 => conv_std_logic_vector(2043, 16),
2532 => conv_std_logic_vector(2052, 16),
2533 => conv_std_logic_vector(2061, 16),
2534 => conv_std_logic_vector(2070, 16),
2535 => conv_std_logic_vector(2079, 16),
2536 => conv_std_logic_vector(2088, 16),
2537 => conv_std_logic_vector(2097, 16),
2538 => conv_std_logic_vector(2106, 16),
2539 => conv_std_logic_vector(2115, 16),
2540 => conv_std_logic_vector(2124, 16),
2541 => conv_std_logic_vector(2133, 16),
2542 => conv_std_logic_vector(2142, 16),
2543 => conv_std_logic_vector(2151, 16),
2544 => conv_std_logic_vector(2160, 16),
2545 => conv_std_logic_vector(2169, 16),
2546 => conv_std_logic_vector(2178, 16),
2547 => conv_std_logic_vector(2187, 16),
2548 => conv_std_logic_vector(2196, 16),
2549 => conv_std_logic_vector(2205, 16),
2550 => conv_std_logic_vector(2214, 16),
2551 => conv_std_logic_vector(2223, 16),
2552 => conv_std_logic_vector(2232, 16),
2553 => conv_std_logic_vector(2241, 16),
2554 => conv_std_logic_vector(2250, 16),
2555 => conv_std_logic_vector(2259, 16),
2556 => conv_std_logic_vector(2268, 16),
2557 => conv_std_logic_vector(2277, 16),
2558 => conv_std_logic_vector(2286, 16),
2559 => conv_std_logic_vector(2295, 16),
2560 => conv_std_logic_vector(0, 16),
2561 => conv_std_logic_vector(10, 16),
2562 => conv_std_logic_vector(20, 16),
2563 => conv_std_logic_vector(30, 16),
2564 => conv_std_logic_vector(40, 16),
2565 => conv_std_logic_vector(50, 16),
2566 => conv_std_logic_vector(60, 16),
2567 => conv_std_logic_vector(70, 16),
2568 => conv_std_logic_vector(80, 16),
2569 => conv_std_logic_vector(90, 16),
2570 => conv_std_logic_vector(100, 16),
2571 => conv_std_logic_vector(110, 16),
2572 => conv_std_logic_vector(120, 16),
2573 => conv_std_logic_vector(130, 16),
2574 => conv_std_logic_vector(140, 16),
2575 => conv_std_logic_vector(150, 16),
2576 => conv_std_logic_vector(160, 16),
2577 => conv_std_logic_vector(170, 16),
2578 => conv_std_logic_vector(180, 16),
2579 => conv_std_logic_vector(190, 16),
2580 => conv_std_logic_vector(200, 16),
2581 => conv_std_logic_vector(210, 16),
2582 => conv_std_logic_vector(220, 16),
2583 => conv_std_logic_vector(230, 16),
2584 => conv_std_logic_vector(240, 16),
2585 => conv_std_logic_vector(250, 16),
2586 => conv_std_logic_vector(260, 16),
2587 => conv_std_logic_vector(270, 16),
2588 => conv_std_logic_vector(280, 16),
2589 => conv_std_logic_vector(290, 16),
2590 => conv_std_logic_vector(300, 16),
2591 => conv_std_logic_vector(310, 16),
2592 => conv_std_logic_vector(320, 16),
2593 => conv_std_logic_vector(330, 16),
2594 => conv_std_logic_vector(340, 16),
2595 => conv_std_logic_vector(350, 16),
2596 => conv_std_logic_vector(360, 16),
2597 => conv_std_logic_vector(370, 16),
2598 => conv_std_logic_vector(380, 16),
2599 => conv_std_logic_vector(390, 16),
2600 => conv_std_logic_vector(400, 16),
2601 => conv_std_logic_vector(410, 16),
2602 => conv_std_logic_vector(420, 16),
2603 => conv_std_logic_vector(430, 16),
2604 => conv_std_logic_vector(440, 16),
2605 => conv_std_logic_vector(450, 16),
2606 => conv_std_logic_vector(460, 16),
2607 => conv_std_logic_vector(470, 16),
2608 => conv_std_logic_vector(480, 16),
2609 => conv_std_logic_vector(490, 16),
2610 => conv_std_logic_vector(500, 16),
2611 => conv_std_logic_vector(510, 16),
2612 => conv_std_logic_vector(520, 16),
2613 => conv_std_logic_vector(530, 16),
2614 => conv_std_logic_vector(540, 16),
2615 => conv_std_logic_vector(550, 16),
2616 => conv_std_logic_vector(560, 16),
2617 => conv_std_logic_vector(570, 16),
2618 => conv_std_logic_vector(580, 16),
2619 => conv_std_logic_vector(590, 16),
2620 => conv_std_logic_vector(600, 16),
2621 => conv_std_logic_vector(610, 16),
2622 => conv_std_logic_vector(620, 16),
2623 => conv_std_logic_vector(630, 16),
2624 => conv_std_logic_vector(640, 16),
2625 => conv_std_logic_vector(650, 16),
2626 => conv_std_logic_vector(660, 16),
2627 => conv_std_logic_vector(670, 16),
2628 => conv_std_logic_vector(680, 16),
2629 => conv_std_logic_vector(690, 16),
2630 => conv_std_logic_vector(700, 16),
2631 => conv_std_logic_vector(710, 16),
2632 => conv_std_logic_vector(720, 16),
2633 => conv_std_logic_vector(730, 16),
2634 => conv_std_logic_vector(740, 16),
2635 => conv_std_logic_vector(750, 16),
2636 => conv_std_logic_vector(760, 16),
2637 => conv_std_logic_vector(770, 16),
2638 => conv_std_logic_vector(780, 16),
2639 => conv_std_logic_vector(790, 16),
2640 => conv_std_logic_vector(800, 16),
2641 => conv_std_logic_vector(810, 16),
2642 => conv_std_logic_vector(820, 16),
2643 => conv_std_logic_vector(830, 16),
2644 => conv_std_logic_vector(840, 16),
2645 => conv_std_logic_vector(850, 16),
2646 => conv_std_logic_vector(860, 16),
2647 => conv_std_logic_vector(870, 16),
2648 => conv_std_logic_vector(880, 16),
2649 => conv_std_logic_vector(890, 16),
2650 => conv_std_logic_vector(900, 16),
2651 => conv_std_logic_vector(910, 16),
2652 => conv_std_logic_vector(920, 16),
2653 => conv_std_logic_vector(930, 16),
2654 => conv_std_logic_vector(940, 16),
2655 => conv_std_logic_vector(950, 16),
2656 => conv_std_logic_vector(960, 16),
2657 => conv_std_logic_vector(970, 16),
2658 => conv_std_logic_vector(980, 16),
2659 => conv_std_logic_vector(990, 16),
2660 => conv_std_logic_vector(1000, 16),
2661 => conv_std_logic_vector(1010, 16),
2662 => conv_std_logic_vector(1020, 16),
2663 => conv_std_logic_vector(1030, 16),
2664 => conv_std_logic_vector(1040, 16),
2665 => conv_std_logic_vector(1050, 16),
2666 => conv_std_logic_vector(1060, 16),
2667 => conv_std_logic_vector(1070, 16),
2668 => conv_std_logic_vector(1080, 16),
2669 => conv_std_logic_vector(1090, 16),
2670 => conv_std_logic_vector(1100, 16),
2671 => conv_std_logic_vector(1110, 16),
2672 => conv_std_logic_vector(1120, 16),
2673 => conv_std_logic_vector(1130, 16),
2674 => conv_std_logic_vector(1140, 16),
2675 => conv_std_logic_vector(1150, 16),
2676 => conv_std_logic_vector(1160, 16),
2677 => conv_std_logic_vector(1170, 16),
2678 => conv_std_logic_vector(1180, 16),
2679 => conv_std_logic_vector(1190, 16),
2680 => conv_std_logic_vector(1200, 16),
2681 => conv_std_logic_vector(1210, 16),
2682 => conv_std_logic_vector(1220, 16),
2683 => conv_std_logic_vector(1230, 16),
2684 => conv_std_logic_vector(1240, 16),
2685 => conv_std_logic_vector(1250, 16),
2686 => conv_std_logic_vector(1260, 16),
2687 => conv_std_logic_vector(1270, 16),
2688 => conv_std_logic_vector(1280, 16),
2689 => conv_std_logic_vector(1290, 16),
2690 => conv_std_logic_vector(1300, 16),
2691 => conv_std_logic_vector(1310, 16),
2692 => conv_std_logic_vector(1320, 16),
2693 => conv_std_logic_vector(1330, 16),
2694 => conv_std_logic_vector(1340, 16),
2695 => conv_std_logic_vector(1350, 16),
2696 => conv_std_logic_vector(1360, 16),
2697 => conv_std_logic_vector(1370, 16),
2698 => conv_std_logic_vector(1380, 16),
2699 => conv_std_logic_vector(1390, 16),
2700 => conv_std_logic_vector(1400, 16),
2701 => conv_std_logic_vector(1410, 16),
2702 => conv_std_logic_vector(1420, 16),
2703 => conv_std_logic_vector(1430, 16),
2704 => conv_std_logic_vector(1440, 16),
2705 => conv_std_logic_vector(1450, 16),
2706 => conv_std_logic_vector(1460, 16),
2707 => conv_std_logic_vector(1470, 16),
2708 => conv_std_logic_vector(1480, 16),
2709 => conv_std_logic_vector(1490, 16),
2710 => conv_std_logic_vector(1500, 16),
2711 => conv_std_logic_vector(1510, 16),
2712 => conv_std_logic_vector(1520, 16),
2713 => conv_std_logic_vector(1530, 16),
2714 => conv_std_logic_vector(1540, 16),
2715 => conv_std_logic_vector(1550, 16),
2716 => conv_std_logic_vector(1560, 16),
2717 => conv_std_logic_vector(1570, 16),
2718 => conv_std_logic_vector(1580, 16),
2719 => conv_std_logic_vector(1590, 16),
2720 => conv_std_logic_vector(1600, 16),
2721 => conv_std_logic_vector(1610, 16),
2722 => conv_std_logic_vector(1620, 16),
2723 => conv_std_logic_vector(1630, 16),
2724 => conv_std_logic_vector(1640, 16),
2725 => conv_std_logic_vector(1650, 16),
2726 => conv_std_logic_vector(1660, 16),
2727 => conv_std_logic_vector(1670, 16),
2728 => conv_std_logic_vector(1680, 16),
2729 => conv_std_logic_vector(1690, 16),
2730 => conv_std_logic_vector(1700, 16),
2731 => conv_std_logic_vector(1710, 16),
2732 => conv_std_logic_vector(1720, 16),
2733 => conv_std_logic_vector(1730, 16),
2734 => conv_std_logic_vector(1740, 16),
2735 => conv_std_logic_vector(1750, 16),
2736 => conv_std_logic_vector(1760, 16),
2737 => conv_std_logic_vector(1770, 16),
2738 => conv_std_logic_vector(1780, 16),
2739 => conv_std_logic_vector(1790, 16),
2740 => conv_std_logic_vector(1800, 16),
2741 => conv_std_logic_vector(1810, 16),
2742 => conv_std_logic_vector(1820, 16),
2743 => conv_std_logic_vector(1830, 16),
2744 => conv_std_logic_vector(1840, 16),
2745 => conv_std_logic_vector(1850, 16),
2746 => conv_std_logic_vector(1860, 16),
2747 => conv_std_logic_vector(1870, 16),
2748 => conv_std_logic_vector(1880, 16),
2749 => conv_std_logic_vector(1890, 16),
2750 => conv_std_logic_vector(1900, 16),
2751 => conv_std_logic_vector(1910, 16),
2752 => conv_std_logic_vector(1920, 16),
2753 => conv_std_logic_vector(1930, 16),
2754 => conv_std_logic_vector(1940, 16),
2755 => conv_std_logic_vector(1950, 16),
2756 => conv_std_logic_vector(1960, 16),
2757 => conv_std_logic_vector(1970, 16),
2758 => conv_std_logic_vector(1980, 16),
2759 => conv_std_logic_vector(1990, 16),
2760 => conv_std_logic_vector(2000, 16),
2761 => conv_std_logic_vector(2010, 16),
2762 => conv_std_logic_vector(2020, 16),
2763 => conv_std_logic_vector(2030, 16),
2764 => conv_std_logic_vector(2040, 16),
2765 => conv_std_logic_vector(2050, 16),
2766 => conv_std_logic_vector(2060, 16),
2767 => conv_std_logic_vector(2070, 16),
2768 => conv_std_logic_vector(2080, 16),
2769 => conv_std_logic_vector(2090, 16),
2770 => conv_std_logic_vector(2100, 16),
2771 => conv_std_logic_vector(2110, 16),
2772 => conv_std_logic_vector(2120, 16),
2773 => conv_std_logic_vector(2130, 16),
2774 => conv_std_logic_vector(2140, 16),
2775 => conv_std_logic_vector(2150, 16),
2776 => conv_std_logic_vector(2160, 16),
2777 => conv_std_logic_vector(2170, 16),
2778 => conv_std_logic_vector(2180, 16),
2779 => conv_std_logic_vector(2190, 16),
2780 => conv_std_logic_vector(2200, 16),
2781 => conv_std_logic_vector(2210, 16),
2782 => conv_std_logic_vector(2220, 16),
2783 => conv_std_logic_vector(2230, 16),
2784 => conv_std_logic_vector(2240, 16),
2785 => conv_std_logic_vector(2250, 16),
2786 => conv_std_logic_vector(2260, 16),
2787 => conv_std_logic_vector(2270, 16),
2788 => conv_std_logic_vector(2280, 16),
2789 => conv_std_logic_vector(2290, 16),
2790 => conv_std_logic_vector(2300, 16),
2791 => conv_std_logic_vector(2310, 16),
2792 => conv_std_logic_vector(2320, 16),
2793 => conv_std_logic_vector(2330, 16),
2794 => conv_std_logic_vector(2340, 16),
2795 => conv_std_logic_vector(2350, 16),
2796 => conv_std_logic_vector(2360, 16),
2797 => conv_std_logic_vector(2370, 16),
2798 => conv_std_logic_vector(2380, 16),
2799 => conv_std_logic_vector(2390, 16),
2800 => conv_std_logic_vector(2400, 16),
2801 => conv_std_logic_vector(2410, 16),
2802 => conv_std_logic_vector(2420, 16),
2803 => conv_std_logic_vector(2430, 16),
2804 => conv_std_logic_vector(2440, 16),
2805 => conv_std_logic_vector(2450, 16),
2806 => conv_std_logic_vector(2460, 16),
2807 => conv_std_logic_vector(2470, 16),
2808 => conv_std_logic_vector(2480, 16),
2809 => conv_std_logic_vector(2490, 16),
2810 => conv_std_logic_vector(2500, 16),
2811 => conv_std_logic_vector(2510, 16),
2812 => conv_std_logic_vector(2520, 16),
2813 => conv_std_logic_vector(2530, 16),
2814 => conv_std_logic_vector(2540, 16),
2815 => conv_std_logic_vector(2550, 16),
2816 => conv_std_logic_vector(0, 16),
2817 => conv_std_logic_vector(11, 16),
2818 => conv_std_logic_vector(22, 16),
2819 => conv_std_logic_vector(33, 16),
2820 => conv_std_logic_vector(44, 16),
2821 => conv_std_logic_vector(55, 16),
2822 => conv_std_logic_vector(66, 16),
2823 => conv_std_logic_vector(77, 16),
2824 => conv_std_logic_vector(88, 16),
2825 => conv_std_logic_vector(99, 16),
2826 => conv_std_logic_vector(110, 16),
2827 => conv_std_logic_vector(121, 16),
2828 => conv_std_logic_vector(132, 16),
2829 => conv_std_logic_vector(143, 16),
2830 => conv_std_logic_vector(154, 16),
2831 => conv_std_logic_vector(165, 16),
2832 => conv_std_logic_vector(176, 16),
2833 => conv_std_logic_vector(187, 16),
2834 => conv_std_logic_vector(198, 16),
2835 => conv_std_logic_vector(209, 16),
2836 => conv_std_logic_vector(220, 16),
2837 => conv_std_logic_vector(231, 16),
2838 => conv_std_logic_vector(242, 16),
2839 => conv_std_logic_vector(253, 16),
2840 => conv_std_logic_vector(264, 16),
2841 => conv_std_logic_vector(275, 16),
2842 => conv_std_logic_vector(286, 16),
2843 => conv_std_logic_vector(297, 16),
2844 => conv_std_logic_vector(308, 16),
2845 => conv_std_logic_vector(319, 16),
2846 => conv_std_logic_vector(330, 16),
2847 => conv_std_logic_vector(341, 16),
2848 => conv_std_logic_vector(352, 16),
2849 => conv_std_logic_vector(363, 16),
2850 => conv_std_logic_vector(374, 16),
2851 => conv_std_logic_vector(385, 16),
2852 => conv_std_logic_vector(396, 16),
2853 => conv_std_logic_vector(407, 16),
2854 => conv_std_logic_vector(418, 16),
2855 => conv_std_logic_vector(429, 16),
2856 => conv_std_logic_vector(440, 16),
2857 => conv_std_logic_vector(451, 16),
2858 => conv_std_logic_vector(462, 16),
2859 => conv_std_logic_vector(473, 16),
2860 => conv_std_logic_vector(484, 16),
2861 => conv_std_logic_vector(495, 16),
2862 => conv_std_logic_vector(506, 16),
2863 => conv_std_logic_vector(517, 16),
2864 => conv_std_logic_vector(528, 16),
2865 => conv_std_logic_vector(539, 16),
2866 => conv_std_logic_vector(550, 16),
2867 => conv_std_logic_vector(561, 16),
2868 => conv_std_logic_vector(572, 16),
2869 => conv_std_logic_vector(583, 16),
2870 => conv_std_logic_vector(594, 16),
2871 => conv_std_logic_vector(605, 16),
2872 => conv_std_logic_vector(616, 16),
2873 => conv_std_logic_vector(627, 16),
2874 => conv_std_logic_vector(638, 16),
2875 => conv_std_logic_vector(649, 16),
2876 => conv_std_logic_vector(660, 16),
2877 => conv_std_logic_vector(671, 16),
2878 => conv_std_logic_vector(682, 16),
2879 => conv_std_logic_vector(693, 16),
2880 => conv_std_logic_vector(704, 16),
2881 => conv_std_logic_vector(715, 16),
2882 => conv_std_logic_vector(726, 16),
2883 => conv_std_logic_vector(737, 16),
2884 => conv_std_logic_vector(748, 16),
2885 => conv_std_logic_vector(759, 16),
2886 => conv_std_logic_vector(770, 16),
2887 => conv_std_logic_vector(781, 16),
2888 => conv_std_logic_vector(792, 16),
2889 => conv_std_logic_vector(803, 16),
2890 => conv_std_logic_vector(814, 16),
2891 => conv_std_logic_vector(825, 16),
2892 => conv_std_logic_vector(836, 16),
2893 => conv_std_logic_vector(847, 16),
2894 => conv_std_logic_vector(858, 16),
2895 => conv_std_logic_vector(869, 16),
2896 => conv_std_logic_vector(880, 16),
2897 => conv_std_logic_vector(891, 16),
2898 => conv_std_logic_vector(902, 16),
2899 => conv_std_logic_vector(913, 16),
2900 => conv_std_logic_vector(924, 16),
2901 => conv_std_logic_vector(935, 16),
2902 => conv_std_logic_vector(946, 16),
2903 => conv_std_logic_vector(957, 16),
2904 => conv_std_logic_vector(968, 16),
2905 => conv_std_logic_vector(979, 16),
2906 => conv_std_logic_vector(990, 16),
2907 => conv_std_logic_vector(1001, 16),
2908 => conv_std_logic_vector(1012, 16),
2909 => conv_std_logic_vector(1023, 16),
2910 => conv_std_logic_vector(1034, 16),
2911 => conv_std_logic_vector(1045, 16),
2912 => conv_std_logic_vector(1056, 16),
2913 => conv_std_logic_vector(1067, 16),
2914 => conv_std_logic_vector(1078, 16),
2915 => conv_std_logic_vector(1089, 16),
2916 => conv_std_logic_vector(1100, 16),
2917 => conv_std_logic_vector(1111, 16),
2918 => conv_std_logic_vector(1122, 16),
2919 => conv_std_logic_vector(1133, 16),
2920 => conv_std_logic_vector(1144, 16),
2921 => conv_std_logic_vector(1155, 16),
2922 => conv_std_logic_vector(1166, 16),
2923 => conv_std_logic_vector(1177, 16),
2924 => conv_std_logic_vector(1188, 16),
2925 => conv_std_logic_vector(1199, 16),
2926 => conv_std_logic_vector(1210, 16),
2927 => conv_std_logic_vector(1221, 16),
2928 => conv_std_logic_vector(1232, 16),
2929 => conv_std_logic_vector(1243, 16),
2930 => conv_std_logic_vector(1254, 16),
2931 => conv_std_logic_vector(1265, 16),
2932 => conv_std_logic_vector(1276, 16),
2933 => conv_std_logic_vector(1287, 16),
2934 => conv_std_logic_vector(1298, 16),
2935 => conv_std_logic_vector(1309, 16),
2936 => conv_std_logic_vector(1320, 16),
2937 => conv_std_logic_vector(1331, 16),
2938 => conv_std_logic_vector(1342, 16),
2939 => conv_std_logic_vector(1353, 16),
2940 => conv_std_logic_vector(1364, 16),
2941 => conv_std_logic_vector(1375, 16),
2942 => conv_std_logic_vector(1386, 16),
2943 => conv_std_logic_vector(1397, 16),
2944 => conv_std_logic_vector(1408, 16),
2945 => conv_std_logic_vector(1419, 16),
2946 => conv_std_logic_vector(1430, 16),
2947 => conv_std_logic_vector(1441, 16),
2948 => conv_std_logic_vector(1452, 16),
2949 => conv_std_logic_vector(1463, 16),
2950 => conv_std_logic_vector(1474, 16),
2951 => conv_std_logic_vector(1485, 16),
2952 => conv_std_logic_vector(1496, 16),
2953 => conv_std_logic_vector(1507, 16),
2954 => conv_std_logic_vector(1518, 16),
2955 => conv_std_logic_vector(1529, 16),
2956 => conv_std_logic_vector(1540, 16),
2957 => conv_std_logic_vector(1551, 16),
2958 => conv_std_logic_vector(1562, 16),
2959 => conv_std_logic_vector(1573, 16),
2960 => conv_std_logic_vector(1584, 16),
2961 => conv_std_logic_vector(1595, 16),
2962 => conv_std_logic_vector(1606, 16),
2963 => conv_std_logic_vector(1617, 16),
2964 => conv_std_logic_vector(1628, 16),
2965 => conv_std_logic_vector(1639, 16),
2966 => conv_std_logic_vector(1650, 16),
2967 => conv_std_logic_vector(1661, 16),
2968 => conv_std_logic_vector(1672, 16),
2969 => conv_std_logic_vector(1683, 16),
2970 => conv_std_logic_vector(1694, 16),
2971 => conv_std_logic_vector(1705, 16),
2972 => conv_std_logic_vector(1716, 16),
2973 => conv_std_logic_vector(1727, 16),
2974 => conv_std_logic_vector(1738, 16),
2975 => conv_std_logic_vector(1749, 16),
2976 => conv_std_logic_vector(1760, 16),
2977 => conv_std_logic_vector(1771, 16),
2978 => conv_std_logic_vector(1782, 16),
2979 => conv_std_logic_vector(1793, 16),
2980 => conv_std_logic_vector(1804, 16),
2981 => conv_std_logic_vector(1815, 16),
2982 => conv_std_logic_vector(1826, 16),
2983 => conv_std_logic_vector(1837, 16),
2984 => conv_std_logic_vector(1848, 16),
2985 => conv_std_logic_vector(1859, 16),
2986 => conv_std_logic_vector(1870, 16),
2987 => conv_std_logic_vector(1881, 16),
2988 => conv_std_logic_vector(1892, 16),
2989 => conv_std_logic_vector(1903, 16),
2990 => conv_std_logic_vector(1914, 16),
2991 => conv_std_logic_vector(1925, 16),
2992 => conv_std_logic_vector(1936, 16),
2993 => conv_std_logic_vector(1947, 16),
2994 => conv_std_logic_vector(1958, 16),
2995 => conv_std_logic_vector(1969, 16),
2996 => conv_std_logic_vector(1980, 16),
2997 => conv_std_logic_vector(1991, 16),
2998 => conv_std_logic_vector(2002, 16),
2999 => conv_std_logic_vector(2013, 16),
3000 => conv_std_logic_vector(2024, 16),
3001 => conv_std_logic_vector(2035, 16),
3002 => conv_std_logic_vector(2046, 16),
3003 => conv_std_logic_vector(2057, 16),
3004 => conv_std_logic_vector(2068, 16),
3005 => conv_std_logic_vector(2079, 16),
3006 => conv_std_logic_vector(2090, 16),
3007 => conv_std_logic_vector(2101, 16),
3008 => conv_std_logic_vector(2112, 16),
3009 => conv_std_logic_vector(2123, 16),
3010 => conv_std_logic_vector(2134, 16),
3011 => conv_std_logic_vector(2145, 16),
3012 => conv_std_logic_vector(2156, 16),
3013 => conv_std_logic_vector(2167, 16),
3014 => conv_std_logic_vector(2178, 16),
3015 => conv_std_logic_vector(2189, 16),
3016 => conv_std_logic_vector(2200, 16),
3017 => conv_std_logic_vector(2211, 16),
3018 => conv_std_logic_vector(2222, 16),
3019 => conv_std_logic_vector(2233, 16),
3020 => conv_std_logic_vector(2244, 16),
3021 => conv_std_logic_vector(2255, 16),
3022 => conv_std_logic_vector(2266, 16),
3023 => conv_std_logic_vector(2277, 16),
3024 => conv_std_logic_vector(2288, 16),
3025 => conv_std_logic_vector(2299, 16),
3026 => conv_std_logic_vector(2310, 16),
3027 => conv_std_logic_vector(2321, 16),
3028 => conv_std_logic_vector(2332, 16),
3029 => conv_std_logic_vector(2343, 16),
3030 => conv_std_logic_vector(2354, 16),
3031 => conv_std_logic_vector(2365, 16),
3032 => conv_std_logic_vector(2376, 16),
3033 => conv_std_logic_vector(2387, 16),
3034 => conv_std_logic_vector(2398, 16),
3035 => conv_std_logic_vector(2409, 16),
3036 => conv_std_logic_vector(2420, 16),
3037 => conv_std_logic_vector(2431, 16),
3038 => conv_std_logic_vector(2442, 16),
3039 => conv_std_logic_vector(2453, 16),
3040 => conv_std_logic_vector(2464, 16),
3041 => conv_std_logic_vector(2475, 16),
3042 => conv_std_logic_vector(2486, 16),
3043 => conv_std_logic_vector(2497, 16),
3044 => conv_std_logic_vector(2508, 16),
3045 => conv_std_logic_vector(2519, 16),
3046 => conv_std_logic_vector(2530, 16),
3047 => conv_std_logic_vector(2541, 16),
3048 => conv_std_logic_vector(2552, 16),
3049 => conv_std_logic_vector(2563, 16),
3050 => conv_std_logic_vector(2574, 16),
3051 => conv_std_logic_vector(2585, 16),
3052 => conv_std_logic_vector(2596, 16),
3053 => conv_std_logic_vector(2607, 16),
3054 => conv_std_logic_vector(2618, 16),
3055 => conv_std_logic_vector(2629, 16),
3056 => conv_std_logic_vector(2640, 16),
3057 => conv_std_logic_vector(2651, 16),
3058 => conv_std_logic_vector(2662, 16),
3059 => conv_std_logic_vector(2673, 16),
3060 => conv_std_logic_vector(2684, 16),
3061 => conv_std_logic_vector(2695, 16),
3062 => conv_std_logic_vector(2706, 16),
3063 => conv_std_logic_vector(2717, 16),
3064 => conv_std_logic_vector(2728, 16),
3065 => conv_std_logic_vector(2739, 16),
3066 => conv_std_logic_vector(2750, 16),
3067 => conv_std_logic_vector(2761, 16),
3068 => conv_std_logic_vector(2772, 16),
3069 => conv_std_logic_vector(2783, 16),
3070 => conv_std_logic_vector(2794, 16),
3071 => conv_std_logic_vector(2805, 16),
3072 => conv_std_logic_vector(0, 16),
3073 => conv_std_logic_vector(12, 16),
3074 => conv_std_logic_vector(24, 16),
3075 => conv_std_logic_vector(36, 16),
3076 => conv_std_logic_vector(48, 16),
3077 => conv_std_logic_vector(60, 16),
3078 => conv_std_logic_vector(72, 16),
3079 => conv_std_logic_vector(84, 16),
3080 => conv_std_logic_vector(96, 16),
3081 => conv_std_logic_vector(108, 16),
3082 => conv_std_logic_vector(120, 16),
3083 => conv_std_logic_vector(132, 16),
3084 => conv_std_logic_vector(144, 16),
3085 => conv_std_logic_vector(156, 16),
3086 => conv_std_logic_vector(168, 16),
3087 => conv_std_logic_vector(180, 16),
3088 => conv_std_logic_vector(192, 16),
3089 => conv_std_logic_vector(204, 16),
3090 => conv_std_logic_vector(216, 16),
3091 => conv_std_logic_vector(228, 16),
3092 => conv_std_logic_vector(240, 16),
3093 => conv_std_logic_vector(252, 16),
3094 => conv_std_logic_vector(264, 16),
3095 => conv_std_logic_vector(276, 16),
3096 => conv_std_logic_vector(288, 16),
3097 => conv_std_logic_vector(300, 16),
3098 => conv_std_logic_vector(312, 16),
3099 => conv_std_logic_vector(324, 16),
3100 => conv_std_logic_vector(336, 16),
3101 => conv_std_logic_vector(348, 16),
3102 => conv_std_logic_vector(360, 16),
3103 => conv_std_logic_vector(372, 16),
3104 => conv_std_logic_vector(384, 16),
3105 => conv_std_logic_vector(396, 16),
3106 => conv_std_logic_vector(408, 16),
3107 => conv_std_logic_vector(420, 16),
3108 => conv_std_logic_vector(432, 16),
3109 => conv_std_logic_vector(444, 16),
3110 => conv_std_logic_vector(456, 16),
3111 => conv_std_logic_vector(468, 16),
3112 => conv_std_logic_vector(480, 16),
3113 => conv_std_logic_vector(492, 16),
3114 => conv_std_logic_vector(504, 16),
3115 => conv_std_logic_vector(516, 16),
3116 => conv_std_logic_vector(528, 16),
3117 => conv_std_logic_vector(540, 16),
3118 => conv_std_logic_vector(552, 16),
3119 => conv_std_logic_vector(564, 16),
3120 => conv_std_logic_vector(576, 16),
3121 => conv_std_logic_vector(588, 16),
3122 => conv_std_logic_vector(600, 16),
3123 => conv_std_logic_vector(612, 16),
3124 => conv_std_logic_vector(624, 16),
3125 => conv_std_logic_vector(636, 16),
3126 => conv_std_logic_vector(648, 16),
3127 => conv_std_logic_vector(660, 16),
3128 => conv_std_logic_vector(672, 16),
3129 => conv_std_logic_vector(684, 16),
3130 => conv_std_logic_vector(696, 16),
3131 => conv_std_logic_vector(708, 16),
3132 => conv_std_logic_vector(720, 16),
3133 => conv_std_logic_vector(732, 16),
3134 => conv_std_logic_vector(744, 16),
3135 => conv_std_logic_vector(756, 16),
3136 => conv_std_logic_vector(768, 16),
3137 => conv_std_logic_vector(780, 16),
3138 => conv_std_logic_vector(792, 16),
3139 => conv_std_logic_vector(804, 16),
3140 => conv_std_logic_vector(816, 16),
3141 => conv_std_logic_vector(828, 16),
3142 => conv_std_logic_vector(840, 16),
3143 => conv_std_logic_vector(852, 16),
3144 => conv_std_logic_vector(864, 16),
3145 => conv_std_logic_vector(876, 16),
3146 => conv_std_logic_vector(888, 16),
3147 => conv_std_logic_vector(900, 16),
3148 => conv_std_logic_vector(912, 16),
3149 => conv_std_logic_vector(924, 16),
3150 => conv_std_logic_vector(936, 16),
3151 => conv_std_logic_vector(948, 16),
3152 => conv_std_logic_vector(960, 16),
3153 => conv_std_logic_vector(972, 16),
3154 => conv_std_logic_vector(984, 16),
3155 => conv_std_logic_vector(996, 16),
3156 => conv_std_logic_vector(1008, 16),
3157 => conv_std_logic_vector(1020, 16),
3158 => conv_std_logic_vector(1032, 16),
3159 => conv_std_logic_vector(1044, 16),
3160 => conv_std_logic_vector(1056, 16),
3161 => conv_std_logic_vector(1068, 16),
3162 => conv_std_logic_vector(1080, 16),
3163 => conv_std_logic_vector(1092, 16),
3164 => conv_std_logic_vector(1104, 16),
3165 => conv_std_logic_vector(1116, 16),
3166 => conv_std_logic_vector(1128, 16),
3167 => conv_std_logic_vector(1140, 16),
3168 => conv_std_logic_vector(1152, 16),
3169 => conv_std_logic_vector(1164, 16),
3170 => conv_std_logic_vector(1176, 16),
3171 => conv_std_logic_vector(1188, 16),
3172 => conv_std_logic_vector(1200, 16),
3173 => conv_std_logic_vector(1212, 16),
3174 => conv_std_logic_vector(1224, 16),
3175 => conv_std_logic_vector(1236, 16),
3176 => conv_std_logic_vector(1248, 16),
3177 => conv_std_logic_vector(1260, 16),
3178 => conv_std_logic_vector(1272, 16),
3179 => conv_std_logic_vector(1284, 16),
3180 => conv_std_logic_vector(1296, 16),
3181 => conv_std_logic_vector(1308, 16),
3182 => conv_std_logic_vector(1320, 16),
3183 => conv_std_logic_vector(1332, 16),
3184 => conv_std_logic_vector(1344, 16),
3185 => conv_std_logic_vector(1356, 16),
3186 => conv_std_logic_vector(1368, 16),
3187 => conv_std_logic_vector(1380, 16),
3188 => conv_std_logic_vector(1392, 16),
3189 => conv_std_logic_vector(1404, 16),
3190 => conv_std_logic_vector(1416, 16),
3191 => conv_std_logic_vector(1428, 16),
3192 => conv_std_logic_vector(1440, 16),
3193 => conv_std_logic_vector(1452, 16),
3194 => conv_std_logic_vector(1464, 16),
3195 => conv_std_logic_vector(1476, 16),
3196 => conv_std_logic_vector(1488, 16),
3197 => conv_std_logic_vector(1500, 16),
3198 => conv_std_logic_vector(1512, 16),
3199 => conv_std_logic_vector(1524, 16),
3200 => conv_std_logic_vector(1536, 16),
3201 => conv_std_logic_vector(1548, 16),
3202 => conv_std_logic_vector(1560, 16),
3203 => conv_std_logic_vector(1572, 16),
3204 => conv_std_logic_vector(1584, 16),
3205 => conv_std_logic_vector(1596, 16),
3206 => conv_std_logic_vector(1608, 16),
3207 => conv_std_logic_vector(1620, 16),
3208 => conv_std_logic_vector(1632, 16),
3209 => conv_std_logic_vector(1644, 16),
3210 => conv_std_logic_vector(1656, 16),
3211 => conv_std_logic_vector(1668, 16),
3212 => conv_std_logic_vector(1680, 16),
3213 => conv_std_logic_vector(1692, 16),
3214 => conv_std_logic_vector(1704, 16),
3215 => conv_std_logic_vector(1716, 16),
3216 => conv_std_logic_vector(1728, 16),
3217 => conv_std_logic_vector(1740, 16),
3218 => conv_std_logic_vector(1752, 16),
3219 => conv_std_logic_vector(1764, 16),
3220 => conv_std_logic_vector(1776, 16),
3221 => conv_std_logic_vector(1788, 16),
3222 => conv_std_logic_vector(1800, 16),
3223 => conv_std_logic_vector(1812, 16),
3224 => conv_std_logic_vector(1824, 16),
3225 => conv_std_logic_vector(1836, 16),
3226 => conv_std_logic_vector(1848, 16),
3227 => conv_std_logic_vector(1860, 16),
3228 => conv_std_logic_vector(1872, 16),
3229 => conv_std_logic_vector(1884, 16),
3230 => conv_std_logic_vector(1896, 16),
3231 => conv_std_logic_vector(1908, 16),
3232 => conv_std_logic_vector(1920, 16),
3233 => conv_std_logic_vector(1932, 16),
3234 => conv_std_logic_vector(1944, 16),
3235 => conv_std_logic_vector(1956, 16),
3236 => conv_std_logic_vector(1968, 16),
3237 => conv_std_logic_vector(1980, 16),
3238 => conv_std_logic_vector(1992, 16),
3239 => conv_std_logic_vector(2004, 16),
3240 => conv_std_logic_vector(2016, 16),
3241 => conv_std_logic_vector(2028, 16),
3242 => conv_std_logic_vector(2040, 16),
3243 => conv_std_logic_vector(2052, 16),
3244 => conv_std_logic_vector(2064, 16),
3245 => conv_std_logic_vector(2076, 16),
3246 => conv_std_logic_vector(2088, 16),
3247 => conv_std_logic_vector(2100, 16),
3248 => conv_std_logic_vector(2112, 16),
3249 => conv_std_logic_vector(2124, 16),
3250 => conv_std_logic_vector(2136, 16),
3251 => conv_std_logic_vector(2148, 16),
3252 => conv_std_logic_vector(2160, 16),
3253 => conv_std_logic_vector(2172, 16),
3254 => conv_std_logic_vector(2184, 16),
3255 => conv_std_logic_vector(2196, 16),
3256 => conv_std_logic_vector(2208, 16),
3257 => conv_std_logic_vector(2220, 16),
3258 => conv_std_logic_vector(2232, 16),
3259 => conv_std_logic_vector(2244, 16),
3260 => conv_std_logic_vector(2256, 16),
3261 => conv_std_logic_vector(2268, 16),
3262 => conv_std_logic_vector(2280, 16),
3263 => conv_std_logic_vector(2292, 16),
3264 => conv_std_logic_vector(2304, 16),
3265 => conv_std_logic_vector(2316, 16),
3266 => conv_std_logic_vector(2328, 16),
3267 => conv_std_logic_vector(2340, 16),
3268 => conv_std_logic_vector(2352, 16),
3269 => conv_std_logic_vector(2364, 16),
3270 => conv_std_logic_vector(2376, 16),
3271 => conv_std_logic_vector(2388, 16),
3272 => conv_std_logic_vector(2400, 16),
3273 => conv_std_logic_vector(2412, 16),
3274 => conv_std_logic_vector(2424, 16),
3275 => conv_std_logic_vector(2436, 16),
3276 => conv_std_logic_vector(2448, 16),
3277 => conv_std_logic_vector(2460, 16),
3278 => conv_std_logic_vector(2472, 16),
3279 => conv_std_logic_vector(2484, 16),
3280 => conv_std_logic_vector(2496, 16),
3281 => conv_std_logic_vector(2508, 16),
3282 => conv_std_logic_vector(2520, 16),
3283 => conv_std_logic_vector(2532, 16),
3284 => conv_std_logic_vector(2544, 16),
3285 => conv_std_logic_vector(2556, 16),
3286 => conv_std_logic_vector(2568, 16),
3287 => conv_std_logic_vector(2580, 16),
3288 => conv_std_logic_vector(2592, 16),
3289 => conv_std_logic_vector(2604, 16),
3290 => conv_std_logic_vector(2616, 16),
3291 => conv_std_logic_vector(2628, 16),
3292 => conv_std_logic_vector(2640, 16),
3293 => conv_std_logic_vector(2652, 16),
3294 => conv_std_logic_vector(2664, 16),
3295 => conv_std_logic_vector(2676, 16),
3296 => conv_std_logic_vector(2688, 16),
3297 => conv_std_logic_vector(2700, 16),
3298 => conv_std_logic_vector(2712, 16),
3299 => conv_std_logic_vector(2724, 16),
3300 => conv_std_logic_vector(2736, 16),
3301 => conv_std_logic_vector(2748, 16),
3302 => conv_std_logic_vector(2760, 16),
3303 => conv_std_logic_vector(2772, 16),
3304 => conv_std_logic_vector(2784, 16),
3305 => conv_std_logic_vector(2796, 16),
3306 => conv_std_logic_vector(2808, 16),
3307 => conv_std_logic_vector(2820, 16),
3308 => conv_std_logic_vector(2832, 16),
3309 => conv_std_logic_vector(2844, 16),
3310 => conv_std_logic_vector(2856, 16),
3311 => conv_std_logic_vector(2868, 16),
3312 => conv_std_logic_vector(2880, 16),
3313 => conv_std_logic_vector(2892, 16),
3314 => conv_std_logic_vector(2904, 16),
3315 => conv_std_logic_vector(2916, 16),
3316 => conv_std_logic_vector(2928, 16),
3317 => conv_std_logic_vector(2940, 16),
3318 => conv_std_logic_vector(2952, 16),
3319 => conv_std_logic_vector(2964, 16),
3320 => conv_std_logic_vector(2976, 16),
3321 => conv_std_logic_vector(2988, 16),
3322 => conv_std_logic_vector(3000, 16),
3323 => conv_std_logic_vector(3012, 16),
3324 => conv_std_logic_vector(3024, 16),
3325 => conv_std_logic_vector(3036, 16),
3326 => conv_std_logic_vector(3048, 16),
3327 => conv_std_logic_vector(3060, 16),
3328 => conv_std_logic_vector(0, 16),
3329 => conv_std_logic_vector(13, 16),
3330 => conv_std_logic_vector(26, 16),
3331 => conv_std_logic_vector(39, 16),
3332 => conv_std_logic_vector(52, 16),
3333 => conv_std_logic_vector(65, 16),
3334 => conv_std_logic_vector(78, 16),
3335 => conv_std_logic_vector(91, 16),
3336 => conv_std_logic_vector(104, 16),
3337 => conv_std_logic_vector(117, 16),
3338 => conv_std_logic_vector(130, 16),
3339 => conv_std_logic_vector(143, 16),
3340 => conv_std_logic_vector(156, 16),
3341 => conv_std_logic_vector(169, 16),
3342 => conv_std_logic_vector(182, 16),
3343 => conv_std_logic_vector(195, 16),
3344 => conv_std_logic_vector(208, 16),
3345 => conv_std_logic_vector(221, 16),
3346 => conv_std_logic_vector(234, 16),
3347 => conv_std_logic_vector(247, 16),
3348 => conv_std_logic_vector(260, 16),
3349 => conv_std_logic_vector(273, 16),
3350 => conv_std_logic_vector(286, 16),
3351 => conv_std_logic_vector(299, 16),
3352 => conv_std_logic_vector(312, 16),
3353 => conv_std_logic_vector(325, 16),
3354 => conv_std_logic_vector(338, 16),
3355 => conv_std_logic_vector(351, 16),
3356 => conv_std_logic_vector(364, 16),
3357 => conv_std_logic_vector(377, 16),
3358 => conv_std_logic_vector(390, 16),
3359 => conv_std_logic_vector(403, 16),
3360 => conv_std_logic_vector(416, 16),
3361 => conv_std_logic_vector(429, 16),
3362 => conv_std_logic_vector(442, 16),
3363 => conv_std_logic_vector(455, 16),
3364 => conv_std_logic_vector(468, 16),
3365 => conv_std_logic_vector(481, 16),
3366 => conv_std_logic_vector(494, 16),
3367 => conv_std_logic_vector(507, 16),
3368 => conv_std_logic_vector(520, 16),
3369 => conv_std_logic_vector(533, 16),
3370 => conv_std_logic_vector(546, 16),
3371 => conv_std_logic_vector(559, 16),
3372 => conv_std_logic_vector(572, 16),
3373 => conv_std_logic_vector(585, 16),
3374 => conv_std_logic_vector(598, 16),
3375 => conv_std_logic_vector(611, 16),
3376 => conv_std_logic_vector(624, 16),
3377 => conv_std_logic_vector(637, 16),
3378 => conv_std_logic_vector(650, 16),
3379 => conv_std_logic_vector(663, 16),
3380 => conv_std_logic_vector(676, 16),
3381 => conv_std_logic_vector(689, 16),
3382 => conv_std_logic_vector(702, 16),
3383 => conv_std_logic_vector(715, 16),
3384 => conv_std_logic_vector(728, 16),
3385 => conv_std_logic_vector(741, 16),
3386 => conv_std_logic_vector(754, 16),
3387 => conv_std_logic_vector(767, 16),
3388 => conv_std_logic_vector(780, 16),
3389 => conv_std_logic_vector(793, 16),
3390 => conv_std_logic_vector(806, 16),
3391 => conv_std_logic_vector(819, 16),
3392 => conv_std_logic_vector(832, 16),
3393 => conv_std_logic_vector(845, 16),
3394 => conv_std_logic_vector(858, 16),
3395 => conv_std_logic_vector(871, 16),
3396 => conv_std_logic_vector(884, 16),
3397 => conv_std_logic_vector(897, 16),
3398 => conv_std_logic_vector(910, 16),
3399 => conv_std_logic_vector(923, 16),
3400 => conv_std_logic_vector(936, 16),
3401 => conv_std_logic_vector(949, 16),
3402 => conv_std_logic_vector(962, 16),
3403 => conv_std_logic_vector(975, 16),
3404 => conv_std_logic_vector(988, 16),
3405 => conv_std_logic_vector(1001, 16),
3406 => conv_std_logic_vector(1014, 16),
3407 => conv_std_logic_vector(1027, 16),
3408 => conv_std_logic_vector(1040, 16),
3409 => conv_std_logic_vector(1053, 16),
3410 => conv_std_logic_vector(1066, 16),
3411 => conv_std_logic_vector(1079, 16),
3412 => conv_std_logic_vector(1092, 16),
3413 => conv_std_logic_vector(1105, 16),
3414 => conv_std_logic_vector(1118, 16),
3415 => conv_std_logic_vector(1131, 16),
3416 => conv_std_logic_vector(1144, 16),
3417 => conv_std_logic_vector(1157, 16),
3418 => conv_std_logic_vector(1170, 16),
3419 => conv_std_logic_vector(1183, 16),
3420 => conv_std_logic_vector(1196, 16),
3421 => conv_std_logic_vector(1209, 16),
3422 => conv_std_logic_vector(1222, 16),
3423 => conv_std_logic_vector(1235, 16),
3424 => conv_std_logic_vector(1248, 16),
3425 => conv_std_logic_vector(1261, 16),
3426 => conv_std_logic_vector(1274, 16),
3427 => conv_std_logic_vector(1287, 16),
3428 => conv_std_logic_vector(1300, 16),
3429 => conv_std_logic_vector(1313, 16),
3430 => conv_std_logic_vector(1326, 16),
3431 => conv_std_logic_vector(1339, 16),
3432 => conv_std_logic_vector(1352, 16),
3433 => conv_std_logic_vector(1365, 16),
3434 => conv_std_logic_vector(1378, 16),
3435 => conv_std_logic_vector(1391, 16),
3436 => conv_std_logic_vector(1404, 16),
3437 => conv_std_logic_vector(1417, 16),
3438 => conv_std_logic_vector(1430, 16),
3439 => conv_std_logic_vector(1443, 16),
3440 => conv_std_logic_vector(1456, 16),
3441 => conv_std_logic_vector(1469, 16),
3442 => conv_std_logic_vector(1482, 16),
3443 => conv_std_logic_vector(1495, 16),
3444 => conv_std_logic_vector(1508, 16),
3445 => conv_std_logic_vector(1521, 16),
3446 => conv_std_logic_vector(1534, 16),
3447 => conv_std_logic_vector(1547, 16),
3448 => conv_std_logic_vector(1560, 16),
3449 => conv_std_logic_vector(1573, 16),
3450 => conv_std_logic_vector(1586, 16),
3451 => conv_std_logic_vector(1599, 16),
3452 => conv_std_logic_vector(1612, 16),
3453 => conv_std_logic_vector(1625, 16),
3454 => conv_std_logic_vector(1638, 16),
3455 => conv_std_logic_vector(1651, 16),
3456 => conv_std_logic_vector(1664, 16),
3457 => conv_std_logic_vector(1677, 16),
3458 => conv_std_logic_vector(1690, 16),
3459 => conv_std_logic_vector(1703, 16),
3460 => conv_std_logic_vector(1716, 16),
3461 => conv_std_logic_vector(1729, 16),
3462 => conv_std_logic_vector(1742, 16),
3463 => conv_std_logic_vector(1755, 16),
3464 => conv_std_logic_vector(1768, 16),
3465 => conv_std_logic_vector(1781, 16),
3466 => conv_std_logic_vector(1794, 16),
3467 => conv_std_logic_vector(1807, 16),
3468 => conv_std_logic_vector(1820, 16),
3469 => conv_std_logic_vector(1833, 16),
3470 => conv_std_logic_vector(1846, 16),
3471 => conv_std_logic_vector(1859, 16),
3472 => conv_std_logic_vector(1872, 16),
3473 => conv_std_logic_vector(1885, 16),
3474 => conv_std_logic_vector(1898, 16),
3475 => conv_std_logic_vector(1911, 16),
3476 => conv_std_logic_vector(1924, 16),
3477 => conv_std_logic_vector(1937, 16),
3478 => conv_std_logic_vector(1950, 16),
3479 => conv_std_logic_vector(1963, 16),
3480 => conv_std_logic_vector(1976, 16),
3481 => conv_std_logic_vector(1989, 16),
3482 => conv_std_logic_vector(2002, 16),
3483 => conv_std_logic_vector(2015, 16),
3484 => conv_std_logic_vector(2028, 16),
3485 => conv_std_logic_vector(2041, 16),
3486 => conv_std_logic_vector(2054, 16),
3487 => conv_std_logic_vector(2067, 16),
3488 => conv_std_logic_vector(2080, 16),
3489 => conv_std_logic_vector(2093, 16),
3490 => conv_std_logic_vector(2106, 16),
3491 => conv_std_logic_vector(2119, 16),
3492 => conv_std_logic_vector(2132, 16),
3493 => conv_std_logic_vector(2145, 16),
3494 => conv_std_logic_vector(2158, 16),
3495 => conv_std_logic_vector(2171, 16),
3496 => conv_std_logic_vector(2184, 16),
3497 => conv_std_logic_vector(2197, 16),
3498 => conv_std_logic_vector(2210, 16),
3499 => conv_std_logic_vector(2223, 16),
3500 => conv_std_logic_vector(2236, 16),
3501 => conv_std_logic_vector(2249, 16),
3502 => conv_std_logic_vector(2262, 16),
3503 => conv_std_logic_vector(2275, 16),
3504 => conv_std_logic_vector(2288, 16),
3505 => conv_std_logic_vector(2301, 16),
3506 => conv_std_logic_vector(2314, 16),
3507 => conv_std_logic_vector(2327, 16),
3508 => conv_std_logic_vector(2340, 16),
3509 => conv_std_logic_vector(2353, 16),
3510 => conv_std_logic_vector(2366, 16),
3511 => conv_std_logic_vector(2379, 16),
3512 => conv_std_logic_vector(2392, 16),
3513 => conv_std_logic_vector(2405, 16),
3514 => conv_std_logic_vector(2418, 16),
3515 => conv_std_logic_vector(2431, 16),
3516 => conv_std_logic_vector(2444, 16),
3517 => conv_std_logic_vector(2457, 16),
3518 => conv_std_logic_vector(2470, 16),
3519 => conv_std_logic_vector(2483, 16),
3520 => conv_std_logic_vector(2496, 16),
3521 => conv_std_logic_vector(2509, 16),
3522 => conv_std_logic_vector(2522, 16),
3523 => conv_std_logic_vector(2535, 16),
3524 => conv_std_logic_vector(2548, 16),
3525 => conv_std_logic_vector(2561, 16),
3526 => conv_std_logic_vector(2574, 16),
3527 => conv_std_logic_vector(2587, 16),
3528 => conv_std_logic_vector(2600, 16),
3529 => conv_std_logic_vector(2613, 16),
3530 => conv_std_logic_vector(2626, 16),
3531 => conv_std_logic_vector(2639, 16),
3532 => conv_std_logic_vector(2652, 16),
3533 => conv_std_logic_vector(2665, 16),
3534 => conv_std_logic_vector(2678, 16),
3535 => conv_std_logic_vector(2691, 16),
3536 => conv_std_logic_vector(2704, 16),
3537 => conv_std_logic_vector(2717, 16),
3538 => conv_std_logic_vector(2730, 16),
3539 => conv_std_logic_vector(2743, 16),
3540 => conv_std_logic_vector(2756, 16),
3541 => conv_std_logic_vector(2769, 16),
3542 => conv_std_logic_vector(2782, 16),
3543 => conv_std_logic_vector(2795, 16),
3544 => conv_std_logic_vector(2808, 16),
3545 => conv_std_logic_vector(2821, 16),
3546 => conv_std_logic_vector(2834, 16),
3547 => conv_std_logic_vector(2847, 16),
3548 => conv_std_logic_vector(2860, 16),
3549 => conv_std_logic_vector(2873, 16),
3550 => conv_std_logic_vector(2886, 16),
3551 => conv_std_logic_vector(2899, 16),
3552 => conv_std_logic_vector(2912, 16),
3553 => conv_std_logic_vector(2925, 16),
3554 => conv_std_logic_vector(2938, 16),
3555 => conv_std_logic_vector(2951, 16),
3556 => conv_std_logic_vector(2964, 16),
3557 => conv_std_logic_vector(2977, 16),
3558 => conv_std_logic_vector(2990, 16),
3559 => conv_std_logic_vector(3003, 16),
3560 => conv_std_logic_vector(3016, 16),
3561 => conv_std_logic_vector(3029, 16),
3562 => conv_std_logic_vector(3042, 16),
3563 => conv_std_logic_vector(3055, 16),
3564 => conv_std_logic_vector(3068, 16),
3565 => conv_std_logic_vector(3081, 16),
3566 => conv_std_logic_vector(3094, 16),
3567 => conv_std_logic_vector(3107, 16),
3568 => conv_std_logic_vector(3120, 16),
3569 => conv_std_logic_vector(3133, 16),
3570 => conv_std_logic_vector(3146, 16),
3571 => conv_std_logic_vector(3159, 16),
3572 => conv_std_logic_vector(3172, 16),
3573 => conv_std_logic_vector(3185, 16),
3574 => conv_std_logic_vector(3198, 16),
3575 => conv_std_logic_vector(3211, 16),
3576 => conv_std_logic_vector(3224, 16),
3577 => conv_std_logic_vector(3237, 16),
3578 => conv_std_logic_vector(3250, 16),
3579 => conv_std_logic_vector(3263, 16),
3580 => conv_std_logic_vector(3276, 16),
3581 => conv_std_logic_vector(3289, 16),
3582 => conv_std_logic_vector(3302, 16),
3583 => conv_std_logic_vector(3315, 16),
3584 => conv_std_logic_vector(0, 16),
3585 => conv_std_logic_vector(14, 16),
3586 => conv_std_logic_vector(28, 16),
3587 => conv_std_logic_vector(42, 16),
3588 => conv_std_logic_vector(56, 16),
3589 => conv_std_logic_vector(70, 16),
3590 => conv_std_logic_vector(84, 16),
3591 => conv_std_logic_vector(98, 16),
3592 => conv_std_logic_vector(112, 16),
3593 => conv_std_logic_vector(126, 16),
3594 => conv_std_logic_vector(140, 16),
3595 => conv_std_logic_vector(154, 16),
3596 => conv_std_logic_vector(168, 16),
3597 => conv_std_logic_vector(182, 16),
3598 => conv_std_logic_vector(196, 16),
3599 => conv_std_logic_vector(210, 16),
3600 => conv_std_logic_vector(224, 16),
3601 => conv_std_logic_vector(238, 16),
3602 => conv_std_logic_vector(252, 16),
3603 => conv_std_logic_vector(266, 16),
3604 => conv_std_logic_vector(280, 16),
3605 => conv_std_logic_vector(294, 16),
3606 => conv_std_logic_vector(308, 16),
3607 => conv_std_logic_vector(322, 16),
3608 => conv_std_logic_vector(336, 16),
3609 => conv_std_logic_vector(350, 16),
3610 => conv_std_logic_vector(364, 16),
3611 => conv_std_logic_vector(378, 16),
3612 => conv_std_logic_vector(392, 16),
3613 => conv_std_logic_vector(406, 16),
3614 => conv_std_logic_vector(420, 16),
3615 => conv_std_logic_vector(434, 16),
3616 => conv_std_logic_vector(448, 16),
3617 => conv_std_logic_vector(462, 16),
3618 => conv_std_logic_vector(476, 16),
3619 => conv_std_logic_vector(490, 16),
3620 => conv_std_logic_vector(504, 16),
3621 => conv_std_logic_vector(518, 16),
3622 => conv_std_logic_vector(532, 16),
3623 => conv_std_logic_vector(546, 16),
3624 => conv_std_logic_vector(560, 16),
3625 => conv_std_logic_vector(574, 16),
3626 => conv_std_logic_vector(588, 16),
3627 => conv_std_logic_vector(602, 16),
3628 => conv_std_logic_vector(616, 16),
3629 => conv_std_logic_vector(630, 16),
3630 => conv_std_logic_vector(644, 16),
3631 => conv_std_logic_vector(658, 16),
3632 => conv_std_logic_vector(672, 16),
3633 => conv_std_logic_vector(686, 16),
3634 => conv_std_logic_vector(700, 16),
3635 => conv_std_logic_vector(714, 16),
3636 => conv_std_logic_vector(728, 16),
3637 => conv_std_logic_vector(742, 16),
3638 => conv_std_logic_vector(756, 16),
3639 => conv_std_logic_vector(770, 16),
3640 => conv_std_logic_vector(784, 16),
3641 => conv_std_logic_vector(798, 16),
3642 => conv_std_logic_vector(812, 16),
3643 => conv_std_logic_vector(826, 16),
3644 => conv_std_logic_vector(840, 16),
3645 => conv_std_logic_vector(854, 16),
3646 => conv_std_logic_vector(868, 16),
3647 => conv_std_logic_vector(882, 16),
3648 => conv_std_logic_vector(896, 16),
3649 => conv_std_logic_vector(910, 16),
3650 => conv_std_logic_vector(924, 16),
3651 => conv_std_logic_vector(938, 16),
3652 => conv_std_logic_vector(952, 16),
3653 => conv_std_logic_vector(966, 16),
3654 => conv_std_logic_vector(980, 16),
3655 => conv_std_logic_vector(994, 16),
3656 => conv_std_logic_vector(1008, 16),
3657 => conv_std_logic_vector(1022, 16),
3658 => conv_std_logic_vector(1036, 16),
3659 => conv_std_logic_vector(1050, 16),
3660 => conv_std_logic_vector(1064, 16),
3661 => conv_std_logic_vector(1078, 16),
3662 => conv_std_logic_vector(1092, 16),
3663 => conv_std_logic_vector(1106, 16),
3664 => conv_std_logic_vector(1120, 16),
3665 => conv_std_logic_vector(1134, 16),
3666 => conv_std_logic_vector(1148, 16),
3667 => conv_std_logic_vector(1162, 16),
3668 => conv_std_logic_vector(1176, 16),
3669 => conv_std_logic_vector(1190, 16),
3670 => conv_std_logic_vector(1204, 16),
3671 => conv_std_logic_vector(1218, 16),
3672 => conv_std_logic_vector(1232, 16),
3673 => conv_std_logic_vector(1246, 16),
3674 => conv_std_logic_vector(1260, 16),
3675 => conv_std_logic_vector(1274, 16),
3676 => conv_std_logic_vector(1288, 16),
3677 => conv_std_logic_vector(1302, 16),
3678 => conv_std_logic_vector(1316, 16),
3679 => conv_std_logic_vector(1330, 16),
3680 => conv_std_logic_vector(1344, 16),
3681 => conv_std_logic_vector(1358, 16),
3682 => conv_std_logic_vector(1372, 16),
3683 => conv_std_logic_vector(1386, 16),
3684 => conv_std_logic_vector(1400, 16),
3685 => conv_std_logic_vector(1414, 16),
3686 => conv_std_logic_vector(1428, 16),
3687 => conv_std_logic_vector(1442, 16),
3688 => conv_std_logic_vector(1456, 16),
3689 => conv_std_logic_vector(1470, 16),
3690 => conv_std_logic_vector(1484, 16),
3691 => conv_std_logic_vector(1498, 16),
3692 => conv_std_logic_vector(1512, 16),
3693 => conv_std_logic_vector(1526, 16),
3694 => conv_std_logic_vector(1540, 16),
3695 => conv_std_logic_vector(1554, 16),
3696 => conv_std_logic_vector(1568, 16),
3697 => conv_std_logic_vector(1582, 16),
3698 => conv_std_logic_vector(1596, 16),
3699 => conv_std_logic_vector(1610, 16),
3700 => conv_std_logic_vector(1624, 16),
3701 => conv_std_logic_vector(1638, 16),
3702 => conv_std_logic_vector(1652, 16),
3703 => conv_std_logic_vector(1666, 16),
3704 => conv_std_logic_vector(1680, 16),
3705 => conv_std_logic_vector(1694, 16),
3706 => conv_std_logic_vector(1708, 16),
3707 => conv_std_logic_vector(1722, 16),
3708 => conv_std_logic_vector(1736, 16),
3709 => conv_std_logic_vector(1750, 16),
3710 => conv_std_logic_vector(1764, 16),
3711 => conv_std_logic_vector(1778, 16),
3712 => conv_std_logic_vector(1792, 16),
3713 => conv_std_logic_vector(1806, 16),
3714 => conv_std_logic_vector(1820, 16),
3715 => conv_std_logic_vector(1834, 16),
3716 => conv_std_logic_vector(1848, 16),
3717 => conv_std_logic_vector(1862, 16),
3718 => conv_std_logic_vector(1876, 16),
3719 => conv_std_logic_vector(1890, 16),
3720 => conv_std_logic_vector(1904, 16),
3721 => conv_std_logic_vector(1918, 16),
3722 => conv_std_logic_vector(1932, 16),
3723 => conv_std_logic_vector(1946, 16),
3724 => conv_std_logic_vector(1960, 16),
3725 => conv_std_logic_vector(1974, 16),
3726 => conv_std_logic_vector(1988, 16),
3727 => conv_std_logic_vector(2002, 16),
3728 => conv_std_logic_vector(2016, 16),
3729 => conv_std_logic_vector(2030, 16),
3730 => conv_std_logic_vector(2044, 16),
3731 => conv_std_logic_vector(2058, 16),
3732 => conv_std_logic_vector(2072, 16),
3733 => conv_std_logic_vector(2086, 16),
3734 => conv_std_logic_vector(2100, 16),
3735 => conv_std_logic_vector(2114, 16),
3736 => conv_std_logic_vector(2128, 16),
3737 => conv_std_logic_vector(2142, 16),
3738 => conv_std_logic_vector(2156, 16),
3739 => conv_std_logic_vector(2170, 16),
3740 => conv_std_logic_vector(2184, 16),
3741 => conv_std_logic_vector(2198, 16),
3742 => conv_std_logic_vector(2212, 16),
3743 => conv_std_logic_vector(2226, 16),
3744 => conv_std_logic_vector(2240, 16),
3745 => conv_std_logic_vector(2254, 16),
3746 => conv_std_logic_vector(2268, 16),
3747 => conv_std_logic_vector(2282, 16),
3748 => conv_std_logic_vector(2296, 16),
3749 => conv_std_logic_vector(2310, 16),
3750 => conv_std_logic_vector(2324, 16),
3751 => conv_std_logic_vector(2338, 16),
3752 => conv_std_logic_vector(2352, 16),
3753 => conv_std_logic_vector(2366, 16),
3754 => conv_std_logic_vector(2380, 16),
3755 => conv_std_logic_vector(2394, 16),
3756 => conv_std_logic_vector(2408, 16),
3757 => conv_std_logic_vector(2422, 16),
3758 => conv_std_logic_vector(2436, 16),
3759 => conv_std_logic_vector(2450, 16),
3760 => conv_std_logic_vector(2464, 16),
3761 => conv_std_logic_vector(2478, 16),
3762 => conv_std_logic_vector(2492, 16),
3763 => conv_std_logic_vector(2506, 16),
3764 => conv_std_logic_vector(2520, 16),
3765 => conv_std_logic_vector(2534, 16),
3766 => conv_std_logic_vector(2548, 16),
3767 => conv_std_logic_vector(2562, 16),
3768 => conv_std_logic_vector(2576, 16),
3769 => conv_std_logic_vector(2590, 16),
3770 => conv_std_logic_vector(2604, 16),
3771 => conv_std_logic_vector(2618, 16),
3772 => conv_std_logic_vector(2632, 16),
3773 => conv_std_logic_vector(2646, 16),
3774 => conv_std_logic_vector(2660, 16),
3775 => conv_std_logic_vector(2674, 16),
3776 => conv_std_logic_vector(2688, 16),
3777 => conv_std_logic_vector(2702, 16),
3778 => conv_std_logic_vector(2716, 16),
3779 => conv_std_logic_vector(2730, 16),
3780 => conv_std_logic_vector(2744, 16),
3781 => conv_std_logic_vector(2758, 16),
3782 => conv_std_logic_vector(2772, 16),
3783 => conv_std_logic_vector(2786, 16),
3784 => conv_std_logic_vector(2800, 16),
3785 => conv_std_logic_vector(2814, 16),
3786 => conv_std_logic_vector(2828, 16),
3787 => conv_std_logic_vector(2842, 16),
3788 => conv_std_logic_vector(2856, 16),
3789 => conv_std_logic_vector(2870, 16),
3790 => conv_std_logic_vector(2884, 16),
3791 => conv_std_logic_vector(2898, 16),
3792 => conv_std_logic_vector(2912, 16),
3793 => conv_std_logic_vector(2926, 16),
3794 => conv_std_logic_vector(2940, 16),
3795 => conv_std_logic_vector(2954, 16),
3796 => conv_std_logic_vector(2968, 16),
3797 => conv_std_logic_vector(2982, 16),
3798 => conv_std_logic_vector(2996, 16),
3799 => conv_std_logic_vector(3010, 16),
3800 => conv_std_logic_vector(3024, 16),
3801 => conv_std_logic_vector(3038, 16),
3802 => conv_std_logic_vector(3052, 16),
3803 => conv_std_logic_vector(3066, 16),
3804 => conv_std_logic_vector(3080, 16),
3805 => conv_std_logic_vector(3094, 16),
3806 => conv_std_logic_vector(3108, 16),
3807 => conv_std_logic_vector(3122, 16),
3808 => conv_std_logic_vector(3136, 16),
3809 => conv_std_logic_vector(3150, 16),
3810 => conv_std_logic_vector(3164, 16),
3811 => conv_std_logic_vector(3178, 16),
3812 => conv_std_logic_vector(3192, 16),
3813 => conv_std_logic_vector(3206, 16),
3814 => conv_std_logic_vector(3220, 16),
3815 => conv_std_logic_vector(3234, 16),
3816 => conv_std_logic_vector(3248, 16),
3817 => conv_std_logic_vector(3262, 16),
3818 => conv_std_logic_vector(3276, 16),
3819 => conv_std_logic_vector(3290, 16),
3820 => conv_std_logic_vector(3304, 16),
3821 => conv_std_logic_vector(3318, 16),
3822 => conv_std_logic_vector(3332, 16),
3823 => conv_std_logic_vector(3346, 16),
3824 => conv_std_logic_vector(3360, 16),
3825 => conv_std_logic_vector(3374, 16),
3826 => conv_std_logic_vector(3388, 16),
3827 => conv_std_logic_vector(3402, 16),
3828 => conv_std_logic_vector(3416, 16),
3829 => conv_std_logic_vector(3430, 16),
3830 => conv_std_logic_vector(3444, 16),
3831 => conv_std_logic_vector(3458, 16),
3832 => conv_std_logic_vector(3472, 16),
3833 => conv_std_logic_vector(3486, 16),
3834 => conv_std_logic_vector(3500, 16),
3835 => conv_std_logic_vector(3514, 16),
3836 => conv_std_logic_vector(3528, 16),
3837 => conv_std_logic_vector(3542, 16),
3838 => conv_std_logic_vector(3556, 16),
3839 => conv_std_logic_vector(3570, 16),
3840 => conv_std_logic_vector(0, 16),
3841 => conv_std_logic_vector(15, 16),
3842 => conv_std_logic_vector(30, 16),
3843 => conv_std_logic_vector(45, 16),
3844 => conv_std_logic_vector(60, 16),
3845 => conv_std_logic_vector(75, 16),
3846 => conv_std_logic_vector(90, 16),
3847 => conv_std_logic_vector(105, 16),
3848 => conv_std_logic_vector(120, 16),
3849 => conv_std_logic_vector(135, 16),
3850 => conv_std_logic_vector(150, 16),
3851 => conv_std_logic_vector(165, 16),
3852 => conv_std_logic_vector(180, 16),
3853 => conv_std_logic_vector(195, 16),
3854 => conv_std_logic_vector(210, 16),
3855 => conv_std_logic_vector(225, 16),
3856 => conv_std_logic_vector(240, 16),
3857 => conv_std_logic_vector(255, 16),
3858 => conv_std_logic_vector(270, 16),
3859 => conv_std_logic_vector(285, 16),
3860 => conv_std_logic_vector(300, 16),
3861 => conv_std_logic_vector(315, 16),
3862 => conv_std_logic_vector(330, 16),
3863 => conv_std_logic_vector(345, 16),
3864 => conv_std_logic_vector(360, 16),
3865 => conv_std_logic_vector(375, 16),
3866 => conv_std_logic_vector(390, 16),
3867 => conv_std_logic_vector(405, 16),
3868 => conv_std_logic_vector(420, 16),
3869 => conv_std_logic_vector(435, 16),
3870 => conv_std_logic_vector(450, 16),
3871 => conv_std_logic_vector(465, 16),
3872 => conv_std_logic_vector(480, 16),
3873 => conv_std_logic_vector(495, 16),
3874 => conv_std_logic_vector(510, 16),
3875 => conv_std_logic_vector(525, 16),
3876 => conv_std_logic_vector(540, 16),
3877 => conv_std_logic_vector(555, 16),
3878 => conv_std_logic_vector(570, 16),
3879 => conv_std_logic_vector(585, 16),
3880 => conv_std_logic_vector(600, 16),
3881 => conv_std_logic_vector(615, 16),
3882 => conv_std_logic_vector(630, 16),
3883 => conv_std_logic_vector(645, 16),
3884 => conv_std_logic_vector(660, 16),
3885 => conv_std_logic_vector(675, 16),
3886 => conv_std_logic_vector(690, 16),
3887 => conv_std_logic_vector(705, 16),
3888 => conv_std_logic_vector(720, 16),
3889 => conv_std_logic_vector(735, 16),
3890 => conv_std_logic_vector(750, 16),
3891 => conv_std_logic_vector(765, 16),
3892 => conv_std_logic_vector(780, 16),
3893 => conv_std_logic_vector(795, 16),
3894 => conv_std_logic_vector(810, 16),
3895 => conv_std_logic_vector(825, 16),
3896 => conv_std_logic_vector(840, 16),
3897 => conv_std_logic_vector(855, 16),
3898 => conv_std_logic_vector(870, 16),
3899 => conv_std_logic_vector(885, 16),
3900 => conv_std_logic_vector(900, 16),
3901 => conv_std_logic_vector(915, 16),
3902 => conv_std_logic_vector(930, 16),
3903 => conv_std_logic_vector(945, 16),
3904 => conv_std_logic_vector(960, 16),
3905 => conv_std_logic_vector(975, 16),
3906 => conv_std_logic_vector(990, 16),
3907 => conv_std_logic_vector(1005, 16),
3908 => conv_std_logic_vector(1020, 16),
3909 => conv_std_logic_vector(1035, 16),
3910 => conv_std_logic_vector(1050, 16),
3911 => conv_std_logic_vector(1065, 16),
3912 => conv_std_logic_vector(1080, 16),
3913 => conv_std_logic_vector(1095, 16),
3914 => conv_std_logic_vector(1110, 16),
3915 => conv_std_logic_vector(1125, 16),
3916 => conv_std_logic_vector(1140, 16),
3917 => conv_std_logic_vector(1155, 16),
3918 => conv_std_logic_vector(1170, 16),
3919 => conv_std_logic_vector(1185, 16),
3920 => conv_std_logic_vector(1200, 16),
3921 => conv_std_logic_vector(1215, 16),
3922 => conv_std_logic_vector(1230, 16),
3923 => conv_std_logic_vector(1245, 16),
3924 => conv_std_logic_vector(1260, 16),
3925 => conv_std_logic_vector(1275, 16),
3926 => conv_std_logic_vector(1290, 16),
3927 => conv_std_logic_vector(1305, 16),
3928 => conv_std_logic_vector(1320, 16),
3929 => conv_std_logic_vector(1335, 16),
3930 => conv_std_logic_vector(1350, 16),
3931 => conv_std_logic_vector(1365, 16),
3932 => conv_std_logic_vector(1380, 16),
3933 => conv_std_logic_vector(1395, 16),
3934 => conv_std_logic_vector(1410, 16),
3935 => conv_std_logic_vector(1425, 16),
3936 => conv_std_logic_vector(1440, 16),
3937 => conv_std_logic_vector(1455, 16),
3938 => conv_std_logic_vector(1470, 16),
3939 => conv_std_logic_vector(1485, 16),
3940 => conv_std_logic_vector(1500, 16),
3941 => conv_std_logic_vector(1515, 16),
3942 => conv_std_logic_vector(1530, 16),
3943 => conv_std_logic_vector(1545, 16),
3944 => conv_std_logic_vector(1560, 16),
3945 => conv_std_logic_vector(1575, 16),
3946 => conv_std_logic_vector(1590, 16),
3947 => conv_std_logic_vector(1605, 16),
3948 => conv_std_logic_vector(1620, 16),
3949 => conv_std_logic_vector(1635, 16),
3950 => conv_std_logic_vector(1650, 16),
3951 => conv_std_logic_vector(1665, 16),
3952 => conv_std_logic_vector(1680, 16),
3953 => conv_std_logic_vector(1695, 16),
3954 => conv_std_logic_vector(1710, 16),
3955 => conv_std_logic_vector(1725, 16),
3956 => conv_std_logic_vector(1740, 16),
3957 => conv_std_logic_vector(1755, 16),
3958 => conv_std_logic_vector(1770, 16),
3959 => conv_std_logic_vector(1785, 16),
3960 => conv_std_logic_vector(1800, 16),
3961 => conv_std_logic_vector(1815, 16),
3962 => conv_std_logic_vector(1830, 16),
3963 => conv_std_logic_vector(1845, 16),
3964 => conv_std_logic_vector(1860, 16),
3965 => conv_std_logic_vector(1875, 16),
3966 => conv_std_logic_vector(1890, 16),
3967 => conv_std_logic_vector(1905, 16),
3968 => conv_std_logic_vector(1920, 16),
3969 => conv_std_logic_vector(1935, 16),
3970 => conv_std_logic_vector(1950, 16),
3971 => conv_std_logic_vector(1965, 16),
3972 => conv_std_logic_vector(1980, 16),
3973 => conv_std_logic_vector(1995, 16),
3974 => conv_std_logic_vector(2010, 16),
3975 => conv_std_logic_vector(2025, 16),
3976 => conv_std_logic_vector(2040, 16),
3977 => conv_std_logic_vector(2055, 16),
3978 => conv_std_logic_vector(2070, 16),
3979 => conv_std_logic_vector(2085, 16),
3980 => conv_std_logic_vector(2100, 16),
3981 => conv_std_logic_vector(2115, 16),
3982 => conv_std_logic_vector(2130, 16),
3983 => conv_std_logic_vector(2145, 16),
3984 => conv_std_logic_vector(2160, 16),
3985 => conv_std_logic_vector(2175, 16),
3986 => conv_std_logic_vector(2190, 16),
3987 => conv_std_logic_vector(2205, 16),
3988 => conv_std_logic_vector(2220, 16),
3989 => conv_std_logic_vector(2235, 16),
3990 => conv_std_logic_vector(2250, 16),
3991 => conv_std_logic_vector(2265, 16),
3992 => conv_std_logic_vector(2280, 16),
3993 => conv_std_logic_vector(2295, 16),
3994 => conv_std_logic_vector(2310, 16),
3995 => conv_std_logic_vector(2325, 16),
3996 => conv_std_logic_vector(2340, 16),
3997 => conv_std_logic_vector(2355, 16),
3998 => conv_std_logic_vector(2370, 16),
3999 => conv_std_logic_vector(2385, 16),
4000 => conv_std_logic_vector(2400, 16),
4001 => conv_std_logic_vector(2415, 16),
4002 => conv_std_logic_vector(2430, 16),
4003 => conv_std_logic_vector(2445, 16),
4004 => conv_std_logic_vector(2460, 16),
4005 => conv_std_logic_vector(2475, 16),
4006 => conv_std_logic_vector(2490, 16),
4007 => conv_std_logic_vector(2505, 16),
4008 => conv_std_logic_vector(2520, 16),
4009 => conv_std_logic_vector(2535, 16),
4010 => conv_std_logic_vector(2550, 16),
4011 => conv_std_logic_vector(2565, 16),
4012 => conv_std_logic_vector(2580, 16),
4013 => conv_std_logic_vector(2595, 16),
4014 => conv_std_logic_vector(2610, 16),
4015 => conv_std_logic_vector(2625, 16),
4016 => conv_std_logic_vector(2640, 16),
4017 => conv_std_logic_vector(2655, 16),
4018 => conv_std_logic_vector(2670, 16),
4019 => conv_std_logic_vector(2685, 16),
4020 => conv_std_logic_vector(2700, 16),
4021 => conv_std_logic_vector(2715, 16),
4022 => conv_std_logic_vector(2730, 16),
4023 => conv_std_logic_vector(2745, 16),
4024 => conv_std_logic_vector(2760, 16),
4025 => conv_std_logic_vector(2775, 16),
4026 => conv_std_logic_vector(2790, 16),
4027 => conv_std_logic_vector(2805, 16),
4028 => conv_std_logic_vector(2820, 16),
4029 => conv_std_logic_vector(2835, 16),
4030 => conv_std_logic_vector(2850, 16),
4031 => conv_std_logic_vector(2865, 16),
4032 => conv_std_logic_vector(2880, 16),
4033 => conv_std_logic_vector(2895, 16),
4034 => conv_std_logic_vector(2910, 16),
4035 => conv_std_logic_vector(2925, 16),
4036 => conv_std_logic_vector(2940, 16),
4037 => conv_std_logic_vector(2955, 16),
4038 => conv_std_logic_vector(2970, 16),
4039 => conv_std_logic_vector(2985, 16),
4040 => conv_std_logic_vector(3000, 16),
4041 => conv_std_logic_vector(3015, 16),
4042 => conv_std_logic_vector(3030, 16),
4043 => conv_std_logic_vector(3045, 16),
4044 => conv_std_logic_vector(3060, 16),
4045 => conv_std_logic_vector(3075, 16),
4046 => conv_std_logic_vector(3090, 16),
4047 => conv_std_logic_vector(3105, 16),
4048 => conv_std_logic_vector(3120, 16),
4049 => conv_std_logic_vector(3135, 16),
4050 => conv_std_logic_vector(3150, 16),
4051 => conv_std_logic_vector(3165, 16),
4052 => conv_std_logic_vector(3180, 16),
4053 => conv_std_logic_vector(3195, 16),
4054 => conv_std_logic_vector(3210, 16),
4055 => conv_std_logic_vector(3225, 16),
4056 => conv_std_logic_vector(3240, 16),
4057 => conv_std_logic_vector(3255, 16),
4058 => conv_std_logic_vector(3270, 16),
4059 => conv_std_logic_vector(3285, 16),
4060 => conv_std_logic_vector(3300, 16),
4061 => conv_std_logic_vector(3315, 16),
4062 => conv_std_logic_vector(3330, 16),
4063 => conv_std_logic_vector(3345, 16),
4064 => conv_std_logic_vector(3360, 16),
4065 => conv_std_logic_vector(3375, 16),
4066 => conv_std_logic_vector(3390, 16),
4067 => conv_std_logic_vector(3405, 16),
4068 => conv_std_logic_vector(3420, 16),
4069 => conv_std_logic_vector(3435, 16),
4070 => conv_std_logic_vector(3450, 16),
4071 => conv_std_logic_vector(3465, 16),
4072 => conv_std_logic_vector(3480, 16),
4073 => conv_std_logic_vector(3495, 16),
4074 => conv_std_logic_vector(3510, 16),
4075 => conv_std_logic_vector(3525, 16),
4076 => conv_std_logic_vector(3540, 16),
4077 => conv_std_logic_vector(3555, 16),
4078 => conv_std_logic_vector(3570, 16),
4079 => conv_std_logic_vector(3585, 16),
4080 => conv_std_logic_vector(3600, 16),
4081 => conv_std_logic_vector(3615, 16),
4082 => conv_std_logic_vector(3630, 16),
4083 => conv_std_logic_vector(3645, 16),
4084 => conv_std_logic_vector(3660, 16),
4085 => conv_std_logic_vector(3675, 16),
4086 => conv_std_logic_vector(3690, 16),
4087 => conv_std_logic_vector(3705, 16),
4088 => conv_std_logic_vector(3720, 16),
4089 => conv_std_logic_vector(3735, 16),
4090 => conv_std_logic_vector(3750, 16),
4091 => conv_std_logic_vector(3765, 16),
4092 => conv_std_logic_vector(3780, 16),
4093 => conv_std_logic_vector(3795, 16),
4094 => conv_std_logic_vector(3810, 16),
4095 => conv_std_logic_vector(3825, 16),
4096 => conv_std_logic_vector(0, 16),
4097 => conv_std_logic_vector(16, 16),
4098 => conv_std_logic_vector(32, 16),
4099 => conv_std_logic_vector(48, 16),
4100 => conv_std_logic_vector(64, 16),
4101 => conv_std_logic_vector(80, 16),
4102 => conv_std_logic_vector(96, 16),
4103 => conv_std_logic_vector(112, 16),
4104 => conv_std_logic_vector(128, 16),
4105 => conv_std_logic_vector(144, 16),
4106 => conv_std_logic_vector(160, 16),
4107 => conv_std_logic_vector(176, 16),
4108 => conv_std_logic_vector(192, 16),
4109 => conv_std_logic_vector(208, 16),
4110 => conv_std_logic_vector(224, 16),
4111 => conv_std_logic_vector(240, 16),
4112 => conv_std_logic_vector(256, 16),
4113 => conv_std_logic_vector(272, 16),
4114 => conv_std_logic_vector(288, 16),
4115 => conv_std_logic_vector(304, 16),
4116 => conv_std_logic_vector(320, 16),
4117 => conv_std_logic_vector(336, 16),
4118 => conv_std_logic_vector(352, 16),
4119 => conv_std_logic_vector(368, 16),
4120 => conv_std_logic_vector(384, 16),
4121 => conv_std_logic_vector(400, 16),
4122 => conv_std_logic_vector(416, 16),
4123 => conv_std_logic_vector(432, 16),
4124 => conv_std_logic_vector(448, 16),
4125 => conv_std_logic_vector(464, 16),
4126 => conv_std_logic_vector(480, 16),
4127 => conv_std_logic_vector(496, 16),
4128 => conv_std_logic_vector(512, 16),
4129 => conv_std_logic_vector(528, 16),
4130 => conv_std_logic_vector(544, 16),
4131 => conv_std_logic_vector(560, 16),
4132 => conv_std_logic_vector(576, 16),
4133 => conv_std_logic_vector(592, 16),
4134 => conv_std_logic_vector(608, 16),
4135 => conv_std_logic_vector(624, 16),
4136 => conv_std_logic_vector(640, 16),
4137 => conv_std_logic_vector(656, 16),
4138 => conv_std_logic_vector(672, 16),
4139 => conv_std_logic_vector(688, 16),
4140 => conv_std_logic_vector(704, 16),
4141 => conv_std_logic_vector(720, 16),
4142 => conv_std_logic_vector(736, 16),
4143 => conv_std_logic_vector(752, 16),
4144 => conv_std_logic_vector(768, 16),
4145 => conv_std_logic_vector(784, 16),
4146 => conv_std_logic_vector(800, 16),
4147 => conv_std_logic_vector(816, 16),
4148 => conv_std_logic_vector(832, 16),
4149 => conv_std_logic_vector(848, 16),
4150 => conv_std_logic_vector(864, 16),
4151 => conv_std_logic_vector(880, 16),
4152 => conv_std_logic_vector(896, 16),
4153 => conv_std_logic_vector(912, 16),
4154 => conv_std_logic_vector(928, 16),
4155 => conv_std_logic_vector(944, 16),
4156 => conv_std_logic_vector(960, 16),
4157 => conv_std_logic_vector(976, 16),
4158 => conv_std_logic_vector(992, 16),
4159 => conv_std_logic_vector(1008, 16),
4160 => conv_std_logic_vector(1024, 16),
4161 => conv_std_logic_vector(1040, 16),
4162 => conv_std_logic_vector(1056, 16),
4163 => conv_std_logic_vector(1072, 16),
4164 => conv_std_logic_vector(1088, 16),
4165 => conv_std_logic_vector(1104, 16),
4166 => conv_std_logic_vector(1120, 16),
4167 => conv_std_logic_vector(1136, 16),
4168 => conv_std_logic_vector(1152, 16),
4169 => conv_std_logic_vector(1168, 16),
4170 => conv_std_logic_vector(1184, 16),
4171 => conv_std_logic_vector(1200, 16),
4172 => conv_std_logic_vector(1216, 16),
4173 => conv_std_logic_vector(1232, 16),
4174 => conv_std_logic_vector(1248, 16),
4175 => conv_std_logic_vector(1264, 16),
4176 => conv_std_logic_vector(1280, 16),
4177 => conv_std_logic_vector(1296, 16),
4178 => conv_std_logic_vector(1312, 16),
4179 => conv_std_logic_vector(1328, 16),
4180 => conv_std_logic_vector(1344, 16),
4181 => conv_std_logic_vector(1360, 16),
4182 => conv_std_logic_vector(1376, 16),
4183 => conv_std_logic_vector(1392, 16),
4184 => conv_std_logic_vector(1408, 16),
4185 => conv_std_logic_vector(1424, 16),
4186 => conv_std_logic_vector(1440, 16),
4187 => conv_std_logic_vector(1456, 16),
4188 => conv_std_logic_vector(1472, 16),
4189 => conv_std_logic_vector(1488, 16),
4190 => conv_std_logic_vector(1504, 16),
4191 => conv_std_logic_vector(1520, 16),
4192 => conv_std_logic_vector(1536, 16),
4193 => conv_std_logic_vector(1552, 16),
4194 => conv_std_logic_vector(1568, 16),
4195 => conv_std_logic_vector(1584, 16),
4196 => conv_std_logic_vector(1600, 16),
4197 => conv_std_logic_vector(1616, 16),
4198 => conv_std_logic_vector(1632, 16),
4199 => conv_std_logic_vector(1648, 16),
4200 => conv_std_logic_vector(1664, 16),
4201 => conv_std_logic_vector(1680, 16),
4202 => conv_std_logic_vector(1696, 16),
4203 => conv_std_logic_vector(1712, 16),
4204 => conv_std_logic_vector(1728, 16),
4205 => conv_std_logic_vector(1744, 16),
4206 => conv_std_logic_vector(1760, 16),
4207 => conv_std_logic_vector(1776, 16),
4208 => conv_std_logic_vector(1792, 16),
4209 => conv_std_logic_vector(1808, 16),
4210 => conv_std_logic_vector(1824, 16),
4211 => conv_std_logic_vector(1840, 16),
4212 => conv_std_logic_vector(1856, 16),
4213 => conv_std_logic_vector(1872, 16),
4214 => conv_std_logic_vector(1888, 16),
4215 => conv_std_logic_vector(1904, 16),
4216 => conv_std_logic_vector(1920, 16),
4217 => conv_std_logic_vector(1936, 16),
4218 => conv_std_logic_vector(1952, 16),
4219 => conv_std_logic_vector(1968, 16),
4220 => conv_std_logic_vector(1984, 16),
4221 => conv_std_logic_vector(2000, 16),
4222 => conv_std_logic_vector(2016, 16),
4223 => conv_std_logic_vector(2032, 16),
4224 => conv_std_logic_vector(2048, 16),
4225 => conv_std_logic_vector(2064, 16),
4226 => conv_std_logic_vector(2080, 16),
4227 => conv_std_logic_vector(2096, 16),
4228 => conv_std_logic_vector(2112, 16),
4229 => conv_std_logic_vector(2128, 16),
4230 => conv_std_logic_vector(2144, 16),
4231 => conv_std_logic_vector(2160, 16),
4232 => conv_std_logic_vector(2176, 16),
4233 => conv_std_logic_vector(2192, 16),
4234 => conv_std_logic_vector(2208, 16),
4235 => conv_std_logic_vector(2224, 16),
4236 => conv_std_logic_vector(2240, 16),
4237 => conv_std_logic_vector(2256, 16),
4238 => conv_std_logic_vector(2272, 16),
4239 => conv_std_logic_vector(2288, 16),
4240 => conv_std_logic_vector(2304, 16),
4241 => conv_std_logic_vector(2320, 16),
4242 => conv_std_logic_vector(2336, 16),
4243 => conv_std_logic_vector(2352, 16),
4244 => conv_std_logic_vector(2368, 16),
4245 => conv_std_logic_vector(2384, 16),
4246 => conv_std_logic_vector(2400, 16),
4247 => conv_std_logic_vector(2416, 16),
4248 => conv_std_logic_vector(2432, 16),
4249 => conv_std_logic_vector(2448, 16),
4250 => conv_std_logic_vector(2464, 16),
4251 => conv_std_logic_vector(2480, 16),
4252 => conv_std_logic_vector(2496, 16),
4253 => conv_std_logic_vector(2512, 16),
4254 => conv_std_logic_vector(2528, 16),
4255 => conv_std_logic_vector(2544, 16),
4256 => conv_std_logic_vector(2560, 16),
4257 => conv_std_logic_vector(2576, 16),
4258 => conv_std_logic_vector(2592, 16),
4259 => conv_std_logic_vector(2608, 16),
4260 => conv_std_logic_vector(2624, 16),
4261 => conv_std_logic_vector(2640, 16),
4262 => conv_std_logic_vector(2656, 16),
4263 => conv_std_logic_vector(2672, 16),
4264 => conv_std_logic_vector(2688, 16),
4265 => conv_std_logic_vector(2704, 16),
4266 => conv_std_logic_vector(2720, 16),
4267 => conv_std_logic_vector(2736, 16),
4268 => conv_std_logic_vector(2752, 16),
4269 => conv_std_logic_vector(2768, 16),
4270 => conv_std_logic_vector(2784, 16),
4271 => conv_std_logic_vector(2800, 16),
4272 => conv_std_logic_vector(2816, 16),
4273 => conv_std_logic_vector(2832, 16),
4274 => conv_std_logic_vector(2848, 16),
4275 => conv_std_logic_vector(2864, 16),
4276 => conv_std_logic_vector(2880, 16),
4277 => conv_std_logic_vector(2896, 16),
4278 => conv_std_logic_vector(2912, 16),
4279 => conv_std_logic_vector(2928, 16),
4280 => conv_std_logic_vector(2944, 16),
4281 => conv_std_logic_vector(2960, 16),
4282 => conv_std_logic_vector(2976, 16),
4283 => conv_std_logic_vector(2992, 16),
4284 => conv_std_logic_vector(3008, 16),
4285 => conv_std_logic_vector(3024, 16),
4286 => conv_std_logic_vector(3040, 16),
4287 => conv_std_logic_vector(3056, 16),
4288 => conv_std_logic_vector(3072, 16),
4289 => conv_std_logic_vector(3088, 16),
4290 => conv_std_logic_vector(3104, 16),
4291 => conv_std_logic_vector(3120, 16),
4292 => conv_std_logic_vector(3136, 16),
4293 => conv_std_logic_vector(3152, 16),
4294 => conv_std_logic_vector(3168, 16),
4295 => conv_std_logic_vector(3184, 16),
4296 => conv_std_logic_vector(3200, 16),
4297 => conv_std_logic_vector(3216, 16),
4298 => conv_std_logic_vector(3232, 16),
4299 => conv_std_logic_vector(3248, 16),
4300 => conv_std_logic_vector(3264, 16),
4301 => conv_std_logic_vector(3280, 16),
4302 => conv_std_logic_vector(3296, 16),
4303 => conv_std_logic_vector(3312, 16),
4304 => conv_std_logic_vector(3328, 16),
4305 => conv_std_logic_vector(3344, 16),
4306 => conv_std_logic_vector(3360, 16),
4307 => conv_std_logic_vector(3376, 16),
4308 => conv_std_logic_vector(3392, 16),
4309 => conv_std_logic_vector(3408, 16),
4310 => conv_std_logic_vector(3424, 16),
4311 => conv_std_logic_vector(3440, 16),
4312 => conv_std_logic_vector(3456, 16),
4313 => conv_std_logic_vector(3472, 16),
4314 => conv_std_logic_vector(3488, 16),
4315 => conv_std_logic_vector(3504, 16),
4316 => conv_std_logic_vector(3520, 16),
4317 => conv_std_logic_vector(3536, 16),
4318 => conv_std_logic_vector(3552, 16),
4319 => conv_std_logic_vector(3568, 16),
4320 => conv_std_logic_vector(3584, 16),
4321 => conv_std_logic_vector(3600, 16),
4322 => conv_std_logic_vector(3616, 16),
4323 => conv_std_logic_vector(3632, 16),
4324 => conv_std_logic_vector(3648, 16),
4325 => conv_std_logic_vector(3664, 16),
4326 => conv_std_logic_vector(3680, 16),
4327 => conv_std_logic_vector(3696, 16),
4328 => conv_std_logic_vector(3712, 16),
4329 => conv_std_logic_vector(3728, 16),
4330 => conv_std_logic_vector(3744, 16),
4331 => conv_std_logic_vector(3760, 16),
4332 => conv_std_logic_vector(3776, 16),
4333 => conv_std_logic_vector(3792, 16),
4334 => conv_std_logic_vector(3808, 16),
4335 => conv_std_logic_vector(3824, 16),
4336 => conv_std_logic_vector(3840, 16),
4337 => conv_std_logic_vector(3856, 16),
4338 => conv_std_logic_vector(3872, 16),
4339 => conv_std_logic_vector(3888, 16),
4340 => conv_std_logic_vector(3904, 16),
4341 => conv_std_logic_vector(3920, 16),
4342 => conv_std_logic_vector(3936, 16),
4343 => conv_std_logic_vector(3952, 16),
4344 => conv_std_logic_vector(3968, 16),
4345 => conv_std_logic_vector(3984, 16),
4346 => conv_std_logic_vector(4000, 16),
4347 => conv_std_logic_vector(4016, 16),
4348 => conv_std_logic_vector(4032, 16),
4349 => conv_std_logic_vector(4048, 16),
4350 => conv_std_logic_vector(4064, 16),
4351 => conv_std_logic_vector(4080, 16),
4352 => conv_std_logic_vector(0, 16),
4353 => conv_std_logic_vector(17, 16),
4354 => conv_std_logic_vector(34, 16),
4355 => conv_std_logic_vector(51, 16),
4356 => conv_std_logic_vector(68, 16),
4357 => conv_std_logic_vector(85, 16),
4358 => conv_std_logic_vector(102, 16),
4359 => conv_std_logic_vector(119, 16),
4360 => conv_std_logic_vector(136, 16),
4361 => conv_std_logic_vector(153, 16),
4362 => conv_std_logic_vector(170, 16),
4363 => conv_std_logic_vector(187, 16),
4364 => conv_std_logic_vector(204, 16),
4365 => conv_std_logic_vector(221, 16),
4366 => conv_std_logic_vector(238, 16),
4367 => conv_std_logic_vector(255, 16),
4368 => conv_std_logic_vector(272, 16),
4369 => conv_std_logic_vector(289, 16),
4370 => conv_std_logic_vector(306, 16),
4371 => conv_std_logic_vector(323, 16),
4372 => conv_std_logic_vector(340, 16),
4373 => conv_std_logic_vector(357, 16),
4374 => conv_std_logic_vector(374, 16),
4375 => conv_std_logic_vector(391, 16),
4376 => conv_std_logic_vector(408, 16),
4377 => conv_std_logic_vector(425, 16),
4378 => conv_std_logic_vector(442, 16),
4379 => conv_std_logic_vector(459, 16),
4380 => conv_std_logic_vector(476, 16),
4381 => conv_std_logic_vector(493, 16),
4382 => conv_std_logic_vector(510, 16),
4383 => conv_std_logic_vector(527, 16),
4384 => conv_std_logic_vector(544, 16),
4385 => conv_std_logic_vector(561, 16),
4386 => conv_std_logic_vector(578, 16),
4387 => conv_std_logic_vector(595, 16),
4388 => conv_std_logic_vector(612, 16),
4389 => conv_std_logic_vector(629, 16),
4390 => conv_std_logic_vector(646, 16),
4391 => conv_std_logic_vector(663, 16),
4392 => conv_std_logic_vector(680, 16),
4393 => conv_std_logic_vector(697, 16),
4394 => conv_std_logic_vector(714, 16),
4395 => conv_std_logic_vector(731, 16),
4396 => conv_std_logic_vector(748, 16),
4397 => conv_std_logic_vector(765, 16),
4398 => conv_std_logic_vector(782, 16),
4399 => conv_std_logic_vector(799, 16),
4400 => conv_std_logic_vector(816, 16),
4401 => conv_std_logic_vector(833, 16),
4402 => conv_std_logic_vector(850, 16),
4403 => conv_std_logic_vector(867, 16),
4404 => conv_std_logic_vector(884, 16),
4405 => conv_std_logic_vector(901, 16),
4406 => conv_std_logic_vector(918, 16),
4407 => conv_std_logic_vector(935, 16),
4408 => conv_std_logic_vector(952, 16),
4409 => conv_std_logic_vector(969, 16),
4410 => conv_std_logic_vector(986, 16),
4411 => conv_std_logic_vector(1003, 16),
4412 => conv_std_logic_vector(1020, 16),
4413 => conv_std_logic_vector(1037, 16),
4414 => conv_std_logic_vector(1054, 16),
4415 => conv_std_logic_vector(1071, 16),
4416 => conv_std_logic_vector(1088, 16),
4417 => conv_std_logic_vector(1105, 16),
4418 => conv_std_logic_vector(1122, 16),
4419 => conv_std_logic_vector(1139, 16),
4420 => conv_std_logic_vector(1156, 16),
4421 => conv_std_logic_vector(1173, 16),
4422 => conv_std_logic_vector(1190, 16),
4423 => conv_std_logic_vector(1207, 16),
4424 => conv_std_logic_vector(1224, 16),
4425 => conv_std_logic_vector(1241, 16),
4426 => conv_std_logic_vector(1258, 16),
4427 => conv_std_logic_vector(1275, 16),
4428 => conv_std_logic_vector(1292, 16),
4429 => conv_std_logic_vector(1309, 16),
4430 => conv_std_logic_vector(1326, 16),
4431 => conv_std_logic_vector(1343, 16),
4432 => conv_std_logic_vector(1360, 16),
4433 => conv_std_logic_vector(1377, 16),
4434 => conv_std_logic_vector(1394, 16),
4435 => conv_std_logic_vector(1411, 16),
4436 => conv_std_logic_vector(1428, 16),
4437 => conv_std_logic_vector(1445, 16),
4438 => conv_std_logic_vector(1462, 16),
4439 => conv_std_logic_vector(1479, 16),
4440 => conv_std_logic_vector(1496, 16),
4441 => conv_std_logic_vector(1513, 16),
4442 => conv_std_logic_vector(1530, 16),
4443 => conv_std_logic_vector(1547, 16),
4444 => conv_std_logic_vector(1564, 16),
4445 => conv_std_logic_vector(1581, 16),
4446 => conv_std_logic_vector(1598, 16),
4447 => conv_std_logic_vector(1615, 16),
4448 => conv_std_logic_vector(1632, 16),
4449 => conv_std_logic_vector(1649, 16),
4450 => conv_std_logic_vector(1666, 16),
4451 => conv_std_logic_vector(1683, 16),
4452 => conv_std_logic_vector(1700, 16),
4453 => conv_std_logic_vector(1717, 16),
4454 => conv_std_logic_vector(1734, 16),
4455 => conv_std_logic_vector(1751, 16),
4456 => conv_std_logic_vector(1768, 16),
4457 => conv_std_logic_vector(1785, 16),
4458 => conv_std_logic_vector(1802, 16),
4459 => conv_std_logic_vector(1819, 16),
4460 => conv_std_logic_vector(1836, 16),
4461 => conv_std_logic_vector(1853, 16),
4462 => conv_std_logic_vector(1870, 16),
4463 => conv_std_logic_vector(1887, 16),
4464 => conv_std_logic_vector(1904, 16),
4465 => conv_std_logic_vector(1921, 16),
4466 => conv_std_logic_vector(1938, 16),
4467 => conv_std_logic_vector(1955, 16),
4468 => conv_std_logic_vector(1972, 16),
4469 => conv_std_logic_vector(1989, 16),
4470 => conv_std_logic_vector(2006, 16),
4471 => conv_std_logic_vector(2023, 16),
4472 => conv_std_logic_vector(2040, 16),
4473 => conv_std_logic_vector(2057, 16),
4474 => conv_std_logic_vector(2074, 16),
4475 => conv_std_logic_vector(2091, 16),
4476 => conv_std_logic_vector(2108, 16),
4477 => conv_std_logic_vector(2125, 16),
4478 => conv_std_logic_vector(2142, 16),
4479 => conv_std_logic_vector(2159, 16),
4480 => conv_std_logic_vector(2176, 16),
4481 => conv_std_logic_vector(2193, 16),
4482 => conv_std_logic_vector(2210, 16),
4483 => conv_std_logic_vector(2227, 16),
4484 => conv_std_logic_vector(2244, 16),
4485 => conv_std_logic_vector(2261, 16),
4486 => conv_std_logic_vector(2278, 16),
4487 => conv_std_logic_vector(2295, 16),
4488 => conv_std_logic_vector(2312, 16),
4489 => conv_std_logic_vector(2329, 16),
4490 => conv_std_logic_vector(2346, 16),
4491 => conv_std_logic_vector(2363, 16),
4492 => conv_std_logic_vector(2380, 16),
4493 => conv_std_logic_vector(2397, 16),
4494 => conv_std_logic_vector(2414, 16),
4495 => conv_std_logic_vector(2431, 16),
4496 => conv_std_logic_vector(2448, 16),
4497 => conv_std_logic_vector(2465, 16),
4498 => conv_std_logic_vector(2482, 16),
4499 => conv_std_logic_vector(2499, 16),
4500 => conv_std_logic_vector(2516, 16),
4501 => conv_std_logic_vector(2533, 16),
4502 => conv_std_logic_vector(2550, 16),
4503 => conv_std_logic_vector(2567, 16),
4504 => conv_std_logic_vector(2584, 16),
4505 => conv_std_logic_vector(2601, 16),
4506 => conv_std_logic_vector(2618, 16),
4507 => conv_std_logic_vector(2635, 16),
4508 => conv_std_logic_vector(2652, 16),
4509 => conv_std_logic_vector(2669, 16),
4510 => conv_std_logic_vector(2686, 16),
4511 => conv_std_logic_vector(2703, 16),
4512 => conv_std_logic_vector(2720, 16),
4513 => conv_std_logic_vector(2737, 16),
4514 => conv_std_logic_vector(2754, 16),
4515 => conv_std_logic_vector(2771, 16),
4516 => conv_std_logic_vector(2788, 16),
4517 => conv_std_logic_vector(2805, 16),
4518 => conv_std_logic_vector(2822, 16),
4519 => conv_std_logic_vector(2839, 16),
4520 => conv_std_logic_vector(2856, 16),
4521 => conv_std_logic_vector(2873, 16),
4522 => conv_std_logic_vector(2890, 16),
4523 => conv_std_logic_vector(2907, 16),
4524 => conv_std_logic_vector(2924, 16),
4525 => conv_std_logic_vector(2941, 16),
4526 => conv_std_logic_vector(2958, 16),
4527 => conv_std_logic_vector(2975, 16),
4528 => conv_std_logic_vector(2992, 16),
4529 => conv_std_logic_vector(3009, 16),
4530 => conv_std_logic_vector(3026, 16),
4531 => conv_std_logic_vector(3043, 16),
4532 => conv_std_logic_vector(3060, 16),
4533 => conv_std_logic_vector(3077, 16),
4534 => conv_std_logic_vector(3094, 16),
4535 => conv_std_logic_vector(3111, 16),
4536 => conv_std_logic_vector(3128, 16),
4537 => conv_std_logic_vector(3145, 16),
4538 => conv_std_logic_vector(3162, 16),
4539 => conv_std_logic_vector(3179, 16),
4540 => conv_std_logic_vector(3196, 16),
4541 => conv_std_logic_vector(3213, 16),
4542 => conv_std_logic_vector(3230, 16),
4543 => conv_std_logic_vector(3247, 16),
4544 => conv_std_logic_vector(3264, 16),
4545 => conv_std_logic_vector(3281, 16),
4546 => conv_std_logic_vector(3298, 16),
4547 => conv_std_logic_vector(3315, 16),
4548 => conv_std_logic_vector(3332, 16),
4549 => conv_std_logic_vector(3349, 16),
4550 => conv_std_logic_vector(3366, 16),
4551 => conv_std_logic_vector(3383, 16),
4552 => conv_std_logic_vector(3400, 16),
4553 => conv_std_logic_vector(3417, 16),
4554 => conv_std_logic_vector(3434, 16),
4555 => conv_std_logic_vector(3451, 16),
4556 => conv_std_logic_vector(3468, 16),
4557 => conv_std_logic_vector(3485, 16),
4558 => conv_std_logic_vector(3502, 16),
4559 => conv_std_logic_vector(3519, 16),
4560 => conv_std_logic_vector(3536, 16),
4561 => conv_std_logic_vector(3553, 16),
4562 => conv_std_logic_vector(3570, 16),
4563 => conv_std_logic_vector(3587, 16),
4564 => conv_std_logic_vector(3604, 16),
4565 => conv_std_logic_vector(3621, 16),
4566 => conv_std_logic_vector(3638, 16),
4567 => conv_std_logic_vector(3655, 16),
4568 => conv_std_logic_vector(3672, 16),
4569 => conv_std_logic_vector(3689, 16),
4570 => conv_std_logic_vector(3706, 16),
4571 => conv_std_logic_vector(3723, 16),
4572 => conv_std_logic_vector(3740, 16),
4573 => conv_std_logic_vector(3757, 16),
4574 => conv_std_logic_vector(3774, 16),
4575 => conv_std_logic_vector(3791, 16),
4576 => conv_std_logic_vector(3808, 16),
4577 => conv_std_logic_vector(3825, 16),
4578 => conv_std_logic_vector(3842, 16),
4579 => conv_std_logic_vector(3859, 16),
4580 => conv_std_logic_vector(3876, 16),
4581 => conv_std_logic_vector(3893, 16),
4582 => conv_std_logic_vector(3910, 16),
4583 => conv_std_logic_vector(3927, 16),
4584 => conv_std_logic_vector(3944, 16),
4585 => conv_std_logic_vector(3961, 16),
4586 => conv_std_logic_vector(3978, 16),
4587 => conv_std_logic_vector(3995, 16),
4588 => conv_std_logic_vector(4012, 16),
4589 => conv_std_logic_vector(4029, 16),
4590 => conv_std_logic_vector(4046, 16),
4591 => conv_std_logic_vector(4063, 16),
4592 => conv_std_logic_vector(4080, 16),
4593 => conv_std_logic_vector(4097, 16),
4594 => conv_std_logic_vector(4114, 16),
4595 => conv_std_logic_vector(4131, 16),
4596 => conv_std_logic_vector(4148, 16),
4597 => conv_std_logic_vector(4165, 16),
4598 => conv_std_logic_vector(4182, 16),
4599 => conv_std_logic_vector(4199, 16),
4600 => conv_std_logic_vector(4216, 16),
4601 => conv_std_logic_vector(4233, 16),
4602 => conv_std_logic_vector(4250, 16),
4603 => conv_std_logic_vector(4267, 16),
4604 => conv_std_logic_vector(4284, 16),
4605 => conv_std_logic_vector(4301, 16),
4606 => conv_std_logic_vector(4318, 16),
4607 => conv_std_logic_vector(4335, 16),
4608 => conv_std_logic_vector(0, 16),
4609 => conv_std_logic_vector(18, 16),
4610 => conv_std_logic_vector(36, 16),
4611 => conv_std_logic_vector(54, 16),
4612 => conv_std_logic_vector(72, 16),
4613 => conv_std_logic_vector(90, 16),
4614 => conv_std_logic_vector(108, 16),
4615 => conv_std_logic_vector(126, 16),
4616 => conv_std_logic_vector(144, 16),
4617 => conv_std_logic_vector(162, 16),
4618 => conv_std_logic_vector(180, 16),
4619 => conv_std_logic_vector(198, 16),
4620 => conv_std_logic_vector(216, 16),
4621 => conv_std_logic_vector(234, 16),
4622 => conv_std_logic_vector(252, 16),
4623 => conv_std_logic_vector(270, 16),
4624 => conv_std_logic_vector(288, 16),
4625 => conv_std_logic_vector(306, 16),
4626 => conv_std_logic_vector(324, 16),
4627 => conv_std_logic_vector(342, 16),
4628 => conv_std_logic_vector(360, 16),
4629 => conv_std_logic_vector(378, 16),
4630 => conv_std_logic_vector(396, 16),
4631 => conv_std_logic_vector(414, 16),
4632 => conv_std_logic_vector(432, 16),
4633 => conv_std_logic_vector(450, 16),
4634 => conv_std_logic_vector(468, 16),
4635 => conv_std_logic_vector(486, 16),
4636 => conv_std_logic_vector(504, 16),
4637 => conv_std_logic_vector(522, 16),
4638 => conv_std_logic_vector(540, 16),
4639 => conv_std_logic_vector(558, 16),
4640 => conv_std_logic_vector(576, 16),
4641 => conv_std_logic_vector(594, 16),
4642 => conv_std_logic_vector(612, 16),
4643 => conv_std_logic_vector(630, 16),
4644 => conv_std_logic_vector(648, 16),
4645 => conv_std_logic_vector(666, 16),
4646 => conv_std_logic_vector(684, 16),
4647 => conv_std_logic_vector(702, 16),
4648 => conv_std_logic_vector(720, 16),
4649 => conv_std_logic_vector(738, 16),
4650 => conv_std_logic_vector(756, 16),
4651 => conv_std_logic_vector(774, 16),
4652 => conv_std_logic_vector(792, 16),
4653 => conv_std_logic_vector(810, 16),
4654 => conv_std_logic_vector(828, 16),
4655 => conv_std_logic_vector(846, 16),
4656 => conv_std_logic_vector(864, 16),
4657 => conv_std_logic_vector(882, 16),
4658 => conv_std_logic_vector(900, 16),
4659 => conv_std_logic_vector(918, 16),
4660 => conv_std_logic_vector(936, 16),
4661 => conv_std_logic_vector(954, 16),
4662 => conv_std_logic_vector(972, 16),
4663 => conv_std_logic_vector(990, 16),
4664 => conv_std_logic_vector(1008, 16),
4665 => conv_std_logic_vector(1026, 16),
4666 => conv_std_logic_vector(1044, 16),
4667 => conv_std_logic_vector(1062, 16),
4668 => conv_std_logic_vector(1080, 16),
4669 => conv_std_logic_vector(1098, 16),
4670 => conv_std_logic_vector(1116, 16),
4671 => conv_std_logic_vector(1134, 16),
4672 => conv_std_logic_vector(1152, 16),
4673 => conv_std_logic_vector(1170, 16),
4674 => conv_std_logic_vector(1188, 16),
4675 => conv_std_logic_vector(1206, 16),
4676 => conv_std_logic_vector(1224, 16),
4677 => conv_std_logic_vector(1242, 16),
4678 => conv_std_logic_vector(1260, 16),
4679 => conv_std_logic_vector(1278, 16),
4680 => conv_std_logic_vector(1296, 16),
4681 => conv_std_logic_vector(1314, 16),
4682 => conv_std_logic_vector(1332, 16),
4683 => conv_std_logic_vector(1350, 16),
4684 => conv_std_logic_vector(1368, 16),
4685 => conv_std_logic_vector(1386, 16),
4686 => conv_std_logic_vector(1404, 16),
4687 => conv_std_logic_vector(1422, 16),
4688 => conv_std_logic_vector(1440, 16),
4689 => conv_std_logic_vector(1458, 16),
4690 => conv_std_logic_vector(1476, 16),
4691 => conv_std_logic_vector(1494, 16),
4692 => conv_std_logic_vector(1512, 16),
4693 => conv_std_logic_vector(1530, 16),
4694 => conv_std_logic_vector(1548, 16),
4695 => conv_std_logic_vector(1566, 16),
4696 => conv_std_logic_vector(1584, 16),
4697 => conv_std_logic_vector(1602, 16),
4698 => conv_std_logic_vector(1620, 16),
4699 => conv_std_logic_vector(1638, 16),
4700 => conv_std_logic_vector(1656, 16),
4701 => conv_std_logic_vector(1674, 16),
4702 => conv_std_logic_vector(1692, 16),
4703 => conv_std_logic_vector(1710, 16),
4704 => conv_std_logic_vector(1728, 16),
4705 => conv_std_logic_vector(1746, 16),
4706 => conv_std_logic_vector(1764, 16),
4707 => conv_std_logic_vector(1782, 16),
4708 => conv_std_logic_vector(1800, 16),
4709 => conv_std_logic_vector(1818, 16),
4710 => conv_std_logic_vector(1836, 16),
4711 => conv_std_logic_vector(1854, 16),
4712 => conv_std_logic_vector(1872, 16),
4713 => conv_std_logic_vector(1890, 16),
4714 => conv_std_logic_vector(1908, 16),
4715 => conv_std_logic_vector(1926, 16),
4716 => conv_std_logic_vector(1944, 16),
4717 => conv_std_logic_vector(1962, 16),
4718 => conv_std_logic_vector(1980, 16),
4719 => conv_std_logic_vector(1998, 16),
4720 => conv_std_logic_vector(2016, 16),
4721 => conv_std_logic_vector(2034, 16),
4722 => conv_std_logic_vector(2052, 16),
4723 => conv_std_logic_vector(2070, 16),
4724 => conv_std_logic_vector(2088, 16),
4725 => conv_std_logic_vector(2106, 16),
4726 => conv_std_logic_vector(2124, 16),
4727 => conv_std_logic_vector(2142, 16),
4728 => conv_std_logic_vector(2160, 16),
4729 => conv_std_logic_vector(2178, 16),
4730 => conv_std_logic_vector(2196, 16),
4731 => conv_std_logic_vector(2214, 16),
4732 => conv_std_logic_vector(2232, 16),
4733 => conv_std_logic_vector(2250, 16),
4734 => conv_std_logic_vector(2268, 16),
4735 => conv_std_logic_vector(2286, 16),
4736 => conv_std_logic_vector(2304, 16),
4737 => conv_std_logic_vector(2322, 16),
4738 => conv_std_logic_vector(2340, 16),
4739 => conv_std_logic_vector(2358, 16),
4740 => conv_std_logic_vector(2376, 16),
4741 => conv_std_logic_vector(2394, 16),
4742 => conv_std_logic_vector(2412, 16),
4743 => conv_std_logic_vector(2430, 16),
4744 => conv_std_logic_vector(2448, 16),
4745 => conv_std_logic_vector(2466, 16),
4746 => conv_std_logic_vector(2484, 16),
4747 => conv_std_logic_vector(2502, 16),
4748 => conv_std_logic_vector(2520, 16),
4749 => conv_std_logic_vector(2538, 16),
4750 => conv_std_logic_vector(2556, 16),
4751 => conv_std_logic_vector(2574, 16),
4752 => conv_std_logic_vector(2592, 16),
4753 => conv_std_logic_vector(2610, 16),
4754 => conv_std_logic_vector(2628, 16),
4755 => conv_std_logic_vector(2646, 16),
4756 => conv_std_logic_vector(2664, 16),
4757 => conv_std_logic_vector(2682, 16),
4758 => conv_std_logic_vector(2700, 16),
4759 => conv_std_logic_vector(2718, 16),
4760 => conv_std_logic_vector(2736, 16),
4761 => conv_std_logic_vector(2754, 16),
4762 => conv_std_logic_vector(2772, 16),
4763 => conv_std_logic_vector(2790, 16),
4764 => conv_std_logic_vector(2808, 16),
4765 => conv_std_logic_vector(2826, 16),
4766 => conv_std_logic_vector(2844, 16),
4767 => conv_std_logic_vector(2862, 16),
4768 => conv_std_logic_vector(2880, 16),
4769 => conv_std_logic_vector(2898, 16),
4770 => conv_std_logic_vector(2916, 16),
4771 => conv_std_logic_vector(2934, 16),
4772 => conv_std_logic_vector(2952, 16),
4773 => conv_std_logic_vector(2970, 16),
4774 => conv_std_logic_vector(2988, 16),
4775 => conv_std_logic_vector(3006, 16),
4776 => conv_std_logic_vector(3024, 16),
4777 => conv_std_logic_vector(3042, 16),
4778 => conv_std_logic_vector(3060, 16),
4779 => conv_std_logic_vector(3078, 16),
4780 => conv_std_logic_vector(3096, 16),
4781 => conv_std_logic_vector(3114, 16),
4782 => conv_std_logic_vector(3132, 16),
4783 => conv_std_logic_vector(3150, 16),
4784 => conv_std_logic_vector(3168, 16),
4785 => conv_std_logic_vector(3186, 16),
4786 => conv_std_logic_vector(3204, 16),
4787 => conv_std_logic_vector(3222, 16),
4788 => conv_std_logic_vector(3240, 16),
4789 => conv_std_logic_vector(3258, 16),
4790 => conv_std_logic_vector(3276, 16),
4791 => conv_std_logic_vector(3294, 16),
4792 => conv_std_logic_vector(3312, 16),
4793 => conv_std_logic_vector(3330, 16),
4794 => conv_std_logic_vector(3348, 16),
4795 => conv_std_logic_vector(3366, 16),
4796 => conv_std_logic_vector(3384, 16),
4797 => conv_std_logic_vector(3402, 16),
4798 => conv_std_logic_vector(3420, 16),
4799 => conv_std_logic_vector(3438, 16),
4800 => conv_std_logic_vector(3456, 16),
4801 => conv_std_logic_vector(3474, 16),
4802 => conv_std_logic_vector(3492, 16),
4803 => conv_std_logic_vector(3510, 16),
4804 => conv_std_logic_vector(3528, 16),
4805 => conv_std_logic_vector(3546, 16),
4806 => conv_std_logic_vector(3564, 16),
4807 => conv_std_logic_vector(3582, 16),
4808 => conv_std_logic_vector(3600, 16),
4809 => conv_std_logic_vector(3618, 16),
4810 => conv_std_logic_vector(3636, 16),
4811 => conv_std_logic_vector(3654, 16),
4812 => conv_std_logic_vector(3672, 16),
4813 => conv_std_logic_vector(3690, 16),
4814 => conv_std_logic_vector(3708, 16),
4815 => conv_std_logic_vector(3726, 16),
4816 => conv_std_logic_vector(3744, 16),
4817 => conv_std_logic_vector(3762, 16),
4818 => conv_std_logic_vector(3780, 16),
4819 => conv_std_logic_vector(3798, 16),
4820 => conv_std_logic_vector(3816, 16),
4821 => conv_std_logic_vector(3834, 16),
4822 => conv_std_logic_vector(3852, 16),
4823 => conv_std_logic_vector(3870, 16),
4824 => conv_std_logic_vector(3888, 16),
4825 => conv_std_logic_vector(3906, 16),
4826 => conv_std_logic_vector(3924, 16),
4827 => conv_std_logic_vector(3942, 16),
4828 => conv_std_logic_vector(3960, 16),
4829 => conv_std_logic_vector(3978, 16),
4830 => conv_std_logic_vector(3996, 16),
4831 => conv_std_logic_vector(4014, 16),
4832 => conv_std_logic_vector(4032, 16),
4833 => conv_std_logic_vector(4050, 16),
4834 => conv_std_logic_vector(4068, 16),
4835 => conv_std_logic_vector(4086, 16),
4836 => conv_std_logic_vector(4104, 16),
4837 => conv_std_logic_vector(4122, 16),
4838 => conv_std_logic_vector(4140, 16),
4839 => conv_std_logic_vector(4158, 16),
4840 => conv_std_logic_vector(4176, 16),
4841 => conv_std_logic_vector(4194, 16),
4842 => conv_std_logic_vector(4212, 16),
4843 => conv_std_logic_vector(4230, 16),
4844 => conv_std_logic_vector(4248, 16),
4845 => conv_std_logic_vector(4266, 16),
4846 => conv_std_logic_vector(4284, 16),
4847 => conv_std_logic_vector(4302, 16),
4848 => conv_std_logic_vector(4320, 16),
4849 => conv_std_logic_vector(4338, 16),
4850 => conv_std_logic_vector(4356, 16),
4851 => conv_std_logic_vector(4374, 16),
4852 => conv_std_logic_vector(4392, 16),
4853 => conv_std_logic_vector(4410, 16),
4854 => conv_std_logic_vector(4428, 16),
4855 => conv_std_logic_vector(4446, 16),
4856 => conv_std_logic_vector(4464, 16),
4857 => conv_std_logic_vector(4482, 16),
4858 => conv_std_logic_vector(4500, 16),
4859 => conv_std_logic_vector(4518, 16),
4860 => conv_std_logic_vector(4536, 16),
4861 => conv_std_logic_vector(4554, 16),
4862 => conv_std_logic_vector(4572, 16),
4863 => conv_std_logic_vector(4590, 16),
4864 => conv_std_logic_vector(0, 16),
4865 => conv_std_logic_vector(19, 16),
4866 => conv_std_logic_vector(38, 16),
4867 => conv_std_logic_vector(57, 16),
4868 => conv_std_logic_vector(76, 16),
4869 => conv_std_logic_vector(95, 16),
4870 => conv_std_logic_vector(114, 16),
4871 => conv_std_logic_vector(133, 16),
4872 => conv_std_logic_vector(152, 16),
4873 => conv_std_logic_vector(171, 16),
4874 => conv_std_logic_vector(190, 16),
4875 => conv_std_logic_vector(209, 16),
4876 => conv_std_logic_vector(228, 16),
4877 => conv_std_logic_vector(247, 16),
4878 => conv_std_logic_vector(266, 16),
4879 => conv_std_logic_vector(285, 16),
4880 => conv_std_logic_vector(304, 16),
4881 => conv_std_logic_vector(323, 16),
4882 => conv_std_logic_vector(342, 16),
4883 => conv_std_logic_vector(361, 16),
4884 => conv_std_logic_vector(380, 16),
4885 => conv_std_logic_vector(399, 16),
4886 => conv_std_logic_vector(418, 16),
4887 => conv_std_logic_vector(437, 16),
4888 => conv_std_logic_vector(456, 16),
4889 => conv_std_logic_vector(475, 16),
4890 => conv_std_logic_vector(494, 16),
4891 => conv_std_logic_vector(513, 16),
4892 => conv_std_logic_vector(532, 16),
4893 => conv_std_logic_vector(551, 16),
4894 => conv_std_logic_vector(570, 16),
4895 => conv_std_logic_vector(589, 16),
4896 => conv_std_logic_vector(608, 16),
4897 => conv_std_logic_vector(627, 16),
4898 => conv_std_logic_vector(646, 16),
4899 => conv_std_logic_vector(665, 16),
4900 => conv_std_logic_vector(684, 16),
4901 => conv_std_logic_vector(703, 16),
4902 => conv_std_logic_vector(722, 16),
4903 => conv_std_logic_vector(741, 16),
4904 => conv_std_logic_vector(760, 16),
4905 => conv_std_logic_vector(779, 16),
4906 => conv_std_logic_vector(798, 16),
4907 => conv_std_logic_vector(817, 16),
4908 => conv_std_logic_vector(836, 16),
4909 => conv_std_logic_vector(855, 16),
4910 => conv_std_logic_vector(874, 16),
4911 => conv_std_logic_vector(893, 16),
4912 => conv_std_logic_vector(912, 16),
4913 => conv_std_logic_vector(931, 16),
4914 => conv_std_logic_vector(950, 16),
4915 => conv_std_logic_vector(969, 16),
4916 => conv_std_logic_vector(988, 16),
4917 => conv_std_logic_vector(1007, 16),
4918 => conv_std_logic_vector(1026, 16),
4919 => conv_std_logic_vector(1045, 16),
4920 => conv_std_logic_vector(1064, 16),
4921 => conv_std_logic_vector(1083, 16),
4922 => conv_std_logic_vector(1102, 16),
4923 => conv_std_logic_vector(1121, 16),
4924 => conv_std_logic_vector(1140, 16),
4925 => conv_std_logic_vector(1159, 16),
4926 => conv_std_logic_vector(1178, 16),
4927 => conv_std_logic_vector(1197, 16),
4928 => conv_std_logic_vector(1216, 16),
4929 => conv_std_logic_vector(1235, 16),
4930 => conv_std_logic_vector(1254, 16),
4931 => conv_std_logic_vector(1273, 16),
4932 => conv_std_logic_vector(1292, 16),
4933 => conv_std_logic_vector(1311, 16),
4934 => conv_std_logic_vector(1330, 16),
4935 => conv_std_logic_vector(1349, 16),
4936 => conv_std_logic_vector(1368, 16),
4937 => conv_std_logic_vector(1387, 16),
4938 => conv_std_logic_vector(1406, 16),
4939 => conv_std_logic_vector(1425, 16),
4940 => conv_std_logic_vector(1444, 16),
4941 => conv_std_logic_vector(1463, 16),
4942 => conv_std_logic_vector(1482, 16),
4943 => conv_std_logic_vector(1501, 16),
4944 => conv_std_logic_vector(1520, 16),
4945 => conv_std_logic_vector(1539, 16),
4946 => conv_std_logic_vector(1558, 16),
4947 => conv_std_logic_vector(1577, 16),
4948 => conv_std_logic_vector(1596, 16),
4949 => conv_std_logic_vector(1615, 16),
4950 => conv_std_logic_vector(1634, 16),
4951 => conv_std_logic_vector(1653, 16),
4952 => conv_std_logic_vector(1672, 16),
4953 => conv_std_logic_vector(1691, 16),
4954 => conv_std_logic_vector(1710, 16),
4955 => conv_std_logic_vector(1729, 16),
4956 => conv_std_logic_vector(1748, 16),
4957 => conv_std_logic_vector(1767, 16),
4958 => conv_std_logic_vector(1786, 16),
4959 => conv_std_logic_vector(1805, 16),
4960 => conv_std_logic_vector(1824, 16),
4961 => conv_std_logic_vector(1843, 16),
4962 => conv_std_logic_vector(1862, 16),
4963 => conv_std_logic_vector(1881, 16),
4964 => conv_std_logic_vector(1900, 16),
4965 => conv_std_logic_vector(1919, 16),
4966 => conv_std_logic_vector(1938, 16),
4967 => conv_std_logic_vector(1957, 16),
4968 => conv_std_logic_vector(1976, 16),
4969 => conv_std_logic_vector(1995, 16),
4970 => conv_std_logic_vector(2014, 16),
4971 => conv_std_logic_vector(2033, 16),
4972 => conv_std_logic_vector(2052, 16),
4973 => conv_std_logic_vector(2071, 16),
4974 => conv_std_logic_vector(2090, 16),
4975 => conv_std_logic_vector(2109, 16),
4976 => conv_std_logic_vector(2128, 16),
4977 => conv_std_logic_vector(2147, 16),
4978 => conv_std_logic_vector(2166, 16),
4979 => conv_std_logic_vector(2185, 16),
4980 => conv_std_logic_vector(2204, 16),
4981 => conv_std_logic_vector(2223, 16),
4982 => conv_std_logic_vector(2242, 16),
4983 => conv_std_logic_vector(2261, 16),
4984 => conv_std_logic_vector(2280, 16),
4985 => conv_std_logic_vector(2299, 16),
4986 => conv_std_logic_vector(2318, 16),
4987 => conv_std_logic_vector(2337, 16),
4988 => conv_std_logic_vector(2356, 16),
4989 => conv_std_logic_vector(2375, 16),
4990 => conv_std_logic_vector(2394, 16),
4991 => conv_std_logic_vector(2413, 16),
4992 => conv_std_logic_vector(2432, 16),
4993 => conv_std_logic_vector(2451, 16),
4994 => conv_std_logic_vector(2470, 16),
4995 => conv_std_logic_vector(2489, 16),
4996 => conv_std_logic_vector(2508, 16),
4997 => conv_std_logic_vector(2527, 16),
4998 => conv_std_logic_vector(2546, 16),
4999 => conv_std_logic_vector(2565, 16),
5000 => conv_std_logic_vector(2584, 16),
5001 => conv_std_logic_vector(2603, 16),
5002 => conv_std_logic_vector(2622, 16),
5003 => conv_std_logic_vector(2641, 16),
5004 => conv_std_logic_vector(2660, 16),
5005 => conv_std_logic_vector(2679, 16),
5006 => conv_std_logic_vector(2698, 16),
5007 => conv_std_logic_vector(2717, 16),
5008 => conv_std_logic_vector(2736, 16),
5009 => conv_std_logic_vector(2755, 16),
5010 => conv_std_logic_vector(2774, 16),
5011 => conv_std_logic_vector(2793, 16),
5012 => conv_std_logic_vector(2812, 16),
5013 => conv_std_logic_vector(2831, 16),
5014 => conv_std_logic_vector(2850, 16),
5015 => conv_std_logic_vector(2869, 16),
5016 => conv_std_logic_vector(2888, 16),
5017 => conv_std_logic_vector(2907, 16),
5018 => conv_std_logic_vector(2926, 16),
5019 => conv_std_logic_vector(2945, 16),
5020 => conv_std_logic_vector(2964, 16),
5021 => conv_std_logic_vector(2983, 16),
5022 => conv_std_logic_vector(3002, 16),
5023 => conv_std_logic_vector(3021, 16),
5024 => conv_std_logic_vector(3040, 16),
5025 => conv_std_logic_vector(3059, 16),
5026 => conv_std_logic_vector(3078, 16),
5027 => conv_std_logic_vector(3097, 16),
5028 => conv_std_logic_vector(3116, 16),
5029 => conv_std_logic_vector(3135, 16),
5030 => conv_std_logic_vector(3154, 16),
5031 => conv_std_logic_vector(3173, 16),
5032 => conv_std_logic_vector(3192, 16),
5033 => conv_std_logic_vector(3211, 16),
5034 => conv_std_logic_vector(3230, 16),
5035 => conv_std_logic_vector(3249, 16),
5036 => conv_std_logic_vector(3268, 16),
5037 => conv_std_logic_vector(3287, 16),
5038 => conv_std_logic_vector(3306, 16),
5039 => conv_std_logic_vector(3325, 16),
5040 => conv_std_logic_vector(3344, 16),
5041 => conv_std_logic_vector(3363, 16),
5042 => conv_std_logic_vector(3382, 16),
5043 => conv_std_logic_vector(3401, 16),
5044 => conv_std_logic_vector(3420, 16),
5045 => conv_std_logic_vector(3439, 16),
5046 => conv_std_logic_vector(3458, 16),
5047 => conv_std_logic_vector(3477, 16),
5048 => conv_std_logic_vector(3496, 16),
5049 => conv_std_logic_vector(3515, 16),
5050 => conv_std_logic_vector(3534, 16),
5051 => conv_std_logic_vector(3553, 16),
5052 => conv_std_logic_vector(3572, 16),
5053 => conv_std_logic_vector(3591, 16),
5054 => conv_std_logic_vector(3610, 16),
5055 => conv_std_logic_vector(3629, 16),
5056 => conv_std_logic_vector(3648, 16),
5057 => conv_std_logic_vector(3667, 16),
5058 => conv_std_logic_vector(3686, 16),
5059 => conv_std_logic_vector(3705, 16),
5060 => conv_std_logic_vector(3724, 16),
5061 => conv_std_logic_vector(3743, 16),
5062 => conv_std_logic_vector(3762, 16),
5063 => conv_std_logic_vector(3781, 16),
5064 => conv_std_logic_vector(3800, 16),
5065 => conv_std_logic_vector(3819, 16),
5066 => conv_std_logic_vector(3838, 16),
5067 => conv_std_logic_vector(3857, 16),
5068 => conv_std_logic_vector(3876, 16),
5069 => conv_std_logic_vector(3895, 16),
5070 => conv_std_logic_vector(3914, 16),
5071 => conv_std_logic_vector(3933, 16),
5072 => conv_std_logic_vector(3952, 16),
5073 => conv_std_logic_vector(3971, 16),
5074 => conv_std_logic_vector(3990, 16),
5075 => conv_std_logic_vector(4009, 16),
5076 => conv_std_logic_vector(4028, 16),
5077 => conv_std_logic_vector(4047, 16),
5078 => conv_std_logic_vector(4066, 16),
5079 => conv_std_logic_vector(4085, 16),
5080 => conv_std_logic_vector(4104, 16),
5081 => conv_std_logic_vector(4123, 16),
5082 => conv_std_logic_vector(4142, 16),
5083 => conv_std_logic_vector(4161, 16),
5084 => conv_std_logic_vector(4180, 16),
5085 => conv_std_logic_vector(4199, 16),
5086 => conv_std_logic_vector(4218, 16),
5087 => conv_std_logic_vector(4237, 16),
5088 => conv_std_logic_vector(4256, 16),
5089 => conv_std_logic_vector(4275, 16),
5090 => conv_std_logic_vector(4294, 16),
5091 => conv_std_logic_vector(4313, 16),
5092 => conv_std_logic_vector(4332, 16),
5093 => conv_std_logic_vector(4351, 16),
5094 => conv_std_logic_vector(4370, 16),
5095 => conv_std_logic_vector(4389, 16),
5096 => conv_std_logic_vector(4408, 16),
5097 => conv_std_logic_vector(4427, 16),
5098 => conv_std_logic_vector(4446, 16),
5099 => conv_std_logic_vector(4465, 16),
5100 => conv_std_logic_vector(4484, 16),
5101 => conv_std_logic_vector(4503, 16),
5102 => conv_std_logic_vector(4522, 16),
5103 => conv_std_logic_vector(4541, 16),
5104 => conv_std_logic_vector(4560, 16),
5105 => conv_std_logic_vector(4579, 16),
5106 => conv_std_logic_vector(4598, 16),
5107 => conv_std_logic_vector(4617, 16),
5108 => conv_std_logic_vector(4636, 16),
5109 => conv_std_logic_vector(4655, 16),
5110 => conv_std_logic_vector(4674, 16),
5111 => conv_std_logic_vector(4693, 16),
5112 => conv_std_logic_vector(4712, 16),
5113 => conv_std_logic_vector(4731, 16),
5114 => conv_std_logic_vector(4750, 16),
5115 => conv_std_logic_vector(4769, 16),
5116 => conv_std_logic_vector(4788, 16),
5117 => conv_std_logic_vector(4807, 16),
5118 => conv_std_logic_vector(4826, 16),
5119 => conv_std_logic_vector(4845, 16),
5120 => conv_std_logic_vector(0, 16),
5121 => conv_std_logic_vector(20, 16),
5122 => conv_std_logic_vector(40, 16),
5123 => conv_std_logic_vector(60, 16),
5124 => conv_std_logic_vector(80, 16),
5125 => conv_std_logic_vector(100, 16),
5126 => conv_std_logic_vector(120, 16),
5127 => conv_std_logic_vector(140, 16),
5128 => conv_std_logic_vector(160, 16),
5129 => conv_std_logic_vector(180, 16),
5130 => conv_std_logic_vector(200, 16),
5131 => conv_std_logic_vector(220, 16),
5132 => conv_std_logic_vector(240, 16),
5133 => conv_std_logic_vector(260, 16),
5134 => conv_std_logic_vector(280, 16),
5135 => conv_std_logic_vector(300, 16),
5136 => conv_std_logic_vector(320, 16),
5137 => conv_std_logic_vector(340, 16),
5138 => conv_std_logic_vector(360, 16),
5139 => conv_std_logic_vector(380, 16),
5140 => conv_std_logic_vector(400, 16),
5141 => conv_std_logic_vector(420, 16),
5142 => conv_std_logic_vector(440, 16),
5143 => conv_std_logic_vector(460, 16),
5144 => conv_std_logic_vector(480, 16),
5145 => conv_std_logic_vector(500, 16),
5146 => conv_std_logic_vector(520, 16),
5147 => conv_std_logic_vector(540, 16),
5148 => conv_std_logic_vector(560, 16),
5149 => conv_std_logic_vector(580, 16),
5150 => conv_std_logic_vector(600, 16),
5151 => conv_std_logic_vector(620, 16),
5152 => conv_std_logic_vector(640, 16),
5153 => conv_std_logic_vector(660, 16),
5154 => conv_std_logic_vector(680, 16),
5155 => conv_std_logic_vector(700, 16),
5156 => conv_std_logic_vector(720, 16),
5157 => conv_std_logic_vector(740, 16),
5158 => conv_std_logic_vector(760, 16),
5159 => conv_std_logic_vector(780, 16),
5160 => conv_std_logic_vector(800, 16),
5161 => conv_std_logic_vector(820, 16),
5162 => conv_std_logic_vector(840, 16),
5163 => conv_std_logic_vector(860, 16),
5164 => conv_std_logic_vector(880, 16),
5165 => conv_std_logic_vector(900, 16),
5166 => conv_std_logic_vector(920, 16),
5167 => conv_std_logic_vector(940, 16),
5168 => conv_std_logic_vector(960, 16),
5169 => conv_std_logic_vector(980, 16),
5170 => conv_std_logic_vector(1000, 16),
5171 => conv_std_logic_vector(1020, 16),
5172 => conv_std_logic_vector(1040, 16),
5173 => conv_std_logic_vector(1060, 16),
5174 => conv_std_logic_vector(1080, 16),
5175 => conv_std_logic_vector(1100, 16),
5176 => conv_std_logic_vector(1120, 16),
5177 => conv_std_logic_vector(1140, 16),
5178 => conv_std_logic_vector(1160, 16),
5179 => conv_std_logic_vector(1180, 16),
5180 => conv_std_logic_vector(1200, 16),
5181 => conv_std_logic_vector(1220, 16),
5182 => conv_std_logic_vector(1240, 16),
5183 => conv_std_logic_vector(1260, 16),
5184 => conv_std_logic_vector(1280, 16),
5185 => conv_std_logic_vector(1300, 16),
5186 => conv_std_logic_vector(1320, 16),
5187 => conv_std_logic_vector(1340, 16),
5188 => conv_std_logic_vector(1360, 16),
5189 => conv_std_logic_vector(1380, 16),
5190 => conv_std_logic_vector(1400, 16),
5191 => conv_std_logic_vector(1420, 16),
5192 => conv_std_logic_vector(1440, 16),
5193 => conv_std_logic_vector(1460, 16),
5194 => conv_std_logic_vector(1480, 16),
5195 => conv_std_logic_vector(1500, 16),
5196 => conv_std_logic_vector(1520, 16),
5197 => conv_std_logic_vector(1540, 16),
5198 => conv_std_logic_vector(1560, 16),
5199 => conv_std_logic_vector(1580, 16),
5200 => conv_std_logic_vector(1600, 16),
5201 => conv_std_logic_vector(1620, 16),
5202 => conv_std_logic_vector(1640, 16),
5203 => conv_std_logic_vector(1660, 16),
5204 => conv_std_logic_vector(1680, 16),
5205 => conv_std_logic_vector(1700, 16),
5206 => conv_std_logic_vector(1720, 16),
5207 => conv_std_logic_vector(1740, 16),
5208 => conv_std_logic_vector(1760, 16),
5209 => conv_std_logic_vector(1780, 16),
5210 => conv_std_logic_vector(1800, 16),
5211 => conv_std_logic_vector(1820, 16),
5212 => conv_std_logic_vector(1840, 16),
5213 => conv_std_logic_vector(1860, 16),
5214 => conv_std_logic_vector(1880, 16),
5215 => conv_std_logic_vector(1900, 16),
5216 => conv_std_logic_vector(1920, 16),
5217 => conv_std_logic_vector(1940, 16),
5218 => conv_std_logic_vector(1960, 16),
5219 => conv_std_logic_vector(1980, 16),
5220 => conv_std_logic_vector(2000, 16),
5221 => conv_std_logic_vector(2020, 16),
5222 => conv_std_logic_vector(2040, 16),
5223 => conv_std_logic_vector(2060, 16),
5224 => conv_std_logic_vector(2080, 16),
5225 => conv_std_logic_vector(2100, 16),
5226 => conv_std_logic_vector(2120, 16),
5227 => conv_std_logic_vector(2140, 16),
5228 => conv_std_logic_vector(2160, 16),
5229 => conv_std_logic_vector(2180, 16),
5230 => conv_std_logic_vector(2200, 16),
5231 => conv_std_logic_vector(2220, 16),
5232 => conv_std_logic_vector(2240, 16),
5233 => conv_std_logic_vector(2260, 16),
5234 => conv_std_logic_vector(2280, 16),
5235 => conv_std_logic_vector(2300, 16),
5236 => conv_std_logic_vector(2320, 16),
5237 => conv_std_logic_vector(2340, 16),
5238 => conv_std_logic_vector(2360, 16),
5239 => conv_std_logic_vector(2380, 16),
5240 => conv_std_logic_vector(2400, 16),
5241 => conv_std_logic_vector(2420, 16),
5242 => conv_std_logic_vector(2440, 16),
5243 => conv_std_logic_vector(2460, 16),
5244 => conv_std_logic_vector(2480, 16),
5245 => conv_std_logic_vector(2500, 16),
5246 => conv_std_logic_vector(2520, 16),
5247 => conv_std_logic_vector(2540, 16),
5248 => conv_std_logic_vector(2560, 16),
5249 => conv_std_logic_vector(2580, 16),
5250 => conv_std_logic_vector(2600, 16),
5251 => conv_std_logic_vector(2620, 16),
5252 => conv_std_logic_vector(2640, 16),
5253 => conv_std_logic_vector(2660, 16),
5254 => conv_std_logic_vector(2680, 16),
5255 => conv_std_logic_vector(2700, 16),
5256 => conv_std_logic_vector(2720, 16),
5257 => conv_std_logic_vector(2740, 16),
5258 => conv_std_logic_vector(2760, 16),
5259 => conv_std_logic_vector(2780, 16),
5260 => conv_std_logic_vector(2800, 16),
5261 => conv_std_logic_vector(2820, 16),
5262 => conv_std_logic_vector(2840, 16),
5263 => conv_std_logic_vector(2860, 16),
5264 => conv_std_logic_vector(2880, 16),
5265 => conv_std_logic_vector(2900, 16),
5266 => conv_std_logic_vector(2920, 16),
5267 => conv_std_logic_vector(2940, 16),
5268 => conv_std_logic_vector(2960, 16),
5269 => conv_std_logic_vector(2980, 16),
5270 => conv_std_logic_vector(3000, 16),
5271 => conv_std_logic_vector(3020, 16),
5272 => conv_std_logic_vector(3040, 16),
5273 => conv_std_logic_vector(3060, 16),
5274 => conv_std_logic_vector(3080, 16),
5275 => conv_std_logic_vector(3100, 16),
5276 => conv_std_logic_vector(3120, 16),
5277 => conv_std_logic_vector(3140, 16),
5278 => conv_std_logic_vector(3160, 16),
5279 => conv_std_logic_vector(3180, 16),
5280 => conv_std_logic_vector(3200, 16),
5281 => conv_std_logic_vector(3220, 16),
5282 => conv_std_logic_vector(3240, 16),
5283 => conv_std_logic_vector(3260, 16),
5284 => conv_std_logic_vector(3280, 16),
5285 => conv_std_logic_vector(3300, 16),
5286 => conv_std_logic_vector(3320, 16),
5287 => conv_std_logic_vector(3340, 16),
5288 => conv_std_logic_vector(3360, 16),
5289 => conv_std_logic_vector(3380, 16),
5290 => conv_std_logic_vector(3400, 16),
5291 => conv_std_logic_vector(3420, 16),
5292 => conv_std_logic_vector(3440, 16),
5293 => conv_std_logic_vector(3460, 16),
5294 => conv_std_logic_vector(3480, 16),
5295 => conv_std_logic_vector(3500, 16),
5296 => conv_std_logic_vector(3520, 16),
5297 => conv_std_logic_vector(3540, 16),
5298 => conv_std_logic_vector(3560, 16),
5299 => conv_std_logic_vector(3580, 16),
5300 => conv_std_logic_vector(3600, 16),
5301 => conv_std_logic_vector(3620, 16),
5302 => conv_std_logic_vector(3640, 16),
5303 => conv_std_logic_vector(3660, 16),
5304 => conv_std_logic_vector(3680, 16),
5305 => conv_std_logic_vector(3700, 16),
5306 => conv_std_logic_vector(3720, 16),
5307 => conv_std_logic_vector(3740, 16),
5308 => conv_std_logic_vector(3760, 16),
5309 => conv_std_logic_vector(3780, 16),
5310 => conv_std_logic_vector(3800, 16),
5311 => conv_std_logic_vector(3820, 16),
5312 => conv_std_logic_vector(3840, 16),
5313 => conv_std_logic_vector(3860, 16),
5314 => conv_std_logic_vector(3880, 16),
5315 => conv_std_logic_vector(3900, 16),
5316 => conv_std_logic_vector(3920, 16),
5317 => conv_std_logic_vector(3940, 16),
5318 => conv_std_logic_vector(3960, 16),
5319 => conv_std_logic_vector(3980, 16),
5320 => conv_std_logic_vector(4000, 16),
5321 => conv_std_logic_vector(4020, 16),
5322 => conv_std_logic_vector(4040, 16),
5323 => conv_std_logic_vector(4060, 16),
5324 => conv_std_logic_vector(4080, 16),
5325 => conv_std_logic_vector(4100, 16),
5326 => conv_std_logic_vector(4120, 16),
5327 => conv_std_logic_vector(4140, 16),
5328 => conv_std_logic_vector(4160, 16),
5329 => conv_std_logic_vector(4180, 16),
5330 => conv_std_logic_vector(4200, 16),
5331 => conv_std_logic_vector(4220, 16),
5332 => conv_std_logic_vector(4240, 16),
5333 => conv_std_logic_vector(4260, 16),
5334 => conv_std_logic_vector(4280, 16),
5335 => conv_std_logic_vector(4300, 16),
5336 => conv_std_logic_vector(4320, 16),
5337 => conv_std_logic_vector(4340, 16),
5338 => conv_std_logic_vector(4360, 16),
5339 => conv_std_logic_vector(4380, 16),
5340 => conv_std_logic_vector(4400, 16),
5341 => conv_std_logic_vector(4420, 16),
5342 => conv_std_logic_vector(4440, 16),
5343 => conv_std_logic_vector(4460, 16),
5344 => conv_std_logic_vector(4480, 16),
5345 => conv_std_logic_vector(4500, 16),
5346 => conv_std_logic_vector(4520, 16),
5347 => conv_std_logic_vector(4540, 16),
5348 => conv_std_logic_vector(4560, 16),
5349 => conv_std_logic_vector(4580, 16),
5350 => conv_std_logic_vector(4600, 16),
5351 => conv_std_logic_vector(4620, 16),
5352 => conv_std_logic_vector(4640, 16),
5353 => conv_std_logic_vector(4660, 16),
5354 => conv_std_logic_vector(4680, 16),
5355 => conv_std_logic_vector(4700, 16),
5356 => conv_std_logic_vector(4720, 16),
5357 => conv_std_logic_vector(4740, 16),
5358 => conv_std_logic_vector(4760, 16),
5359 => conv_std_logic_vector(4780, 16),
5360 => conv_std_logic_vector(4800, 16),
5361 => conv_std_logic_vector(4820, 16),
5362 => conv_std_logic_vector(4840, 16),
5363 => conv_std_logic_vector(4860, 16),
5364 => conv_std_logic_vector(4880, 16),
5365 => conv_std_logic_vector(4900, 16),
5366 => conv_std_logic_vector(4920, 16),
5367 => conv_std_logic_vector(4940, 16),
5368 => conv_std_logic_vector(4960, 16),
5369 => conv_std_logic_vector(4980, 16),
5370 => conv_std_logic_vector(5000, 16),
5371 => conv_std_logic_vector(5020, 16),
5372 => conv_std_logic_vector(5040, 16),
5373 => conv_std_logic_vector(5060, 16),
5374 => conv_std_logic_vector(5080, 16),
5375 => conv_std_logic_vector(5100, 16),
5376 => conv_std_logic_vector(0, 16),
5377 => conv_std_logic_vector(21, 16),
5378 => conv_std_logic_vector(42, 16),
5379 => conv_std_logic_vector(63, 16),
5380 => conv_std_logic_vector(84, 16),
5381 => conv_std_logic_vector(105, 16),
5382 => conv_std_logic_vector(126, 16),
5383 => conv_std_logic_vector(147, 16),
5384 => conv_std_logic_vector(168, 16),
5385 => conv_std_logic_vector(189, 16),
5386 => conv_std_logic_vector(210, 16),
5387 => conv_std_logic_vector(231, 16),
5388 => conv_std_logic_vector(252, 16),
5389 => conv_std_logic_vector(273, 16),
5390 => conv_std_logic_vector(294, 16),
5391 => conv_std_logic_vector(315, 16),
5392 => conv_std_logic_vector(336, 16),
5393 => conv_std_logic_vector(357, 16),
5394 => conv_std_logic_vector(378, 16),
5395 => conv_std_logic_vector(399, 16),
5396 => conv_std_logic_vector(420, 16),
5397 => conv_std_logic_vector(441, 16),
5398 => conv_std_logic_vector(462, 16),
5399 => conv_std_logic_vector(483, 16),
5400 => conv_std_logic_vector(504, 16),
5401 => conv_std_logic_vector(525, 16),
5402 => conv_std_logic_vector(546, 16),
5403 => conv_std_logic_vector(567, 16),
5404 => conv_std_logic_vector(588, 16),
5405 => conv_std_logic_vector(609, 16),
5406 => conv_std_logic_vector(630, 16),
5407 => conv_std_logic_vector(651, 16),
5408 => conv_std_logic_vector(672, 16),
5409 => conv_std_logic_vector(693, 16),
5410 => conv_std_logic_vector(714, 16),
5411 => conv_std_logic_vector(735, 16),
5412 => conv_std_logic_vector(756, 16),
5413 => conv_std_logic_vector(777, 16),
5414 => conv_std_logic_vector(798, 16),
5415 => conv_std_logic_vector(819, 16),
5416 => conv_std_logic_vector(840, 16),
5417 => conv_std_logic_vector(861, 16),
5418 => conv_std_logic_vector(882, 16),
5419 => conv_std_logic_vector(903, 16),
5420 => conv_std_logic_vector(924, 16),
5421 => conv_std_logic_vector(945, 16),
5422 => conv_std_logic_vector(966, 16),
5423 => conv_std_logic_vector(987, 16),
5424 => conv_std_logic_vector(1008, 16),
5425 => conv_std_logic_vector(1029, 16),
5426 => conv_std_logic_vector(1050, 16),
5427 => conv_std_logic_vector(1071, 16),
5428 => conv_std_logic_vector(1092, 16),
5429 => conv_std_logic_vector(1113, 16),
5430 => conv_std_logic_vector(1134, 16),
5431 => conv_std_logic_vector(1155, 16),
5432 => conv_std_logic_vector(1176, 16),
5433 => conv_std_logic_vector(1197, 16),
5434 => conv_std_logic_vector(1218, 16),
5435 => conv_std_logic_vector(1239, 16),
5436 => conv_std_logic_vector(1260, 16),
5437 => conv_std_logic_vector(1281, 16),
5438 => conv_std_logic_vector(1302, 16),
5439 => conv_std_logic_vector(1323, 16),
5440 => conv_std_logic_vector(1344, 16),
5441 => conv_std_logic_vector(1365, 16),
5442 => conv_std_logic_vector(1386, 16),
5443 => conv_std_logic_vector(1407, 16),
5444 => conv_std_logic_vector(1428, 16),
5445 => conv_std_logic_vector(1449, 16),
5446 => conv_std_logic_vector(1470, 16),
5447 => conv_std_logic_vector(1491, 16),
5448 => conv_std_logic_vector(1512, 16),
5449 => conv_std_logic_vector(1533, 16),
5450 => conv_std_logic_vector(1554, 16),
5451 => conv_std_logic_vector(1575, 16),
5452 => conv_std_logic_vector(1596, 16),
5453 => conv_std_logic_vector(1617, 16),
5454 => conv_std_logic_vector(1638, 16),
5455 => conv_std_logic_vector(1659, 16),
5456 => conv_std_logic_vector(1680, 16),
5457 => conv_std_logic_vector(1701, 16),
5458 => conv_std_logic_vector(1722, 16),
5459 => conv_std_logic_vector(1743, 16),
5460 => conv_std_logic_vector(1764, 16),
5461 => conv_std_logic_vector(1785, 16),
5462 => conv_std_logic_vector(1806, 16),
5463 => conv_std_logic_vector(1827, 16),
5464 => conv_std_logic_vector(1848, 16),
5465 => conv_std_logic_vector(1869, 16),
5466 => conv_std_logic_vector(1890, 16),
5467 => conv_std_logic_vector(1911, 16),
5468 => conv_std_logic_vector(1932, 16),
5469 => conv_std_logic_vector(1953, 16),
5470 => conv_std_logic_vector(1974, 16),
5471 => conv_std_logic_vector(1995, 16),
5472 => conv_std_logic_vector(2016, 16),
5473 => conv_std_logic_vector(2037, 16),
5474 => conv_std_logic_vector(2058, 16),
5475 => conv_std_logic_vector(2079, 16),
5476 => conv_std_logic_vector(2100, 16),
5477 => conv_std_logic_vector(2121, 16),
5478 => conv_std_logic_vector(2142, 16),
5479 => conv_std_logic_vector(2163, 16),
5480 => conv_std_logic_vector(2184, 16),
5481 => conv_std_logic_vector(2205, 16),
5482 => conv_std_logic_vector(2226, 16),
5483 => conv_std_logic_vector(2247, 16),
5484 => conv_std_logic_vector(2268, 16),
5485 => conv_std_logic_vector(2289, 16),
5486 => conv_std_logic_vector(2310, 16),
5487 => conv_std_logic_vector(2331, 16),
5488 => conv_std_logic_vector(2352, 16),
5489 => conv_std_logic_vector(2373, 16),
5490 => conv_std_logic_vector(2394, 16),
5491 => conv_std_logic_vector(2415, 16),
5492 => conv_std_logic_vector(2436, 16),
5493 => conv_std_logic_vector(2457, 16),
5494 => conv_std_logic_vector(2478, 16),
5495 => conv_std_logic_vector(2499, 16),
5496 => conv_std_logic_vector(2520, 16),
5497 => conv_std_logic_vector(2541, 16),
5498 => conv_std_logic_vector(2562, 16),
5499 => conv_std_logic_vector(2583, 16),
5500 => conv_std_logic_vector(2604, 16),
5501 => conv_std_logic_vector(2625, 16),
5502 => conv_std_logic_vector(2646, 16),
5503 => conv_std_logic_vector(2667, 16),
5504 => conv_std_logic_vector(2688, 16),
5505 => conv_std_logic_vector(2709, 16),
5506 => conv_std_logic_vector(2730, 16),
5507 => conv_std_logic_vector(2751, 16),
5508 => conv_std_logic_vector(2772, 16),
5509 => conv_std_logic_vector(2793, 16),
5510 => conv_std_logic_vector(2814, 16),
5511 => conv_std_logic_vector(2835, 16),
5512 => conv_std_logic_vector(2856, 16),
5513 => conv_std_logic_vector(2877, 16),
5514 => conv_std_logic_vector(2898, 16),
5515 => conv_std_logic_vector(2919, 16),
5516 => conv_std_logic_vector(2940, 16),
5517 => conv_std_logic_vector(2961, 16),
5518 => conv_std_logic_vector(2982, 16),
5519 => conv_std_logic_vector(3003, 16),
5520 => conv_std_logic_vector(3024, 16),
5521 => conv_std_logic_vector(3045, 16),
5522 => conv_std_logic_vector(3066, 16),
5523 => conv_std_logic_vector(3087, 16),
5524 => conv_std_logic_vector(3108, 16),
5525 => conv_std_logic_vector(3129, 16),
5526 => conv_std_logic_vector(3150, 16),
5527 => conv_std_logic_vector(3171, 16),
5528 => conv_std_logic_vector(3192, 16),
5529 => conv_std_logic_vector(3213, 16),
5530 => conv_std_logic_vector(3234, 16),
5531 => conv_std_logic_vector(3255, 16),
5532 => conv_std_logic_vector(3276, 16),
5533 => conv_std_logic_vector(3297, 16),
5534 => conv_std_logic_vector(3318, 16),
5535 => conv_std_logic_vector(3339, 16),
5536 => conv_std_logic_vector(3360, 16),
5537 => conv_std_logic_vector(3381, 16),
5538 => conv_std_logic_vector(3402, 16),
5539 => conv_std_logic_vector(3423, 16),
5540 => conv_std_logic_vector(3444, 16),
5541 => conv_std_logic_vector(3465, 16),
5542 => conv_std_logic_vector(3486, 16),
5543 => conv_std_logic_vector(3507, 16),
5544 => conv_std_logic_vector(3528, 16),
5545 => conv_std_logic_vector(3549, 16),
5546 => conv_std_logic_vector(3570, 16),
5547 => conv_std_logic_vector(3591, 16),
5548 => conv_std_logic_vector(3612, 16),
5549 => conv_std_logic_vector(3633, 16),
5550 => conv_std_logic_vector(3654, 16),
5551 => conv_std_logic_vector(3675, 16),
5552 => conv_std_logic_vector(3696, 16),
5553 => conv_std_logic_vector(3717, 16),
5554 => conv_std_logic_vector(3738, 16),
5555 => conv_std_logic_vector(3759, 16),
5556 => conv_std_logic_vector(3780, 16),
5557 => conv_std_logic_vector(3801, 16),
5558 => conv_std_logic_vector(3822, 16),
5559 => conv_std_logic_vector(3843, 16),
5560 => conv_std_logic_vector(3864, 16),
5561 => conv_std_logic_vector(3885, 16),
5562 => conv_std_logic_vector(3906, 16),
5563 => conv_std_logic_vector(3927, 16),
5564 => conv_std_logic_vector(3948, 16),
5565 => conv_std_logic_vector(3969, 16),
5566 => conv_std_logic_vector(3990, 16),
5567 => conv_std_logic_vector(4011, 16),
5568 => conv_std_logic_vector(4032, 16),
5569 => conv_std_logic_vector(4053, 16),
5570 => conv_std_logic_vector(4074, 16),
5571 => conv_std_logic_vector(4095, 16),
5572 => conv_std_logic_vector(4116, 16),
5573 => conv_std_logic_vector(4137, 16),
5574 => conv_std_logic_vector(4158, 16),
5575 => conv_std_logic_vector(4179, 16),
5576 => conv_std_logic_vector(4200, 16),
5577 => conv_std_logic_vector(4221, 16),
5578 => conv_std_logic_vector(4242, 16),
5579 => conv_std_logic_vector(4263, 16),
5580 => conv_std_logic_vector(4284, 16),
5581 => conv_std_logic_vector(4305, 16),
5582 => conv_std_logic_vector(4326, 16),
5583 => conv_std_logic_vector(4347, 16),
5584 => conv_std_logic_vector(4368, 16),
5585 => conv_std_logic_vector(4389, 16),
5586 => conv_std_logic_vector(4410, 16),
5587 => conv_std_logic_vector(4431, 16),
5588 => conv_std_logic_vector(4452, 16),
5589 => conv_std_logic_vector(4473, 16),
5590 => conv_std_logic_vector(4494, 16),
5591 => conv_std_logic_vector(4515, 16),
5592 => conv_std_logic_vector(4536, 16),
5593 => conv_std_logic_vector(4557, 16),
5594 => conv_std_logic_vector(4578, 16),
5595 => conv_std_logic_vector(4599, 16),
5596 => conv_std_logic_vector(4620, 16),
5597 => conv_std_logic_vector(4641, 16),
5598 => conv_std_logic_vector(4662, 16),
5599 => conv_std_logic_vector(4683, 16),
5600 => conv_std_logic_vector(4704, 16),
5601 => conv_std_logic_vector(4725, 16),
5602 => conv_std_logic_vector(4746, 16),
5603 => conv_std_logic_vector(4767, 16),
5604 => conv_std_logic_vector(4788, 16),
5605 => conv_std_logic_vector(4809, 16),
5606 => conv_std_logic_vector(4830, 16),
5607 => conv_std_logic_vector(4851, 16),
5608 => conv_std_logic_vector(4872, 16),
5609 => conv_std_logic_vector(4893, 16),
5610 => conv_std_logic_vector(4914, 16),
5611 => conv_std_logic_vector(4935, 16),
5612 => conv_std_logic_vector(4956, 16),
5613 => conv_std_logic_vector(4977, 16),
5614 => conv_std_logic_vector(4998, 16),
5615 => conv_std_logic_vector(5019, 16),
5616 => conv_std_logic_vector(5040, 16),
5617 => conv_std_logic_vector(5061, 16),
5618 => conv_std_logic_vector(5082, 16),
5619 => conv_std_logic_vector(5103, 16),
5620 => conv_std_logic_vector(5124, 16),
5621 => conv_std_logic_vector(5145, 16),
5622 => conv_std_logic_vector(5166, 16),
5623 => conv_std_logic_vector(5187, 16),
5624 => conv_std_logic_vector(5208, 16),
5625 => conv_std_logic_vector(5229, 16),
5626 => conv_std_logic_vector(5250, 16),
5627 => conv_std_logic_vector(5271, 16),
5628 => conv_std_logic_vector(5292, 16),
5629 => conv_std_logic_vector(5313, 16),
5630 => conv_std_logic_vector(5334, 16),
5631 => conv_std_logic_vector(5355, 16),
5632 => conv_std_logic_vector(0, 16),
5633 => conv_std_logic_vector(22, 16),
5634 => conv_std_logic_vector(44, 16),
5635 => conv_std_logic_vector(66, 16),
5636 => conv_std_logic_vector(88, 16),
5637 => conv_std_logic_vector(110, 16),
5638 => conv_std_logic_vector(132, 16),
5639 => conv_std_logic_vector(154, 16),
5640 => conv_std_logic_vector(176, 16),
5641 => conv_std_logic_vector(198, 16),
5642 => conv_std_logic_vector(220, 16),
5643 => conv_std_logic_vector(242, 16),
5644 => conv_std_logic_vector(264, 16),
5645 => conv_std_logic_vector(286, 16),
5646 => conv_std_logic_vector(308, 16),
5647 => conv_std_logic_vector(330, 16),
5648 => conv_std_logic_vector(352, 16),
5649 => conv_std_logic_vector(374, 16),
5650 => conv_std_logic_vector(396, 16),
5651 => conv_std_logic_vector(418, 16),
5652 => conv_std_logic_vector(440, 16),
5653 => conv_std_logic_vector(462, 16),
5654 => conv_std_logic_vector(484, 16),
5655 => conv_std_logic_vector(506, 16),
5656 => conv_std_logic_vector(528, 16),
5657 => conv_std_logic_vector(550, 16),
5658 => conv_std_logic_vector(572, 16),
5659 => conv_std_logic_vector(594, 16),
5660 => conv_std_logic_vector(616, 16),
5661 => conv_std_logic_vector(638, 16),
5662 => conv_std_logic_vector(660, 16),
5663 => conv_std_logic_vector(682, 16),
5664 => conv_std_logic_vector(704, 16),
5665 => conv_std_logic_vector(726, 16),
5666 => conv_std_logic_vector(748, 16),
5667 => conv_std_logic_vector(770, 16),
5668 => conv_std_logic_vector(792, 16),
5669 => conv_std_logic_vector(814, 16),
5670 => conv_std_logic_vector(836, 16),
5671 => conv_std_logic_vector(858, 16),
5672 => conv_std_logic_vector(880, 16),
5673 => conv_std_logic_vector(902, 16),
5674 => conv_std_logic_vector(924, 16),
5675 => conv_std_logic_vector(946, 16),
5676 => conv_std_logic_vector(968, 16),
5677 => conv_std_logic_vector(990, 16),
5678 => conv_std_logic_vector(1012, 16),
5679 => conv_std_logic_vector(1034, 16),
5680 => conv_std_logic_vector(1056, 16),
5681 => conv_std_logic_vector(1078, 16),
5682 => conv_std_logic_vector(1100, 16),
5683 => conv_std_logic_vector(1122, 16),
5684 => conv_std_logic_vector(1144, 16),
5685 => conv_std_logic_vector(1166, 16),
5686 => conv_std_logic_vector(1188, 16),
5687 => conv_std_logic_vector(1210, 16),
5688 => conv_std_logic_vector(1232, 16),
5689 => conv_std_logic_vector(1254, 16),
5690 => conv_std_logic_vector(1276, 16),
5691 => conv_std_logic_vector(1298, 16),
5692 => conv_std_logic_vector(1320, 16),
5693 => conv_std_logic_vector(1342, 16),
5694 => conv_std_logic_vector(1364, 16),
5695 => conv_std_logic_vector(1386, 16),
5696 => conv_std_logic_vector(1408, 16),
5697 => conv_std_logic_vector(1430, 16),
5698 => conv_std_logic_vector(1452, 16),
5699 => conv_std_logic_vector(1474, 16),
5700 => conv_std_logic_vector(1496, 16),
5701 => conv_std_logic_vector(1518, 16),
5702 => conv_std_logic_vector(1540, 16),
5703 => conv_std_logic_vector(1562, 16),
5704 => conv_std_logic_vector(1584, 16),
5705 => conv_std_logic_vector(1606, 16),
5706 => conv_std_logic_vector(1628, 16),
5707 => conv_std_logic_vector(1650, 16),
5708 => conv_std_logic_vector(1672, 16),
5709 => conv_std_logic_vector(1694, 16),
5710 => conv_std_logic_vector(1716, 16),
5711 => conv_std_logic_vector(1738, 16),
5712 => conv_std_logic_vector(1760, 16),
5713 => conv_std_logic_vector(1782, 16),
5714 => conv_std_logic_vector(1804, 16),
5715 => conv_std_logic_vector(1826, 16),
5716 => conv_std_logic_vector(1848, 16),
5717 => conv_std_logic_vector(1870, 16),
5718 => conv_std_logic_vector(1892, 16),
5719 => conv_std_logic_vector(1914, 16),
5720 => conv_std_logic_vector(1936, 16),
5721 => conv_std_logic_vector(1958, 16),
5722 => conv_std_logic_vector(1980, 16),
5723 => conv_std_logic_vector(2002, 16),
5724 => conv_std_logic_vector(2024, 16),
5725 => conv_std_logic_vector(2046, 16),
5726 => conv_std_logic_vector(2068, 16),
5727 => conv_std_logic_vector(2090, 16),
5728 => conv_std_logic_vector(2112, 16),
5729 => conv_std_logic_vector(2134, 16),
5730 => conv_std_logic_vector(2156, 16),
5731 => conv_std_logic_vector(2178, 16),
5732 => conv_std_logic_vector(2200, 16),
5733 => conv_std_logic_vector(2222, 16),
5734 => conv_std_logic_vector(2244, 16),
5735 => conv_std_logic_vector(2266, 16),
5736 => conv_std_logic_vector(2288, 16),
5737 => conv_std_logic_vector(2310, 16),
5738 => conv_std_logic_vector(2332, 16),
5739 => conv_std_logic_vector(2354, 16),
5740 => conv_std_logic_vector(2376, 16),
5741 => conv_std_logic_vector(2398, 16),
5742 => conv_std_logic_vector(2420, 16),
5743 => conv_std_logic_vector(2442, 16),
5744 => conv_std_logic_vector(2464, 16),
5745 => conv_std_logic_vector(2486, 16),
5746 => conv_std_logic_vector(2508, 16),
5747 => conv_std_logic_vector(2530, 16),
5748 => conv_std_logic_vector(2552, 16),
5749 => conv_std_logic_vector(2574, 16),
5750 => conv_std_logic_vector(2596, 16),
5751 => conv_std_logic_vector(2618, 16),
5752 => conv_std_logic_vector(2640, 16),
5753 => conv_std_logic_vector(2662, 16),
5754 => conv_std_logic_vector(2684, 16),
5755 => conv_std_logic_vector(2706, 16),
5756 => conv_std_logic_vector(2728, 16),
5757 => conv_std_logic_vector(2750, 16),
5758 => conv_std_logic_vector(2772, 16),
5759 => conv_std_logic_vector(2794, 16),
5760 => conv_std_logic_vector(2816, 16),
5761 => conv_std_logic_vector(2838, 16),
5762 => conv_std_logic_vector(2860, 16),
5763 => conv_std_logic_vector(2882, 16),
5764 => conv_std_logic_vector(2904, 16),
5765 => conv_std_logic_vector(2926, 16),
5766 => conv_std_logic_vector(2948, 16),
5767 => conv_std_logic_vector(2970, 16),
5768 => conv_std_logic_vector(2992, 16),
5769 => conv_std_logic_vector(3014, 16),
5770 => conv_std_logic_vector(3036, 16),
5771 => conv_std_logic_vector(3058, 16),
5772 => conv_std_logic_vector(3080, 16),
5773 => conv_std_logic_vector(3102, 16),
5774 => conv_std_logic_vector(3124, 16),
5775 => conv_std_logic_vector(3146, 16),
5776 => conv_std_logic_vector(3168, 16),
5777 => conv_std_logic_vector(3190, 16),
5778 => conv_std_logic_vector(3212, 16),
5779 => conv_std_logic_vector(3234, 16),
5780 => conv_std_logic_vector(3256, 16),
5781 => conv_std_logic_vector(3278, 16),
5782 => conv_std_logic_vector(3300, 16),
5783 => conv_std_logic_vector(3322, 16),
5784 => conv_std_logic_vector(3344, 16),
5785 => conv_std_logic_vector(3366, 16),
5786 => conv_std_logic_vector(3388, 16),
5787 => conv_std_logic_vector(3410, 16),
5788 => conv_std_logic_vector(3432, 16),
5789 => conv_std_logic_vector(3454, 16),
5790 => conv_std_logic_vector(3476, 16),
5791 => conv_std_logic_vector(3498, 16),
5792 => conv_std_logic_vector(3520, 16),
5793 => conv_std_logic_vector(3542, 16),
5794 => conv_std_logic_vector(3564, 16),
5795 => conv_std_logic_vector(3586, 16),
5796 => conv_std_logic_vector(3608, 16),
5797 => conv_std_logic_vector(3630, 16),
5798 => conv_std_logic_vector(3652, 16),
5799 => conv_std_logic_vector(3674, 16),
5800 => conv_std_logic_vector(3696, 16),
5801 => conv_std_logic_vector(3718, 16),
5802 => conv_std_logic_vector(3740, 16),
5803 => conv_std_logic_vector(3762, 16),
5804 => conv_std_logic_vector(3784, 16),
5805 => conv_std_logic_vector(3806, 16),
5806 => conv_std_logic_vector(3828, 16),
5807 => conv_std_logic_vector(3850, 16),
5808 => conv_std_logic_vector(3872, 16),
5809 => conv_std_logic_vector(3894, 16),
5810 => conv_std_logic_vector(3916, 16),
5811 => conv_std_logic_vector(3938, 16),
5812 => conv_std_logic_vector(3960, 16),
5813 => conv_std_logic_vector(3982, 16),
5814 => conv_std_logic_vector(4004, 16),
5815 => conv_std_logic_vector(4026, 16),
5816 => conv_std_logic_vector(4048, 16),
5817 => conv_std_logic_vector(4070, 16),
5818 => conv_std_logic_vector(4092, 16),
5819 => conv_std_logic_vector(4114, 16),
5820 => conv_std_logic_vector(4136, 16),
5821 => conv_std_logic_vector(4158, 16),
5822 => conv_std_logic_vector(4180, 16),
5823 => conv_std_logic_vector(4202, 16),
5824 => conv_std_logic_vector(4224, 16),
5825 => conv_std_logic_vector(4246, 16),
5826 => conv_std_logic_vector(4268, 16),
5827 => conv_std_logic_vector(4290, 16),
5828 => conv_std_logic_vector(4312, 16),
5829 => conv_std_logic_vector(4334, 16),
5830 => conv_std_logic_vector(4356, 16),
5831 => conv_std_logic_vector(4378, 16),
5832 => conv_std_logic_vector(4400, 16),
5833 => conv_std_logic_vector(4422, 16),
5834 => conv_std_logic_vector(4444, 16),
5835 => conv_std_logic_vector(4466, 16),
5836 => conv_std_logic_vector(4488, 16),
5837 => conv_std_logic_vector(4510, 16),
5838 => conv_std_logic_vector(4532, 16),
5839 => conv_std_logic_vector(4554, 16),
5840 => conv_std_logic_vector(4576, 16),
5841 => conv_std_logic_vector(4598, 16),
5842 => conv_std_logic_vector(4620, 16),
5843 => conv_std_logic_vector(4642, 16),
5844 => conv_std_logic_vector(4664, 16),
5845 => conv_std_logic_vector(4686, 16),
5846 => conv_std_logic_vector(4708, 16),
5847 => conv_std_logic_vector(4730, 16),
5848 => conv_std_logic_vector(4752, 16),
5849 => conv_std_logic_vector(4774, 16),
5850 => conv_std_logic_vector(4796, 16),
5851 => conv_std_logic_vector(4818, 16),
5852 => conv_std_logic_vector(4840, 16),
5853 => conv_std_logic_vector(4862, 16),
5854 => conv_std_logic_vector(4884, 16),
5855 => conv_std_logic_vector(4906, 16),
5856 => conv_std_logic_vector(4928, 16),
5857 => conv_std_logic_vector(4950, 16),
5858 => conv_std_logic_vector(4972, 16),
5859 => conv_std_logic_vector(4994, 16),
5860 => conv_std_logic_vector(5016, 16),
5861 => conv_std_logic_vector(5038, 16),
5862 => conv_std_logic_vector(5060, 16),
5863 => conv_std_logic_vector(5082, 16),
5864 => conv_std_logic_vector(5104, 16),
5865 => conv_std_logic_vector(5126, 16),
5866 => conv_std_logic_vector(5148, 16),
5867 => conv_std_logic_vector(5170, 16),
5868 => conv_std_logic_vector(5192, 16),
5869 => conv_std_logic_vector(5214, 16),
5870 => conv_std_logic_vector(5236, 16),
5871 => conv_std_logic_vector(5258, 16),
5872 => conv_std_logic_vector(5280, 16),
5873 => conv_std_logic_vector(5302, 16),
5874 => conv_std_logic_vector(5324, 16),
5875 => conv_std_logic_vector(5346, 16),
5876 => conv_std_logic_vector(5368, 16),
5877 => conv_std_logic_vector(5390, 16),
5878 => conv_std_logic_vector(5412, 16),
5879 => conv_std_logic_vector(5434, 16),
5880 => conv_std_logic_vector(5456, 16),
5881 => conv_std_logic_vector(5478, 16),
5882 => conv_std_logic_vector(5500, 16),
5883 => conv_std_logic_vector(5522, 16),
5884 => conv_std_logic_vector(5544, 16),
5885 => conv_std_logic_vector(5566, 16),
5886 => conv_std_logic_vector(5588, 16),
5887 => conv_std_logic_vector(5610, 16),
5888 => conv_std_logic_vector(0, 16),
5889 => conv_std_logic_vector(23, 16),
5890 => conv_std_logic_vector(46, 16),
5891 => conv_std_logic_vector(69, 16),
5892 => conv_std_logic_vector(92, 16),
5893 => conv_std_logic_vector(115, 16),
5894 => conv_std_logic_vector(138, 16),
5895 => conv_std_logic_vector(161, 16),
5896 => conv_std_logic_vector(184, 16),
5897 => conv_std_logic_vector(207, 16),
5898 => conv_std_logic_vector(230, 16),
5899 => conv_std_logic_vector(253, 16),
5900 => conv_std_logic_vector(276, 16),
5901 => conv_std_logic_vector(299, 16),
5902 => conv_std_logic_vector(322, 16),
5903 => conv_std_logic_vector(345, 16),
5904 => conv_std_logic_vector(368, 16),
5905 => conv_std_logic_vector(391, 16),
5906 => conv_std_logic_vector(414, 16),
5907 => conv_std_logic_vector(437, 16),
5908 => conv_std_logic_vector(460, 16),
5909 => conv_std_logic_vector(483, 16),
5910 => conv_std_logic_vector(506, 16),
5911 => conv_std_logic_vector(529, 16),
5912 => conv_std_logic_vector(552, 16),
5913 => conv_std_logic_vector(575, 16),
5914 => conv_std_logic_vector(598, 16),
5915 => conv_std_logic_vector(621, 16),
5916 => conv_std_logic_vector(644, 16),
5917 => conv_std_logic_vector(667, 16),
5918 => conv_std_logic_vector(690, 16),
5919 => conv_std_logic_vector(713, 16),
5920 => conv_std_logic_vector(736, 16),
5921 => conv_std_logic_vector(759, 16),
5922 => conv_std_logic_vector(782, 16),
5923 => conv_std_logic_vector(805, 16),
5924 => conv_std_logic_vector(828, 16),
5925 => conv_std_logic_vector(851, 16),
5926 => conv_std_logic_vector(874, 16),
5927 => conv_std_logic_vector(897, 16),
5928 => conv_std_logic_vector(920, 16),
5929 => conv_std_logic_vector(943, 16),
5930 => conv_std_logic_vector(966, 16),
5931 => conv_std_logic_vector(989, 16),
5932 => conv_std_logic_vector(1012, 16),
5933 => conv_std_logic_vector(1035, 16),
5934 => conv_std_logic_vector(1058, 16),
5935 => conv_std_logic_vector(1081, 16),
5936 => conv_std_logic_vector(1104, 16),
5937 => conv_std_logic_vector(1127, 16),
5938 => conv_std_logic_vector(1150, 16),
5939 => conv_std_logic_vector(1173, 16),
5940 => conv_std_logic_vector(1196, 16),
5941 => conv_std_logic_vector(1219, 16),
5942 => conv_std_logic_vector(1242, 16),
5943 => conv_std_logic_vector(1265, 16),
5944 => conv_std_logic_vector(1288, 16),
5945 => conv_std_logic_vector(1311, 16),
5946 => conv_std_logic_vector(1334, 16),
5947 => conv_std_logic_vector(1357, 16),
5948 => conv_std_logic_vector(1380, 16),
5949 => conv_std_logic_vector(1403, 16),
5950 => conv_std_logic_vector(1426, 16),
5951 => conv_std_logic_vector(1449, 16),
5952 => conv_std_logic_vector(1472, 16),
5953 => conv_std_logic_vector(1495, 16),
5954 => conv_std_logic_vector(1518, 16),
5955 => conv_std_logic_vector(1541, 16),
5956 => conv_std_logic_vector(1564, 16),
5957 => conv_std_logic_vector(1587, 16),
5958 => conv_std_logic_vector(1610, 16),
5959 => conv_std_logic_vector(1633, 16),
5960 => conv_std_logic_vector(1656, 16),
5961 => conv_std_logic_vector(1679, 16),
5962 => conv_std_logic_vector(1702, 16),
5963 => conv_std_logic_vector(1725, 16),
5964 => conv_std_logic_vector(1748, 16),
5965 => conv_std_logic_vector(1771, 16),
5966 => conv_std_logic_vector(1794, 16),
5967 => conv_std_logic_vector(1817, 16),
5968 => conv_std_logic_vector(1840, 16),
5969 => conv_std_logic_vector(1863, 16),
5970 => conv_std_logic_vector(1886, 16),
5971 => conv_std_logic_vector(1909, 16),
5972 => conv_std_logic_vector(1932, 16),
5973 => conv_std_logic_vector(1955, 16),
5974 => conv_std_logic_vector(1978, 16),
5975 => conv_std_logic_vector(2001, 16),
5976 => conv_std_logic_vector(2024, 16),
5977 => conv_std_logic_vector(2047, 16),
5978 => conv_std_logic_vector(2070, 16),
5979 => conv_std_logic_vector(2093, 16),
5980 => conv_std_logic_vector(2116, 16),
5981 => conv_std_logic_vector(2139, 16),
5982 => conv_std_logic_vector(2162, 16),
5983 => conv_std_logic_vector(2185, 16),
5984 => conv_std_logic_vector(2208, 16),
5985 => conv_std_logic_vector(2231, 16),
5986 => conv_std_logic_vector(2254, 16),
5987 => conv_std_logic_vector(2277, 16),
5988 => conv_std_logic_vector(2300, 16),
5989 => conv_std_logic_vector(2323, 16),
5990 => conv_std_logic_vector(2346, 16),
5991 => conv_std_logic_vector(2369, 16),
5992 => conv_std_logic_vector(2392, 16),
5993 => conv_std_logic_vector(2415, 16),
5994 => conv_std_logic_vector(2438, 16),
5995 => conv_std_logic_vector(2461, 16),
5996 => conv_std_logic_vector(2484, 16),
5997 => conv_std_logic_vector(2507, 16),
5998 => conv_std_logic_vector(2530, 16),
5999 => conv_std_logic_vector(2553, 16),
6000 => conv_std_logic_vector(2576, 16),
6001 => conv_std_logic_vector(2599, 16),
6002 => conv_std_logic_vector(2622, 16),
6003 => conv_std_logic_vector(2645, 16),
6004 => conv_std_logic_vector(2668, 16),
6005 => conv_std_logic_vector(2691, 16),
6006 => conv_std_logic_vector(2714, 16),
6007 => conv_std_logic_vector(2737, 16),
6008 => conv_std_logic_vector(2760, 16),
6009 => conv_std_logic_vector(2783, 16),
6010 => conv_std_logic_vector(2806, 16),
6011 => conv_std_logic_vector(2829, 16),
6012 => conv_std_logic_vector(2852, 16),
6013 => conv_std_logic_vector(2875, 16),
6014 => conv_std_logic_vector(2898, 16),
6015 => conv_std_logic_vector(2921, 16),
6016 => conv_std_logic_vector(2944, 16),
6017 => conv_std_logic_vector(2967, 16),
6018 => conv_std_logic_vector(2990, 16),
6019 => conv_std_logic_vector(3013, 16),
6020 => conv_std_logic_vector(3036, 16),
6021 => conv_std_logic_vector(3059, 16),
6022 => conv_std_logic_vector(3082, 16),
6023 => conv_std_logic_vector(3105, 16),
6024 => conv_std_logic_vector(3128, 16),
6025 => conv_std_logic_vector(3151, 16),
6026 => conv_std_logic_vector(3174, 16),
6027 => conv_std_logic_vector(3197, 16),
6028 => conv_std_logic_vector(3220, 16),
6029 => conv_std_logic_vector(3243, 16),
6030 => conv_std_logic_vector(3266, 16),
6031 => conv_std_logic_vector(3289, 16),
6032 => conv_std_logic_vector(3312, 16),
6033 => conv_std_logic_vector(3335, 16),
6034 => conv_std_logic_vector(3358, 16),
6035 => conv_std_logic_vector(3381, 16),
6036 => conv_std_logic_vector(3404, 16),
6037 => conv_std_logic_vector(3427, 16),
6038 => conv_std_logic_vector(3450, 16),
6039 => conv_std_logic_vector(3473, 16),
6040 => conv_std_logic_vector(3496, 16),
6041 => conv_std_logic_vector(3519, 16),
6042 => conv_std_logic_vector(3542, 16),
6043 => conv_std_logic_vector(3565, 16),
6044 => conv_std_logic_vector(3588, 16),
6045 => conv_std_logic_vector(3611, 16),
6046 => conv_std_logic_vector(3634, 16),
6047 => conv_std_logic_vector(3657, 16),
6048 => conv_std_logic_vector(3680, 16),
6049 => conv_std_logic_vector(3703, 16),
6050 => conv_std_logic_vector(3726, 16),
6051 => conv_std_logic_vector(3749, 16),
6052 => conv_std_logic_vector(3772, 16),
6053 => conv_std_logic_vector(3795, 16),
6054 => conv_std_logic_vector(3818, 16),
6055 => conv_std_logic_vector(3841, 16),
6056 => conv_std_logic_vector(3864, 16),
6057 => conv_std_logic_vector(3887, 16),
6058 => conv_std_logic_vector(3910, 16),
6059 => conv_std_logic_vector(3933, 16),
6060 => conv_std_logic_vector(3956, 16),
6061 => conv_std_logic_vector(3979, 16),
6062 => conv_std_logic_vector(4002, 16),
6063 => conv_std_logic_vector(4025, 16),
6064 => conv_std_logic_vector(4048, 16),
6065 => conv_std_logic_vector(4071, 16),
6066 => conv_std_logic_vector(4094, 16),
6067 => conv_std_logic_vector(4117, 16),
6068 => conv_std_logic_vector(4140, 16),
6069 => conv_std_logic_vector(4163, 16),
6070 => conv_std_logic_vector(4186, 16),
6071 => conv_std_logic_vector(4209, 16),
6072 => conv_std_logic_vector(4232, 16),
6073 => conv_std_logic_vector(4255, 16),
6074 => conv_std_logic_vector(4278, 16),
6075 => conv_std_logic_vector(4301, 16),
6076 => conv_std_logic_vector(4324, 16),
6077 => conv_std_logic_vector(4347, 16),
6078 => conv_std_logic_vector(4370, 16),
6079 => conv_std_logic_vector(4393, 16),
6080 => conv_std_logic_vector(4416, 16),
6081 => conv_std_logic_vector(4439, 16),
6082 => conv_std_logic_vector(4462, 16),
6083 => conv_std_logic_vector(4485, 16),
6084 => conv_std_logic_vector(4508, 16),
6085 => conv_std_logic_vector(4531, 16),
6086 => conv_std_logic_vector(4554, 16),
6087 => conv_std_logic_vector(4577, 16),
6088 => conv_std_logic_vector(4600, 16),
6089 => conv_std_logic_vector(4623, 16),
6090 => conv_std_logic_vector(4646, 16),
6091 => conv_std_logic_vector(4669, 16),
6092 => conv_std_logic_vector(4692, 16),
6093 => conv_std_logic_vector(4715, 16),
6094 => conv_std_logic_vector(4738, 16),
6095 => conv_std_logic_vector(4761, 16),
6096 => conv_std_logic_vector(4784, 16),
6097 => conv_std_logic_vector(4807, 16),
6098 => conv_std_logic_vector(4830, 16),
6099 => conv_std_logic_vector(4853, 16),
6100 => conv_std_logic_vector(4876, 16),
6101 => conv_std_logic_vector(4899, 16),
6102 => conv_std_logic_vector(4922, 16),
6103 => conv_std_logic_vector(4945, 16),
6104 => conv_std_logic_vector(4968, 16),
6105 => conv_std_logic_vector(4991, 16),
6106 => conv_std_logic_vector(5014, 16),
6107 => conv_std_logic_vector(5037, 16),
6108 => conv_std_logic_vector(5060, 16),
6109 => conv_std_logic_vector(5083, 16),
6110 => conv_std_logic_vector(5106, 16),
6111 => conv_std_logic_vector(5129, 16),
6112 => conv_std_logic_vector(5152, 16),
6113 => conv_std_logic_vector(5175, 16),
6114 => conv_std_logic_vector(5198, 16),
6115 => conv_std_logic_vector(5221, 16),
6116 => conv_std_logic_vector(5244, 16),
6117 => conv_std_logic_vector(5267, 16),
6118 => conv_std_logic_vector(5290, 16),
6119 => conv_std_logic_vector(5313, 16),
6120 => conv_std_logic_vector(5336, 16),
6121 => conv_std_logic_vector(5359, 16),
6122 => conv_std_logic_vector(5382, 16),
6123 => conv_std_logic_vector(5405, 16),
6124 => conv_std_logic_vector(5428, 16),
6125 => conv_std_logic_vector(5451, 16),
6126 => conv_std_logic_vector(5474, 16),
6127 => conv_std_logic_vector(5497, 16),
6128 => conv_std_logic_vector(5520, 16),
6129 => conv_std_logic_vector(5543, 16),
6130 => conv_std_logic_vector(5566, 16),
6131 => conv_std_logic_vector(5589, 16),
6132 => conv_std_logic_vector(5612, 16),
6133 => conv_std_logic_vector(5635, 16),
6134 => conv_std_logic_vector(5658, 16),
6135 => conv_std_logic_vector(5681, 16),
6136 => conv_std_logic_vector(5704, 16),
6137 => conv_std_logic_vector(5727, 16),
6138 => conv_std_logic_vector(5750, 16),
6139 => conv_std_logic_vector(5773, 16),
6140 => conv_std_logic_vector(5796, 16),
6141 => conv_std_logic_vector(5819, 16),
6142 => conv_std_logic_vector(5842, 16),
6143 => conv_std_logic_vector(5865, 16),
6144 => conv_std_logic_vector(0, 16),
6145 => conv_std_logic_vector(24, 16),
6146 => conv_std_logic_vector(48, 16),
6147 => conv_std_logic_vector(72, 16),
6148 => conv_std_logic_vector(96, 16),
6149 => conv_std_logic_vector(120, 16),
6150 => conv_std_logic_vector(144, 16),
6151 => conv_std_logic_vector(168, 16),
6152 => conv_std_logic_vector(192, 16),
6153 => conv_std_logic_vector(216, 16),
6154 => conv_std_logic_vector(240, 16),
6155 => conv_std_logic_vector(264, 16),
6156 => conv_std_logic_vector(288, 16),
6157 => conv_std_logic_vector(312, 16),
6158 => conv_std_logic_vector(336, 16),
6159 => conv_std_logic_vector(360, 16),
6160 => conv_std_logic_vector(384, 16),
6161 => conv_std_logic_vector(408, 16),
6162 => conv_std_logic_vector(432, 16),
6163 => conv_std_logic_vector(456, 16),
6164 => conv_std_logic_vector(480, 16),
6165 => conv_std_logic_vector(504, 16),
6166 => conv_std_logic_vector(528, 16),
6167 => conv_std_logic_vector(552, 16),
6168 => conv_std_logic_vector(576, 16),
6169 => conv_std_logic_vector(600, 16),
6170 => conv_std_logic_vector(624, 16),
6171 => conv_std_logic_vector(648, 16),
6172 => conv_std_logic_vector(672, 16),
6173 => conv_std_logic_vector(696, 16),
6174 => conv_std_logic_vector(720, 16),
6175 => conv_std_logic_vector(744, 16),
6176 => conv_std_logic_vector(768, 16),
6177 => conv_std_logic_vector(792, 16),
6178 => conv_std_logic_vector(816, 16),
6179 => conv_std_logic_vector(840, 16),
6180 => conv_std_logic_vector(864, 16),
6181 => conv_std_logic_vector(888, 16),
6182 => conv_std_logic_vector(912, 16),
6183 => conv_std_logic_vector(936, 16),
6184 => conv_std_logic_vector(960, 16),
6185 => conv_std_logic_vector(984, 16),
6186 => conv_std_logic_vector(1008, 16),
6187 => conv_std_logic_vector(1032, 16),
6188 => conv_std_logic_vector(1056, 16),
6189 => conv_std_logic_vector(1080, 16),
6190 => conv_std_logic_vector(1104, 16),
6191 => conv_std_logic_vector(1128, 16),
6192 => conv_std_logic_vector(1152, 16),
6193 => conv_std_logic_vector(1176, 16),
6194 => conv_std_logic_vector(1200, 16),
6195 => conv_std_logic_vector(1224, 16),
6196 => conv_std_logic_vector(1248, 16),
6197 => conv_std_logic_vector(1272, 16),
6198 => conv_std_logic_vector(1296, 16),
6199 => conv_std_logic_vector(1320, 16),
6200 => conv_std_logic_vector(1344, 16),
6201 => conv_std_logic_vector(1368, 16),
6202 => conv_std_logic_vector(1392, 16),
6203 => conv_std_logic_vector(1416, 16),
6204 => conv_std_logic_vector(1440, 16),
6205 => conv_std_logic_vector(1464, 16),
6206 => conv_std_logic_vector(1488, 16),
6207 => conv_std_logic_vector(1512, 16),
6208 => conv_std_logic_vector(1536, 16),
6209 => conv_std_logic_vector(1560, 16),
6210 => conv_std_logic_vector(1584, 16),
6211 => conv_std_logic_vector(1608, 16),
6212 => conv_std_logic_vector(1632, 16),
6213 => conv_std_logic_vector(1656, 16),
6214 => conv_std_logic_vector(1680, 16),
6215 => conv_std_logic_vector(1704, 16),
6216 => conv_std_logic_vector(1728, 16),
6217 => conv_std_logic_vector(1752, 16),
6218 => conv_std_logic_vector(1776, 16),
6219 => conv_std_logic_vector(1800, 16),
6220 => conv_std_logic_vector(1824, 16),
6221 => conv_std_logic_vector(1848, 16),
6222 => conv_std_logic_vector(1872, 16),
6223 => conv_std_logic_vector(1896, 16),
6224 => conv_std_logic_vector(1920, 16),
6225 => conv_std_logic_vector(1944, 16),
6226 => conv_std_logic_vector(1968, 16),
6227 => conv_std_logic_vector(1992, 16),
6228 => conv_std_logic_vector(2016, 16),
6229 => conv_std_logic_vector(2040, 16),
6230 => conv_std_logic_vector(2064, 16),
6231 => conv_std_logic_vector(2088, 16),
6232 => conv_std_logic_vector(2112, 16),
6233 => conv_std_logic_vector(2136, 16),
6234 => conv_std_logic_vector(2160, 16),
6235 => conv_std_logic_vector(2184, 16),
6236 => conv_std_logic_vector(2208, 16),
6237 => conv_std_logic_vector(2232, 16),
6238 => conv_std_logic_vector(2256, 16),
6239 => conv_std_logic_vector(2280, 16),
6240 => conv_std_logic_vector(2304, 16),
6241 => conv_std_logic_vector(2328, 16),
6242 => conv_std_logic_vector(2352, 16),
6243 => conv_std_logic_vector(2376, 16),
6244 => conv_std_logic_vector(2400, 16),
6245 => conv_std_logic_vector(2424, 16),
6246 => conv_std_logic_vector(2448, 16),
6247 => conv_std_logic_vector(2472, 16),
6248 => conv_std_logic_vector(2496, 16),
6249 => conv_std_logic_vector(2520, 16),
6250 => conv_std_logic_vector(2544, 16),
6251 => conv_std_logic_vector(2568, 16),
6252 => conv_std_logic_vector(2592, 16),
6253 => conv_std_logic_vector(2616, 16),
6254 => conv_std_logic_vector(2640, 16),
6255 => conv_std_logic_vector(2664, 16),
6256 => conv_std_logic_vector(2688, 16),
6257 => conv_std_logic_vector(2712, 16),
6258 => conv_std_logic_vector(2736, 16),
6259 => conv_std_logic_vector(2760, 16),
6260 => conv_std_logic_vector(2784, 16),
6261 => conv_std_logic_vector(2808, 16),
6262 => conv_std_logic_vector(2832, 16),
6263 => conv_std_logic_vector(2856, 16),
6264 => conv_std_logic_vector(2880, 16),
6265 => conv_std_logic_vector(2904, 16),
6266 => conv_std_logic_vector(2928, 16),
6267 => conv_std_logic_vector(2952, 16),
6268 => conv_std_logic_vector(2976, 16),
6269 => conv_std_logic_vector(3000, 16),
6270 => conv_std_logic_vector(3024, 16),
6271 => conv_std_logic_vector(3048, 16),
6272 => conv_std_logic_vector(3072, 16),
6273 => conv_std_logic_vector(3096, 16),
6274 => conv_std_logic_vector(3120, 16),
6275 => conv_std_logic_vector(3144, 16),
6276 => conv_std_logic_vector(3168, 16),
6277 => conv_std_logic_vector(3192, 16),
6278 => conv_std_logic_vector(3216, 16),
6279 => conv_std_logic_vector(3240, 16),
6280 => conv_std_logic_vector(3264, 16),
6281 => conv_std_logic_vector(3288, 16),
6282 => conv_std_logic_vector(3312, 16),
6283 => conv_std_logic_vector(3336, 16),
6284 => conv_std_logic_vector(3360, 16),
6285 => conv_std_logic_vector(3384, 16),
6286 => conv_std_logic_vector(3408, 16),
6287 => conv_std_logic_vector(3432, 16),
6288 => conv_std_logic_vector(3456, 16),
6289 => conv_std_logic_vector(3480, 16),
6290 => conv_std_logic_vector(3504, 16),
6291 => conv_std_logic_vector(3528, 16),
6292 => conv_std_logic_vector(3552, 16),
6293 => conv_std_logic_vector(3576, 16),
6294 => conv_std_logic_vector(3600, 16),
6295 => conv_std_logic_vector(3624, 16),
6296 => conv_std_logic_vector(3648, 16),
6297 => conv_std_logic_vector(3672, 16),
6298 => conv_std_logic_vector(3696, 16),
6299 => conv_std_logic_vector(3720, 16),
6300 => conv_std_logic_vector(3744, 16),
6301 => conv_std_logic_vector(3768, 16),
6302 => conv_std_logic_vector(3792, 16),
6303 => conv_std_logic_vector(3816, 16),
6304 => conv_std_logic_vector(3840, 16),
6305 => conv_std_logic_vector(3864, 16),
6306 => conv_std_logic_vector(3888, 16),
6307 => conv_std_logic_vector(3912, 16),
6308 => conv_std_logic_vector(3936, 16),
6309 => conv_std_logic_vector(3960, 16),
6310 => conv_std_logic_vector(3984, 16),
6311 => conv_std_logic_vector(4008, 16),
6312 => conv_std_logic_vector(4032, 16),
6313 => conv_std_logic_vector(4056, 16),
6314 => conv_std_logic_vector(4080, 16),
6315 => conv_std_logic_vector(4104, 16),
6316 => conv_std_logic_vector(4128, 16),
6317 => conv_std_logic_vector(4152, 16),
6318 => conv_std_logic_vector(4176, 16),
6319 => conv_std_logic_vector(4200, 16),
6320 => conv_std_logic_vector(4224, 16),
6321 => conv_std_logic_vector(4248, 16),
6322 => conv_std_logic_vector(4272, 16),
6323 => conv_std_logic_vector(4296, 16),
6324 => conv_std_logic_vector(4320, 16),
6325 => conv_std_logic_vector(4344, 16),
6326 => conv_std_logic_vector(4368, 16),
6327 => conv_std_logic_vector(4392, 16),
6328 => conv_std_logic_vector(4416, 16),
6329 => conv_std_logic_vector(4440, 16),
6330 => conv_std_logic_vector(4464, 16),
6331 => conv_std_logic_vector(4488, 16),
6332 => conv_std_logic_vector(4512, 16),
6333 => conv_std_logic_vector(4536, 16),
6334 => conv_std_logic_vector(4560, 16),
6335 => conv_std_logic_vector(4584, 16),
6336 => conv_std_logic_vector(4608, 16),
6337 => conv_std_logic_vector(4632, 16),
6338 => conv_std_logic_vector(4656, 16),
6339 => conv_std_logic_vector(4680, 16),
6340 => conv_std_logic_vector(4704, 16),
6341 => conv_std_logic_vector(4728, 16),
6342 => conv_std_logic_vector(4752, 16),
6343 => conv_std_logic_vector(4776, 16),
6344 => conv_std_logic_vector(4800, 16),
6345 => conv_std_logic_vector(4824, 16),
6346 => conv_std_logic_vector(4848, 16),
6347 => conv_std_logic_vector(4872, 16),
6348 => conv_std_logic_vector(4896, 16),
6349 => conv_std_logic_vector(4920, 16),
6350 => conv_std_logic_vector(4944, 16),
6351 => conv_std_logic_vector(4968, 16),
6352 => conv_std_logic_vector(4992, 16),
6353 => conv_std_logic_vector(5016, 16),
6354 => conv_std_logic_vector(5040, 16),
6355 => conv_std_logic_vector(5064, 16),
6356 => conv_std_logic_vector(5088, 16),
6357 => conv_std_logic_vector(5112, 16),
6358 => conv_std_logic_vector(5136, 16),
6359 => conv_std_logic_vector(5160, 16),
6360 => conv_std_logic_vector(5184, 16),
6361 => conv_std_logic_vector(5208, 16),
6362 => conv_std_logic_vector(5232, 16),
6363 => conv_std_logic_vector(5256, 16),
6364 => conv_std_logic_vector(5280, 16),
6365 => conv_std_logic_vector(5304, 16),
6366 => conv_std_logic_vector(5328, 16),
6367 => conv_std_logic_vector(5352, 16),
6368 => conv_std_logic_vector(5376, 16),
6369 => conv_std_logic_vector(5400, 16),
6370 => conv_std_logic_vector(5424, 16),
6371 => conv_std_logic_vector(5448, 16),
6372 => conv_std_logic_vector(5472, 16),
6373 => conv_std_logic_vector(5496, 16),
6374 => conv_std_logic_vector(5520, 16),
6375 => conv_std_logic_vector(5544, 16),
6376 => conv_std_logic_vector(5568, 16),
6377 => conv_std_logic_vector(5592, 16),
6378 => conv_std_logic_vector(5616, 16),
6379 => conv_std_logic_vector(5640, 16),
6380 => conv_std_logic_vector(5664, 16),
6381 => conv_std_logic_vector(5688, 16),
6382 => conv_std_logic_vector(5712, 16),
6383 => conv_std_logic_vector(5736, 16),
6384 => conv_std_logic_vector(5760, 16),
6385 => conv_std_logic_vector(5784, 16),
6386 => conv_std_logic_vector(5808, 16),
6387 => conv_std_logic_vector(5832, 16),
6388 => conv_std_logic_vector(5856, 16),
6389 => conv_std_logic_vector(5880, 16),
6390 => conv_std_logic_vector(5904, 16),
6391 => conv_std_logic_vector(5928, 16),
6392 => conv_std_logic_vector(5952, 16),
6393 => conv_std_logic_vector(5976, 16),
6394 => conv_std_logic_vector(6000, 16),
6395 => conv_std_logic_vector(6024, 16),
6396 => conv_std_logic_vector(6048, 16),
6397 => conv_std_logic_vector(6072, 16),
6398 => conv_std_logic_vector(6096, 16),
6399 => conv_std_logic_vector(6120, 16),
6400 => conv_std_logic_vector(0, 16),
6401 => conv_std_logic_vector(25, 16),
6402 => conv_std_logic_vector(50, 16),
6403 => conv_std_logic_vector(75, 16),
6404 => conv_std_logic_vector(100, 16),
6405 => conv_std_logic_vector(125, 16),
6406 => conv_std_logic_vector(150, 16),
6407 => conv_std_logic_vector(175, 16),
6408 => conv_std_logic_vector(200, 16),
6409 => conv_std_logic_vector(225, 16),
6410 => conv_std_logic_vector(250, 16),
6411 => conv_std_logic_vector(275, 16),
6412 => conv_std_logic_vector(300, 16),
6413 => conv_std_logic_vector(325, 16),
6414 => conv_std_logic_vector(350, 16),
6415 => conv_std_logic_vector(375, 16),
6416 => conv_std_logic_vector(400, 16),
6417 => conv_std_logic_vector(425, 16),
6418 => conv_std_logic_vector(450, 16),
6419 => conv_std_logic_vector(475, 16),
6420 => conv_std_logic_vector(500, 16),
6421 => conv_std_logic_vector(525, 16),
6422 => conv_std_logic_vector(550, 16),
6423 => conv_std_logic_vector(575, 16),
6424 => conv_std_logic_vector(600, 16),
6425 => conv_std_logic_vector(625, 16),
6426 => conv_std_logic_vector(650, 16),
6427 => conv_std_logic_vector(675, 16),
6428 => conv_std_logic_vector(700, 16),
6429 => conv_std_logic_vector(725, 16),
6430 => conv_std_logic_vector(750, 16),
6431 => conv_std_logic_vector(775, 16),
6432 => conv_std_logic_vector(800, 16),
6433 => conv_std_logic_vector(825, 16),
6434 => conv_std_logic_vector(850, 16),
6435 => conv_std_logic_vector(875, 16),
6436 => conv_std_logic_vector(900, 16),
6437 => conv_std_logic_vector(925, 16),
6438 => conv_std_logic_vector(950, 16),
6439 => conv_std_logic_vector(975, 16),
6440 => conv_std_logic_vector(1000, 16),
6441 => conv_std_logic_vector(1025, 16),
6442 => conv_std_logic_vector(1050, 16),
6443 => conv_std_logic_vector(1075, 16),
6444 => conv_std_logic_vector(1100, 16),
6445 => conv_std_logic_vector(1125, 16),
6446 => conv_std_logic_vector(1150, 16),
6447 => conv_std_logic_vector(1175, 16),
6448 => conv_std_logic_vector(1200, 16),
6449 => conv_std_logic_vector(1225, 16),
6450 => conv_std_logic_vector(1250, 16),
6451 => conv_std_logic_vector(1275, 16),
6452 => conv_std_logic_vector(1300, 16),
6453 => conv_std_logic_vector(1325, 16),
6454 => conv_std_logic_vector(1350, 16),
6455 => conv_std_logic_vector(1375, 16),
6456 => conv_std_logic_vector(1400, 16),
6457 => conv_std_logic_vector(1425, 16),
6458 => conv_std_logic_vector(1450, 16),
6459 => conv_std_logic_vector(1475, 16),
6460 => conv_std_logic_vector(1500, 16),
6461 => conv_std_logic_vector(1525, 16),
6462 => conv_std_logic_vector(1550, 16),
6463 => conv_std_logic_vector(1575, 16),
6464 => conv_std_logic_vector(1600, 16),
6465 => conv_std_logic_vector(1625, 16),
6466 => conv_std_logic_vector(1650, 16),
6467 => conv_std_logic_vector(1675, 16),
6468 => conv_std_logic_vector(1700, 16),
6469 => conv_std_logic_vector(1725, 16),
6470 => conv_std_logic_vector(1750, 16),
6471 => conv_std_logic_vector(1775, 16),
6472 => conv_std_logic_vector(1800, 16),
6473 => conv_std_logic_vector(1825, 16),
6474 => conv_std_logic_vector(1850, 16),
6475 => conv_std_logic_vector(1875, 16),
6476 => conv_std_logic_vector(1900, 16),
6477 => conv_std_logic_vector(1925, 16),
6478 => conv_std_logic_vector(1950, 16),
6479 => conv_std_logic_vector(1975, 16),
6480 => conv_std_logic_vector(2000, 16),
6481 => conv_std_logic_vector(2025, 16),
6482 => conv_std_logic_vector(2050, 16),
6483 => conv_std_logic_vector(2075, 16),
6484 => conv_std_logic_vector(2100, 16),
6485 => conv_std_logic_vector(2125, 16),
6486 => conv_std_logic_vector(2150, 16),
6487 => conv_std_logic_vector(2175, 16),
6488 => conv_std_logic_vector(2200, 16),
6489 => conv_std_logic_vector(2225, 16),
6490 => conv_std_logic_vector(2250, 16),
6491 => conv_std_logic_vector(2275, 16),
6492 => conv_std_logic_vector(2300, 16),
6493 => conv_std_logic_vector(2325, 16),
6494 => conv_std_logic_vector(2350, 16),
6495 => conv_std_logic_vector(2375, 16),
6496 => conv_std_logic_vector(2400, 16),
6497 => conv_std_logic_vector(2425, 16),
6498 => conv_std_logic_vector(2450, 16),
6499 => conv_std_logic_vector(2475, 16),
6500 => conv_std_logic_vector(2500, 16),
6501 => conv_std_logic_vector(2525, 16),
6502 => conv_std_logic_vector(2550, 16),
6503 => conv_std_logic_vector(2575, 16),
6504 => conv_std_logic_vector(2600, 16),
6505 => conv_std_logic_vector(2625, 16),
6506 => conv_std_logic_vector(2650, 16),
6507 => conv_std_logic_vector(2675, 16),
6508 => conv_std_logic_vector(2700, 16),
6509 => conv_std_logic_vector(2725, 16),
6510 => conv_std_logic_vector(2750, 16),
6511 => conv_std_logic_vector(2775, 16),
6512 => conv_std_logic_vector(2800, 16),
6513 => conv_std_logic_vector(2825, 16),
6514 => conv_std_logic_vector(2850, 16),
6515 => conv_std_logic_vector(2875, 16),
6516 => conv_std_logic_vector(2900, 16),
6517 => conv_std_logic_vector(2925, 16),
6518 => conv_std_logic_vector(2950, 16),
6519 => conv_std_logic_vector(2975, 16),
6520 => conv_std_logic_vector(3000, 16),
6521 => conv_std_logic_vector(3025, 16),
6522 => conv_std_logic_vector(3050, 16),
6523 => conv_std_logic_vector(3075, 16),
6524 => conv_std_logic_vector(3100, 16),
6525 => conv_std_logic_vector(3125, 16),
6526 => conv_std_logic_vector(3150, 16),
6527 => conv_std_logic_vector(3175, 16),
6528 => conv_std_logic_vector(3200, 16),
6529 => conv_std_logic_vector(3225, 16),
6530 => conv_std_logic_vector(3250, 16),
6531 => conv_std_logic_vector(3275, 16),
6532 => conv_std_logic_vector(3300, 16),
6533 => conv_std_logic_vector(3325, 16),
6534 => conv_std_logic_vector(3350, 16),
6535 => conv_std_logic_vector(3375, 16),
6536 => conv_std_logic_vector(3400, 16),
6537 => conv_std_logic_vector(3425, 16),
6538 => conv_std_logic_vector(3450, 16),
6539 => conv_std_logic_vector(3475, 16),
6540 => conv_std_logic_vector(3500, 16),
6541 => conv_std_logic_vector(3525, 16),
6542 => conv_std_logic_vector(3550, 16),
6543 => conv_std_logic_vector(3575, 16),
6544 => conv_std_logic_vector(3600, 16),
6545 => conv_std_logic_vector(3625, 16),
6546 => conv_std_logic_vector(3650, 16),
6547 => conv_std_logic_vector(3675, 16),
6548 => conv_std_logic_vector(3700, 16),
6549 => conv_std_logic_vector(3725, 16),
6550 => conv_std_logic_vector(3750, 16),
6551 => conv_std_logic_vector(3775, 16),
6552 => conv_std_logic_vector(3800, 16),
6553 => conv_std_logic_vector(3825, 16),
6554 => conv_std_logic_vector(3850, 16),
6555 => conv_std_logic_vector(3875, 16),
6556 => conv_std_logic_vector(3900, 16),
6557 => conv_std_logic_vector(3925, 16),
6558 => conv_std_logic_vector(3950, 16),
6559 => conv_std_logic_vector(3975, 16),
6560 => conv_std_logic_vector(4000, 16),
6561 => conv_std_logic_vector(4025, 16),
6562 => conv_std_logic_vector(4050, 16),
6563 => conv_std_logic_vector(4075, 16),
6564 => conv_std_logic_vector(4100, 16),
6565 => conv_std_logic_vector(4125, 16),
6566 => conv_std_logic_vector(4150, 16),
6567 => conv_std_logic_vector(4175, 16),
6568 => conv_std_logic_vector(4200, 16),
6569 => conv_std_logic_vector(4225, 16),
6570 => conv_std_logic_vector(4250, 16),
6571 => conv_std_logic_vector(4275, 16),
6572 => conv_std_logic_vector(4300, 16),
6573 => conv_std_logic_vector(4325, 16),
6574 => conv_std_logic_vector(4350, 16),
6575 => conv_std_logic_vector(4375, 16),
6576 => conv_std_logic_vector(4400, 16),
6577 => conv_std_logic_vector(4425, 16),
6578 => conv_std_logic_vector(4450, 16),
6579 => conv_std_logic_vector(4475, 16),
6580 => conv_std_logic_vector(4500, 16),
6581 => conv_std_logic_vector(4525, 16),
6582 => conv_std_logic_vector(4550, 16),
6583 => conv_std_logic_vector(4575, 16),
6584 => conv_std_logic_vector(4600, 16),
6585 => conv_std_logic_vector(4625, 16),
6586 => conv_std_logic_vector(4650, 16),
6587 => conv_std_logic_vector(4675, 16),
6588 => conv_std_logic_vector(4700, 16),
6589 => conv_std_logic_vector(4725, 16),
6590 => conv_std_logic_vector(4750, 16),
6591 => conv_std_logic_vector(4775, 16),
6592 => conv_std_logic_vector(4800, 16),
6593 => conv_std_logic_vector(4825, 16),
6594 => conv_std_logic_vector(4850, 16),
6595 => conv_std_logic_vector(4875, 16),
6596 => conv_std_logic_vector(4900, 16),
6597 => conv_std_logic_vector(4925, 16),
6598 => conv_std_logic_vector(4950, 16),
6599 => conv_std_logic_vector(4975, 16),
6600 => conv_std_logic_vector(5000, 16),
6601 => conv_std_logic_vector(5025, 16),
6602 => conv_std_logic_vector(5050, 16),
6603 => conv_std_logic_vector(5075, 16),
6604 => conv_std_logic_vector(5100, 16),
6605 => conv_std_logic_vector(5125, 16),
6606 => conv_std_logic_vector(5150, 16),
6607 => conv_std_logic_vector(5175, 16),
6608 => conv_std_logic_vector(5200, 16),
6609 => conv_std_logic_vector(5225, 16),
6610 => conv_std_logic_vector(5250, 16),
6611 => conv_std_logic_vector(5275, 16),
6612 => conv_std_logic_vector(5300, 16),
6613 => conv_std_logic_vector(5325, 16),
6614 => conv_std_logic_vector(5350, 16),
6615 => conv_std_logic_vector(5375, 16),
6616 => conv_std_logic_vector(5400, 16),
6617 => conv_std_logic_vector(5425, 16),
6618 => conv_std_logic_vector(5450, 16),
6619 => conv_std_logic_vector(5475, 16),
6620 => conv_std_logic_vector(5500, 16),
6621 => conv_std_logic_vector(5525, 16),
6622 => conv_std_logic_vector(5550, 16),
6623 => conv_std_logic_vector(5575, 16),
6624 => conv_std_logic_vector(5600, 16),
6625 => conv_std_logic_vector(5625, 16),
6626 => conv_std_logic_vector(5650, 16),
6627 => conv_std_logic_vector(5675, 16),
6628 => conv_std_logic_vector(5700, 16),
6629 => conv_std_logic_vector(5725, 16),
6630 => conv_std_logic_vector(5750, 16),
6631 => conv_std_logic_vector(5775, 16),
6632 => conv_std_logic_vector(5800, 16),
6633 => conv_std_logic_vector(5825, 16),
6634 => conv_std_logic_vector(5850, 16),
6635 => conv_std_logic_vector(5875, 16),
6636 => conv_std_logic_vector(5900, 16),
6637 => conv_std_logic_vector(5925, 16),
6638 => conv_std_logic_vector(5950, 16),
6639 => conv_std_logic_vector(5975, 16),
6640 => conv_std_logic_vector(6000, 16),
6641 => conv_std_logic_vector(6025, 16),
6642 => conv_std_logic_vector(6050, 16),
6643 => conv_std_logic_vector(6075, 16),
6644 => conv_std_logic_vector(6100, 16),
6645 => conv_std_logic_vector(6125, 16),
6646 => conv_std_logic_vector(6150, 16),
6647 => conv_std_logic_vector(6175, 16),
6648 => conv_std_logic_vector(6200, 16),
6649 => conv_std_logic_vector(6225, 16),
6650 => conv_std_logic_vector(6250, 16),
6651 => conv_std_logic_vector(6275, 16),
6652 => conv_std_logic_vector(6300, 16),
6653 => conv_std_logic_vector(6325, 16),
6654 => conv_std_logic_vector(6350, 16),
6655 => conv_std_logic_vector(6375, 16),
6656 => conv_std_logic_vector(0, 16),
6657 => conv_std_logic_vector(26, 16),
6658 => conv_std_logic_vector(52, 16),
6659 => conv_std_logic_vector(78, 16),
6660 => conv_std_logic_vector(104, 16),
6661 => conv_std_logic_vector(130, 16),
6662 => conv_std_logic_vector(156, 16),
6663 => conv_std_logic_vector(182, 16),
6664 => conv_std_logic_vector(208, 16),
6665 => conv_std_logic_vector(234, 16),
6666 => conv_std_logic_vector(260, 16),
6667 => conv_std_logic_vector(286, 16),
6668 => conv_std_logic_vector(312, 16),
6669 => conv_std_logic_vector(338, 16),
6670 => conv_std_logic_vector(364, 16),
6671 => conv_std_logic_vector(390, 16),
6672 => conv_std_logic_vector(416, 16),
6673 => conv_std_logic_vector(442, 16),
6674 => conv_std_logic_vector(468, 16),
6675 => conv_std_logic_vector(494, 16),
6676 => conv_std_logic_vector(520, 16),
6677 => conv_std_logic_vector(546, 16),
6678 => conv_std_logic_vector(572, 16),
6679 => conv_std_logic_vector(598, 16),
6680 => conv_std_logic_vector(624, 16),
6681 => conv_std_logic_vector(650, 16),
6682 => conv_std_logic_vector(676, 16),
6683 => conv_std_logic_vector(702, 16),
6684 => conv_std_logic_vector(728, 16),
6685 => conv_std_logic_vector(754, 16),
6686 => conv_std_logic_vector(780, 16),
6687 => conv_std_logic_vector(806, 16),
6688 => conv_std_logic_vector(832, 16),
6689 => conv_std_logic_vector(858, 16),
6690 => conv_std_logic_vector(884, 16),
6691 => conv_std_logic_vector(910, 16),
6692 => conv_std_logic_vector(936, 16),
6693 => conv_std_logic_vector(962, 16),
6694 => conv_std_logic_vector(988, 16),
6695 => conv_std_logic_vector(1014, 16),
6696 => conv_std_logic_vector(1040, 16),
6697 => conv_std_logic_vector(1066, 16),
6698 => conv_std_logic_vector(1092, 16),
6699 => conv_std_logic_vector(1118, 16),
6700 => conv_std_logic_vector(1144, 16),
6701 => conv_std_logic_vector(1170, 16),
6702 => conv_std_logic_vector(1196, 16),
6703 => conv_std_logic_vector(1222, 16),
6704 => conv_std_logic_vector(1248, 16),
6705 => conv_std_logic_vector(1274, 16),
6706 => conv_std_logic_vector(1300, 16),
6707 => conv_std_logic_vector(1326, 16),
6708 => conv_std_logic_vector(1352, 16),
6709 => conv_std_logic_vector(1378, 16),
6710 => conv_std_logic_vector(1404, 16),
6711 => conv_std_logic_vector(1430, 16),
6712 => conv_std_logic_vector(1456, 16),
6713 => conv_std_logic_vector(1482, 16),
6714 => conv_std_logic_vector(1508, 16),
6715 => conv_std_logic_vector(1534, 16),
6716 => conv_std_logic_vector(1560, 16),
6717 => conv_std_logic_vector(1586, 16),
6718 => conv_std_logic_vector(1612, 16),
6719 => conv_std_logic_vector(1638, 16),
6720 => conv_std_logic_vector(1664, 16),
6721 => conv_std_logic_vector(1690, 16),
6722 => conv_std_logic_vector(1716, 16),
6723 => conv_std_logic_vector(1742, 16),
6724 => conv_std_logic_vector(1768, 16),
6725 => conv_std_logic_vector(1794, 16),
6726 => conv_std_logic_vector(1820, 16),
6727 => conv_std_logic_vector(1846, 16),
6728 => conv_std_logic_vector(1872, 16),
6729 => conv_std_logic_vector(1898, 16),
6730 => conv_std_logic_vector(1924, 16),
6731 => conv_std_logic_vector(1950, 16),
6732 => conv_std_logic_vector(1976, 16),
6733 => conv_std_logic_vector(2002, 16),
6734 => conv_std_logic_vector(2028, 16),
6735 => conv_std_logic_vector(2054, 16),
6736 => conv_std_logic_vector(2080, 16),
6737 => conv_std_logic_vector(2106, 16),
6738 => conv_std_logic_vector(2132, 16),
6739 => conv_std_logic_vector(2158, 16),
6740 => conv_std_logic_vector(2184, 16),
6741 => conv_std_logic_vector(2210, 16),
6742 => conv_std_logic_vector(2236, 16),
6743 => conv_std_logic_vector(2262, 16),
6744 => conv_std_logic_vector(2288, 16),
6745 => conv_std_logic_vector(2314, 16),
6746 => conv_std_logic_vector(2340, 16),
6747 => conv_std_logic_vector(2366, 16),
6748 => conv_std_logic_vector(2392, 16),
6749 => conv_std_logic_vector(2418, 16),
6750 => conv_std_logic_vector(2444, 16),
6751 => conv_std_logic_vector(2470, 16),
6752 => conv_std_logic_vector(2496, 16),
6753 => conv_std_logic_vector(2522, 16),
6754 => conv_std_logic_vector(2548, 16),
6755 => conv_std_logic_vector(2574, 16),
6756 => conv_std_logic_vector(2600, 16),
6757 => conv_std_logic_vector(2626, 16),
6758 => conv_std_logic_vector(2652, 16),
6759 => conv_std_logic_vector(2678, 16),
6760 => conv_std_logic_vector(2704, 16),
6761 => conv_std_logic_vector(2730, 16),
6762 => conv_std_logic_vector(2756, 16),
6763 => conv_std_logic_vector(2782, 16),
6764 => conv_std_logic_vector(2808, 16),
6765 => conv_std_logic_vector(2834, 16),
6766 => conv_std_logic_vector(2860, 16),
6767 => conv_std_logic_vector(2886, 16),
6768 => conv_std_logic_vector(2912, 16),
6769 => conv_std_logic_vector(2938, 16),
6770 => conv_std_logic_vector(2964, 16),
6771 => conv_std_logic_vector(2990, 16),
6772 => conv_std_logic_vector(3016, 16),
6773 => conv_std_logic_vector(3042, 16),
6774 => conv_std_logic_vector(3068, 16),
6775 => conv_std_logic_vector(3094, 16),
6776 => conv_std_logic_vector(3120, 16),
6777 => conv_std_logic_vector(3146, 16),
6778 => conv_std_logic_vector(3172, 16),
6779 => conv_std_logic_vector(3198, 16),
6780 => conv_std_logic_vector(3224, 16),
6781 => conv_std_logic_vector(3250, 16),
6782 => conv_std_logic_vector(3276, 16),
6783 => conv_std_logic_vector(3302, 16),
6784 => conv_std_logic_vector(3328, 16),
6785 => conv_std_logic_vector(3354, 16),
6786 => conv_std_logic_vector(3380, 16),
6787 => conv_std_logic_vector(3406, 16),
6788 => conv_std_logic_vector(3432, 16),
6789 => conv_std_logic_vector(3458, 16),
6790 => conv_std_logic_vector(3484, 16),
6791 => conv_std_logic_vector(3510, 16),
6792 => conv_std_logic_vector(3536, 16),
6793 => conv_std_logic_vector(3562, 16),
6794 => conv_std_logic_vector(3588, 16),
6795 => conv_std_logic_vector(3614, 16),
6796 => conv_std_logic_vector(3640, 16),
6797 => conv_std_logic_vector(3666, 16),
6798 => conv_std_logic_vector(3692, 16),
6799 => conv_std_logic_vector(3718, 16),
6800 => conv_std_logic_vector(3744, 16),
6801 => conv_std_logic_vector(3770, 16),
6802 => conv_std_logic_vector(3796, 16),
6803 => conv_std_logic_vector(3822, 16),
6804 => conv_std_logic_vector(3848, 16),
6805 => conv_std_logic_vector(3874, 16),
6806 => conv_std_logic_vector(3900, 16),
6807 => conv_std_logic_vector(3926, 16),
6808 => conv_std_logic_vector(3952, 16),
6809 => conv_std_logic_vector(3978, 16),
6810 => conv_std_logic_vector(4004, 16),
6811 => conv_std_logic_vector(4030, 16),
6812 => conv_std_logic_vector(4056, 16),
6813 => conv_std_logic_vector(4082, 16),
6814 => conv_std_logic_vector(4108, 16),
6815 => conv_std_logic_vector(4134, 16),
6816 => conv_std_logic_vector(4160, 16),
6817 => conv_std_logic_vector(4186, 16),
6818 => conv_std_logic_vector(4212, 16),
6819 => conv_std_logic_vector(4238, 16),
6820 => conv_std_logic_vector(4264, 16),
6821 => conv_std_logic_vector(4290, 16),
6822 => conv_std_logic_vector(4316, 16),
6823 => conv_std_logic_vector(4342, 16),
6824 => conv_std_logic_vector(4368, 16),
6825 => conv_std_logic_vector(4394, 16),
6826 => conv_std_logic_vector(4420, 16),
6827 => conv_std_logic_vector(4446, 16),
6828 => conv_std_logic_vector(4472, 16),
6829 => conv_std_logic_vector(4498, 16),
6830 => conv_std_logic_vector(4524, 16),
6831 => conv_std_logic_vector(4550, 16),
6832 => conv_std_logic_vector(4576, 16),
6833 => conv_std_logic_vector(4602, 16),
6834 => conv_std_logic_vector(4628, 16),
6835 => conv_std_logic_vector(4654, 16),
6836 => conv_std_logic_vector(4680, 16),
6837 => conv_std_logic_vector(4706, 16),
6838 => conv_std_logic_vector(4732, 16),
6839 => conv_std_logic_vector(4758, 16),
6840 => conv_std_logic_vector(4784, 16),
6841 => conv_std_logic_vector(4810, 16),
6842 => conv_std_logic_vector(4836, 16),
6843 => conv_std_logic_vector(4862, 16),
6844 => conv_std_logic_vector(4888, 16),
6845 => conv_std_logic_vector(4914, 16),
6846 => conv_std_logic_vector(4940, 16),
6847 => conv_std_logic_vector(4966, 16),
6848 => conv_std_logic_vector(4992, 16),
6849 => conv_std_logic_vector(5018, 16),
6850 => conv_std_logic_vector(5044, 16),
6851 => conv_std_logic_vector(5070, 16),
6852 => conv_std_logic_vector(5096, 16),
6853 => conv_std_logic_vector(5122, 16),
6854 => conv_std_logic_vector(5148, 16),
6855 => conv_std_logic_vector(5174, 16),
6856 => conv_std_logic_vector(5200, 16),
6857 => conv_std_logic_vector(5226, 16),
6858 => conv_std_logic_vector(5252, 16),
6859 => conv_std_logic_vector(5278, 16),
6860 => conv_std_logic_vector(5304, 16),
6861 => conv_std_logic_vector(5330, 16),
6862 => conv_std_logic_vector(5356, 16),
6863 => conv_std_logic_vector(5382, 16),
6864 => conv_std_logic_vector(5408, 16),
6865 => conv_std_logic_vector(5434, 16),
6866 => conv_std_logic_vector(5460, 16),
6867 => conv_std_logic_vector(5486, 16),
6868 => conv_std_logic_vector(5512, 16),
6869 => conv_std_logic_vector(5538, 16),
6870 => conv_std_logic_vector(5564, 16),
6871 => conv_std_logic_vector(5590, 16),
6872 => conv_std_logic_vector(5616, 16),
6873 => conv_std_logic_vector(5642, 16),
6874 => conv_std_logic_vector(5668, 16),
6875 => conv_std_logic_vector(5694, 16),
6876 => conv_std_logic_vector(5720, 16),
6877 => conv_std_logic_vector(5746, 16),
6878 => conv_std_logic_vector(5772, 16),
6879 => conv_std_logic_vector(5798, 16),
6880 => conv_std_logic_vector(5824, 16),
6881 => conv_std_logic_vector(5850, 16),
6882 => conv_std_logic_vector(5876, 16),
6883 => conv_std_logic_vector(5902, 16),
6884 => conv_std_logic_vector(5928, 16),
6885 => conv_std_logic_vector(5954, 16),
6886 => conv_std_logic_vector(5980, 16),
6887 => conv_std_logic_vector(6006, 16),
6888 => conv_std_logic_vector(6032, 16),
6889 => conv_std_logic_vector(6058, 16),
6890 => conv_std_logic_vector(6084, 16),
6891 => conv_std_logic_vector(6110, 16),
6892 => conv_std_logic_vector(6136, 16),
6893 => conv_std_logic_vector(6162, 16),
6894 => conv_std_logic_vector(6188, 16),
6895 => conv_std_logic_vector(6214, 16),
6896 => conv_std_logic_vector(6240, 16),
6897 => conv_std_logic_vector(6266, 16),
6898 => conv_std_logic_vector(6292, 16),
6899 => conv_std_logic_vector(6318, 16),
6900 => conv_std_logic_vector(6344, 16),
6901 => conv_std_logic_vector(6370, 16),
6902 => conv_std_logic_vector(6396, 16),
6903 => conv_std_logic_vector(6422, 16),
6904 => conv_std_logic_vector(6448, 16),
6905 => conv_std_logic_vector(6474, 16),
6906 => conv_std_logic_vector(6500, 16),
6907 => conv_std_logic_vector(6526, 16),
6908 => conv_std_logic_vector(6552, 16),
6909 => conv_std_logic_vector(6578, 16),
6910 => conv_std_logic_vector(6604, 16),
6911 => conv_std_logic_vector(6630, 16),
6912 => conv_std_logic_vector(0, 16),
6913 => conv_std_logic_vector(27, 16),
6914 => conv_std_logic_vector(54, 16),
6915 => conv_std_logic_vector(81, 16),
6916 => conv_std_logic_vector(108, 16),
6917 => conv_std_logic_vector(135, 16),
6918 => conv_std_logic_vector(162, 16),
6919 => conv_std_logic_vector(189, 16),
6920 => conv_std_logic_vector(216, 16),
6921 => conv_std_logic_vector(243, 16),
6922 => conv_std_logic_vector(270, 16),
6923 => conv_std_logic_vector(297, 16),
6924 => conv_std_logic_vector(324, 16),
6925 => conv_std_logic_vector(351, 16),
6926 => conv_std_logic_vector(378, 16),
6927 => conv_std_logic_vector(405, 16),
6928 => conv_std_logic_vector(432, 16),
6929 => conv_std_logic_vector(459, 16),
6930 => conv_std_logic_vector(486, 16),
6931 => conv_std_logic_vector(513, 16),
6932 => conv_std_logic_vector(540, 16),
6933 => conv_std_logic_vector(567, 16),
6934 => conv_std_logic_vector(594, 16),
6935 => conv_std_logic_vector(621, 16),
6936 => conv_std_logic_vector(648, 16),
6937 => conv_std_logic_vector(675, 16),
6938 => conv_std_logic_vector(702, 16),
6939 => conv_std_logic_vector(729, 16),
6940 => conv_std_logic_vector(756, 16),
6941 => conv_std_logic_vector(783, 16),
6942 => conv_std_logic_vector(810, 16),
6943 => conv_std_logic_vector(837, 16),
6944 => conv_std_logic_vector(864, 16),
6945 => conv_std_logic_vector(891, 16),
6946 => conv_std_logic_vector(918, 16),
6947 => conv_std_logic_vector(945, 16),
6948 => conv_std_logic_vector(972, 16),
6949 => conv_std_logic_vector(999, 16),
6950 => conv_std_logic_vector(1026, 16),
6951 => conv_std_logic_vector(1053, 16),
6952 => conv_std_logic_vector(1080, 16),
6953 => conv_std_logic_vector(1107, 16),
6954 => conv_std_logic_vector(1134, 16),
6955 => conv_std_logic_vector(1161, 16),
6956 => conv_std_logic_vector(1188, 16),
6957 => conv_std_logic_vector(1215, 16),
6958 => conv_std_logic_vector(1242, 16),
6959 => conv_std_logic_vector(1269, 16),
6960 => conv_std_logic_vector(1296, 16),
6961 => conv_std_logic_vector(1323, 16),
6962 => conv_std_logic_vector(1350, 16),
6963 => conv_std_logic_vector(1377, 16),
6964 => conv_std_logic_vector(1404, 16),
6965 => conv_std_logic_vector(1431, 16),
6966 => conv_std_logic_vector(1458, 16),
6967 => conv_std_logic_vector(1485, 16),
6968 => conv_std_logic_vector(1512, 16),
6969 => conv_std_logic_vector(1539, 16),
6970 => conv_std_logic_vector(1566, 16),
6971 => conv_std_logic_vector(1593, 16),
6972 => conv_std_logic_vector(1620, 16),
6973 => conv_std_logic_vector(1647, 16),
6974 => conv_std_logic_vector(1674, 16),
6975 => conv_std_logic_vector(1701, 16),
6976 => conv_std_logic_vector(1728, 16),
6977 => conv_std_logic_vector(1755, 16),
6978 => conv_std_logic_vector(1782, 16),
6979 => conv_std_logic_vector(1809, 16),
6980 => conv_std_logic_vector(1836, 16),
6981 => conv_std_logic_vector(1863, 16),
6982 => conv_std_logic_vector(1890, 16),
6983 => conv_std_logic_vector(1917, 16),
6984 => conv_std_logic_vector(1944, 16),
6985 => conv_std_logic_vector(1971, 16),
6986 => conv_std_logic_vector(1998, 16),
6987 => conv_std_logic_vector(2025, 16),
6988 => conv_std_logic_vector(2052, 16),
6989 => conv_std_logic_vector(2079, 16),
6990 => conv_std_logic_vector(2106, 16),
6991 => conv_std_logic_vector(2133, 16),
6992 => conv_std_logic_vector(2160, 16),
6993 => conv_std_logic_vector(2187, 16),
6994 => conv_std_logic_vector(2214, 16),
6995 => conv_std_logic_vector(2241, 16),
6996 => conv_std_logic_vector(2268, 16),
6997 => conv_std_logic_vector(2295, 16),
6998 => conv_std_logic_vector(2322, 16),
6999 => conv_std_logic_vector(2349, 16),
7000 => conv_std_logic_vector(2376, 16),
7001 => conv_std_logic_vector(2403, 16),
7002 => conv_std_logic_vector(2430, 16),
7003 => conv_std_logic_vector(2457, 16),
7004 => conv_std_logic_vector(2484, 16),
7005 => conv_std_logic_vector(2511, 16),
7006 => conv_std_logic_vector(2538, 16),
7007 => conv_std_logic_vector(2565, 16),
7008 => conv_std_logic_vector(2592, 16),
7009 => conv_std_logic_vector(2619, 16),
7010 => conv_std_logic_vector(2646, 16),
7011 => conv_std_logic_vector(2673, 16),
7012 => conv_std_logic_vector(2700, 16),
7013 => conv_std_logic_vector(2727, 16),
7014 => conv_std_logic_vector(2754, 16),
7015 => conv_std_logic_vector(2781, 16),
7016 => conv_std_logic_vector(2808, 16),
7017 => conv_std_logic_vector(2835, 16),
7018 => conv_std_logic_vector(2862, 16),
7019 => conv_std_logic_vector(2889, 16),
7020 => conv_std_logic_vector(2916, 16),
7021 => conv_std_logic_vector(2943, 16),
7022 => conv_std_logic_vector(2970, 16),
7023 => conv_std_logic_vector(2997, 16),
7024 => conv_std_logic_vector(3024, 16),
7025 => conv_std_logic_vector(3051, 16),
7026 => conv_std_logic_vector(3078, 16),
7027 => conv_std_logic_vector(3105, 16),
7028 => conv_std_logic_vector(3132, 16),
7029 => conv_std_logic_vector(3159, 16),
7030 => conv_std_logic_vector(3186, 16),
7031 => conv_std_logic_vector(3213, 16),
7032 => conv_std_logic_vector(3240, 16),
7033 => conv_std_logic_vector(3267, 16),
7034 => conv_std_logic_vector(3294, 16),
7035 => conv_std_logic_vector(3321, 16),
7036 => conv_std_logic_vector(3348, 16),
7037 => conv_std_logic_vector(3375, 16),
7038 => conv_std_logic_vector(3402, 16),
7039 => conv_std_logic_vector(3429, 16),
7040 => conv_std_logic_vector(3456, 16),
7041 => conv_std_logic_vector(3483, 16),
7042 => conv_std_logic_vector(3510, 16),
7043 => conv_std_logic_vector(3537, 16),
7044 => conv_std_logic_vector(3564, 16),
7045 => conv_std_logic_vector(3591, 16),
7046 => conv_std_logic_vector(3618, 16),
7047 => conv_std_logic_vector(3645, 16),
7048 => conv_std_logic_vector(3672, 16),
7049 => conv_std_logic_vector(3699, 16),
7050 => conv_std_logic_vector(3726, 16),
7051 => conv_std_logic_vector(3753, 16),
7052 => conv_std_logic_vector(3780, 16),
7053 => conv_std_logic_vector(3807, 16),
7054 => conv_std_logic_vector(3834, 16),
7055 => conv_std_logic_vector(3861, 16),
7056 => conv_std_logic_vector(3888, 16),
7057 => conv_std_logic_vector(3915, 16),
7058 => conv_std_logic_vector(3942, 16),
7059 => conv_std_logic_vector(3969, 16),
7060 => conv_std_logic_vector(3996, 16),
7061 => conv_std_logic_vector(4023, 16),
7062 => conv_std_logic_vector(4050, 16),
7063 => conv_std_logic_vector(4077, 16),
7064 => conv_std_logic_vector(4104, 16),
7065 => conv_std_logic_vector(4131, 16),
7066 => conv_std_logic_vector(4158, 16),
7067 => conv_std_logic_vector(4185, 16),
7068 => conv_std_logic_vector(4212, 16),
7069 => conv_std_logic_vector(4239, 16),
7070 => conv_std_logic_vector(4266, 16),
7071 => conv_std_logic_vector(4293, 16),
7072 => conv_std_logic_vector(4320, 16),
7073 => conv_std_logic_vector(4347, 16),
7074 => conv_std_logic_vector(4374, 16),
7075 => conv_std_logic_vector(4401, 16),
7076 => conv_std_logic_vector(4428, 16),
7077 => conv_std_logic_vector(4455, 16),
7078 => conv_std_logic_vector(4482, 16),
7079 => conv_std_logic_vector(4509, 16),
7080 => conv_std_logic_vector(4536, 16),
7081 => conv_std_logic_vector(4563, 16),
7082 => conv_std_logic_vector(4590, 16),
7083 => conv_std_logic_vector(4617, 16),
7084 => conv_std_logic_vector(4644, 16),
7085 => conv_std_logic_vector(4671, 16),
7086 => conv_std_logic_vector(4698, 16),
7087 => conv_std_logic_vector(4725, 16),
7088 => conv_std_logic_vector(4752, 16),
7089 => conv_std_logic_vector(4779, 16),
7090 => conv_std_logic_vector(4806, 16),
7091 => conv_std_logic_vector(4833, 16),
7092 => conv_std_logic_vector(4860, 16),
7093 => conv_std_logic_vector(4887, 16),
7094 => conv_std_logic_vector(4914, 16),
7095 => conv_std_logic_vector(4941, 16),
7096 => conv_std_logic_vector(4968, 16),
7097 => conv_std_logic_vector(4995, 16),
7098 => conv_std_logic_vector(5022, 16),
7099 => conv_std_logic_vector(5049, 16),
7100 => conv_std_logic_vector(5076, 16),
7101 => conv_std_logic_vector(5103, 16),
7102 => conv_std_logic_vector(5130, 16),
7103 => conv_std_logic_vector(5157, 16),
7104 => conv_std_logic_vector(5184, 16),
7105 => conv_std_logic_vector(5211, 16),
7106 => conv_std_logic_vector(5238, 16),
7107 => conv_std_logic_vector(5265, 16),
7108 => conv_std_logic_vector(5292, 16),
7109 => conv_std_logic_vector(5319, 16),
7110 => conv_std_logic_vector(5346, 16),
7111 => conv_std_logic_vector(5373, 16),
7112 => conv_std_logic_vector(5400, 16),
7113 => conv_std_logic_vector(5427, 16),
7114 => conv_std_logic_vector(5454, 16),
7115 => conv_std_logic_vector(5481, 16),
7116 => conv_std_logic_vector(5508, 16),
7117 => conv_std_logic_vector(5535, 16),
7118 => conv_std_logic_vector(5562, 16),
7119 => conv_std_logic_vector(5589, 16),
7120 => conv_std_logic_vector(5616, 16),
7121 => conv_std_logic_vector(5643, 16),
7122 => conv_std_logic_vector(5670, 16),
7123 => conv_std_logic_vector(5697, 16),
7124 => conv_std_logic_vector(5724, 16),
7125 => conv_std_logic_vector(5751, 16),
7126 => conv_std_logic_vector(5778, 16),
7127 => conv_std_logic_vector(5805, 16),
7128 => conv_std_logic_vector(5832, 16),
7129 => conv_std_logic_vector(5859, 16),
7130 => conv_std_logic_vector(5886, 16),
7131 => conv_std_logic_vector(5913, 16),
7132 => conv_std_logic_vector(5940, 16),
7133 => conv_std_logic_vector(5967, 16),
7134 => conv_std_logic_vector(5994, 16),
7135 => conv_std_logic_vector(6021, 16),
7136 => conv_std_logic_vector(6048, 16),
7137 => conv_std_logic_vector(6075, 16),
7138 => conv_std_logic_vector(6102, 16),
7139 => conv_std_logic_vector(6129, 16),
7140 => conv_std_logic_vector(6156, 16),
7141 => conv_std_logic_vector(6183, 16),
7142 => conv_std_logic_vector(6210, 16),
7143 => conv_std_logic_vector(6237, 16),
7144 => conv_std_logic_vector(6264, 16),
7145 => conv_std_logic_vector(6291, 16),
7146 => conv_std_logic_vector(6318, 16),
7147 => conv_std_logic_vector(6345, 16),
7148 => conv_std_logic_vector(6372, 16),
7149 => conv_std_logic_vector(6399, 16),
7150 => conv_std_logic_vector(6426, 16),
7151 => conv_std_logic_vector(6453, 16),
7152 => conv_std_logic_vector(6480, 16),
7153 => conv_std_logic_vector(6507, 16),
7154 => conv_std_logic_vector(6534, 16),
7155 => conv_std_logic_vector(6561, 16),
7156 => conv_std_logic_vector(6588, 16),
7157 => conv_std_logic_vector(6615, 16),
7158 => conv_std_logic_vector(6642, 16),
7159 => conv_std_logic_vector(6669, 16),
7160 => conv_std_logic_vector(6696, 16),
7161 => conv_std_logic_vector(6723, 16),
7162 => conv_std_logic_vector(6750, 16),
7163 => conv_std_logic_vector(6777, 16),
7164 => conv_std_logic_vector(6804, 16),
7165 => conv_std_logic_vector(6831, 16),
7166 => conv_std_logic_vector(6858, 16),
7167 => conv_std_logic_vector(6885, 16),
7168 => conv_std_logic_vector(0, 16),
7169 => conv_std_logic_vector(28, 16),
7170 => conv_std_logic_vector(56, 16),
7171 => conv_std_logic_vector(84, 16),
7172 => conv_std_logic_vector(112, 16),
7173 => conv_std_logic_vector(140, 16),
7174 => conv_std_logic_vector(168, 16),
7175 => conv_std_logic_vector(196, 16),
7176 => conv_std_logic_vector(224, 16),
7177 => conv_std_logic_vector(252, 16),
7178 => conv_std_logic_vector(280, 16),
7179 => conv_std_logic_vector(308, 16),
7180 => conv_std_logic_vector(336, 16),
7181 => conv_std_logic_vector(364, 16),
7182 => conv_std_logic_vector(392, 16),
7183 => conv_std_logic_vector(420, 16),
7184 => conv_std_logic_vector(448, 16),
7185 => conv_std_logic_vector(476, 16),
7186 => conv_std_logic_vector(504, 16),
7187 => conv_std_logic_vector(532, 16),
7188 => conv_std_logic_vector(560, 16),
7189 => conv_std_logic_vector(588, 16),
7190 => conv_std_logic_vector(616, 16),
7191 => conv_std_logic_vector(644, 16),
7192 => conv_std_logic_vector(672, 16),
7193 => conv_std_logic_vector(700, 16),
7194 => conv_std_logic_vector(728, 16),
7195 => conv_std_logic_vector(756, 16),
7196 => conv_std_logic_vector(784, 16),
7197 => conv_std_logic_vector(812, 16),
7198 => conv_std_logic_vector(840, 16),
7199 => conv_std_logic_vector(868, 16),
7200 => conv_std_logic_vector(896, 16),
7201 => conv_std_logic_vector(924, 16),
7202 => conv_std_logic_vector(952, 16),
7203 => conv_std_logic_vector(980, 16),
7204 => conv_std_logic_vector(1008, 16),
7205 => conv_std_logic_vector(1036, 16),
7206 => conv_std_logic_vector(1064, 16),
7207 => conv_std_logic_vector(1092, 16),
7208 => conv_std_logic_vector(1120, 16),
7209 => conv_std_logic_vector(1148, 16),
7210 => conv_std_logic_vector(1176, 16),
7211 => conv_std_logic_vector(1204, 16),
7212 => conv_std_logic_vector(1232, 16),
7213 => conv_std_logic_vector(1260, 16),
7214 => conv_std_logic_vector(1288, 16),
7215 => conv_std_logic_vector(1316, 16),
7216 => conv_std_logic_vector(1344, 16),
7217 => conv_std_logic_vector(1372, 16),
7218 => conv_std_logic_vector(1400, 16),
7219 => conv_std_logic_vector(1428, 16),
7220 => conv_std_logic_vector(1456, 16),
7221 => conv_std_logic_vector(1484, 16),
7222 => conv_std_logic_vector(1512, 16),
7223 => conv_std_logic_vector(1540, 16),
7224 => conv_std_logic_vector(1568, 16),
7225 => conv_std_logic_vector(1596, 16),
7226 => conv_std_logic_vector(1624, 16),
7227 => conv_std_logic_vector(1652, 16),
7228 => conv_std_logic_vector(1680, 16),
7229 => conv_std_logic_vector(1708, 16),
7230 => conv_std_logic_vector(1736, 16),
7231 => conv_std_logic_vector(1764, 16),
7232 => conv_std_logic_vector(1792, 16),
7233 => conv_std_logic_vector(1820, 16),
7234 => conv_std_logic_vector(1848, 16),
7235 => conv_std_logic_vector(1876, 16),
7236 => conv_std_logic_vector(1904, 16),
7237 => conv_std_logic_vector(1932, 16),
7238 => conv_std_logic_vector(1960, 16),
7239 => conv_std_logic_vector(1988, 16),
7240 => conv_std_logic_vector(2016, 16),
7241 => conv_std_logic_vector(2044, 16),
7242 => conv_std_logic_vector(2072, 16),
7243 => conv_std_logic_vector(2100, 16),
7244 => conv_std_logic_vector(2128, 16),
7245 => conv_std_logic_vector(2156, 16),
7246 => conv_std_logic_vector(2184, 16),
7247 => conv_std_logic_vector(2212, 16),
7248 => conv_std_logic_vector(2240, 16),
7249 => conv_std_logic_vector(2268, 16),
7250 => conv_std_logic_vector(2296, 16),
7251 => conv_std_logic_vector(2324, 16),
7252 => conv_std_logic_vector(2352, 16),
7253 => conv_std_logic_vector(2380, 16),
7254 => conv_std_logic_vector(2408, 16),
7255 => conv_std_logic_vector(2436, 16),
7256 => conv_std_logic_vector(2464, 16),
7257 => conv_std_logic_vector(2492, 16),
7258 => conv_std_logic_vector(2520, 16),
7259 => conv_std_logic_vector(2548, 16),
7260 => conv_std_logic_vector(2576, 16),
7261 => conv_std_logic_vector(2604, 16),
7262 => conv_std_logic_vector(2632, 16),
7263 => conv_std_logic_vector(2660, 16),
7264 => conv_std_logic_vector(2688, 16),
7265 => conv_std_logic_vector(2716, 16),
7266 => conv_std_logic_vector(2744, 16),
7267 => conv_std_logic_vector(2772, 16),
7268 => conv_std_logic_vector(2800, 16),
7269 => conv_std_logic_vector(2828, 16),
7270 => conv_std_logic_vector(2856, 16),
7271 => conv_std_logic_vector(2884, 16),
7272 => conv_std_logic_vector(2912, 16),
7273 => conv_std_logic_vector(2940, 16),
7274 => conv_std_logic_vector(2968, 16),
7275 => conv_std_logic_vector(2996, 16),
7276 => conv_std_logic_vector(3024, 16),
7277 => conv_std_logic_vector(3052, 16),
7278 => conv_std_logic_vector(3080, 16),
7279 => conv_std_logic_vector(3108, 16),
7280 => conv_std_logic_vector(3136, 16),
7281 => conv_std_logic_vector(3164, 16),
7282 => conv_std_logic_vector(3192, 16),
7283 => conv_std_logic_vector(3220, 16),
7284 => conv_std_logic_vector(3248, 16),
7285 => conv_std_logic_vector(3276, 16),
7286 => conv_std_logic_vector(3304, 16),
7287 => conv_std_logic_vector(3332, 16),
7288 => conv_std_logic_vector(3360, 16),
7289 => conv_std_logic_vector(3388, 16),
7290 => conv_std_logic_vector(3416, 16),
7291 => conv_std_logic_vector(3444, 16),
7292 => conv_std_logic_vector(3472, 16),
7293 => conv_std_logic_vector(3500, 16),
7294 => conv_std_logic_vector(3528, 16),
7295 => conv_std_logic_vector(3556, 16),
7296 => conv_std_logic_vector(3584, 16),
7297 => conv_std_logic_vector(3612, 16),
7298 => conv_std_logic_vector(3640, 16),
7299 => conv_std_logic_vector(3668, 16),
7300 => conv_std_logic_vector(3696, 16),
7301 => conv_std_logic_vector(3724, 16),
7302 => conv_std_logic_vector(3752, 16),
7303 => conv_std_logic_vector(3780, 16),
7304 => conv_std_logic_vector(3808, 16),
7305 => conv_std_logic_vector(3836, 16),
7306 => conv_std_logic_vector(3864, 16),
7307 => conv_std_logic_vector(3892, 16),
7308 => conv_std_logic_vector(3920, 16),
7309 => conv_std_logic_vector(3948, 16),
7310 => conv_std_logic_vector(3976, 16),
7311 => conv_std_logic_vector(4004, 16),
7312 => conv_std_logic_vector(4032, 16),
7313 => conv_std_logic_vector(4060, 16),
7314 => conv_std_logic_vector(4088, 16),
7315 => conv_std_logic_vector(4116, 16),
7316 => conv_std_logic_vector(4144, 16),
7317 => conv_std_logic_vector(4172, 16),
7318 => conv_std_logic_vector(4200, 16),
7319 => conv_std_logic_vector(4228, 16),
7320 => conv_std_logic_vector(4256, 16),
7321 => conv_std_logic_vector(4284, 16),
7322 => conv_std_logic_vector(4312, 16),
7323 => conv_std_logic_vector(4340, 16),
7324 => conv_std_logic_vector(4368, 16),
7325 => conv_std_logic_vector(4396, 16),
7326 => conv_std_logic_vector(4424, 16),
7327 => conv_std_logic_vector(4452, 16),
7328 => conv_std_logic_vector(4480, 16),
7329 => conv_std_logic_vector(4508, 16),
7330 => conv_std_logic_vector(4536, 16),
7331 => conv_std_logic_vector(4564, 16),
7332 => conv_std_logic_vector(4592, 16),
7333 => conv_std_logic_vector(4620, 16),
7334 => conv_std_logic_vector(4648, 16),
7335 => conv_std_logic_vector(4676, 16),
7336 => conv_std_logic_vector(4704, 16),
7337 => conv_std_logic_vector(4732, 16),
7338 => conv_std_logic_vector(4760, 16),
7339 => conv_std_logic_vector(4788, 16),
7340 => conv_std_logic_vector(4816, 16),
7341 => conv_std_logic_vector(4844, 16),
7342 => conv_std_logic_vector(4872, 16),
7343 => conv_std_logic_vector(4900, 16),
7344 => conv_std_logic_vector(4928, 16),
7345 => conv_std_logic_vector(4956, 16),
7346 => conv_std_logic_vector(4984, 16),
7347 => conv_std_logic_vector(5012, 16),
7348 => conv_std_logic_vector(5040, 16),
7349 => conv_std_logic_vector(5068, 16),
7350 => conv_std_logic_vector(5096, 16),
7351 => conv_std_logic_vector(5124, 16),
7352 => conv_std_logic_vector(5152, 16),
7353 => conv_std_logic_vector(5180, 16),
7354 => conv_std_logic_vector(5208, 16),
7355 => conv_std_logic_vector(5236, 16),
7356 => conv_std_logic_vector(5264, 16),
7357 => conv_std_logic_vector(5292, 16),
7358 => conv_std_logic_vector(5320, 16),
7359 => conv_std_logic_vector(5348, 16),
7360 => conv_std_logic_vector(5376, 16),
7361 => conv_std_logic_vector(5404, 16),
7362 => conv_std_logic_vector(5432, 16),
7363 => conv_std_logic_vector(5460, 16),
7364 => conv_std_logic_vector(5488, 16),
7365 => conv_std_logic_vector(5516, 16),
7366 => conv_std_logic_vector(5544, 16),
7367 => conv_std_logic_vector(5572, 16),
7368 => conv_std_logic_vector(5600, 16),
7369 => conv_std_logic_vector(5628, 16),
7370 => conv_std_logic_vector(5656, 16),
7371 => conv_std_logic_vector(5684, 16),
7372 => conv_std_logic_vector(5712, 16),
7373 => conv_std_logic_vector(5740, 16),
7374 => conv_std_logic_vector(5768, 16),
7375 => conv_std_logic_vector(5796, 16),
7376 => conv_std_logic_vector(5824, 16),
7377 => conv_std_logic_vector(5852, 16),
7378 => conv_std_logic_vector(5880, 16),
7379 => conv_std_logic_vector(5908, 16),
7380 => conv_std_logic_vector(5936, 16),
7381 => conv_std_logic_vector(5964, 16),
7382 => conv_std_logic_vector(5992, 16),
7383 => conv_std_logic_vector(6020, 16),
7384 => conv_std_logic_vector(6048, 16),
7385 => conv_std_logic_vector(6076, 16),
7386 => conv_std_logic_vector(6104, 16),
7387 => conv_std_logic_vector(6132, 16),
7388 => conv_std_logic_vector(6160, 16),
7389 => conv_std_logic_vector(6188, 16),
7390 => conv_std_logic_vector(6216, 16),
7391 => conv_std_logic_vector(6244, 16),
7392 => conv_std_logic_vector(6272, 16),
7393 => conv_std_logic_vector(6300, 16),
7394 => conv_std_logic_vector(6328, 16),
7395 => conv_std_logic_vector(6356, 16),
7396 => conv_std_logic_vector(6384, 16),
7397 => conv_std_logic_vector(6412, 16),
7398 => conv_std_logic_vector(6440, 16),
7399 => conv_std_logic_vector(6468, 16),
7400 => conv_std_logic_vector(6496, 16),
7401 => conv_std_logic_vector(6524, 16),
7402 => conv_std_logic_vector(6552, 16),
7403 => conv_std_logic_vector(6580, 16),
7404 => conv_std_logic_vector(6608, 16),
7405 => conv_std_logic_vector(6636, 16),
7406 => conv_std_logic_vector(6664, 16),
7407 => conv_std_logic_vector(6692, 16),
7408 => conv_std_logic_vector(6720, 16),
7409 => conv_std_logic_vector(6748, 16),
7410 => conv_std_logic_vector(6776, 16),
7411 => conv_std_logic_vector(6804, 16),
7412 => conv_std_logic_vector(6832, 16),
7413 => conv_std_logic_vector(6860, 16),
7414 => conv_std_logic_vector(6888, 16),
7415 => conv_std_logic_vector(6916, 16),
7416 => conv_std_logic_vector(6944, 16),
7417 => conv_std_logic_vector(6972, 16),
7418 => conv_std_logic_vector(7000, 16),
7419 => conv_std_logic_vector(7028, 16),
7420 => conv_std_logic_vector(7056, 16),
7421 => conv_std_logic_vector(7084, 16),
7422 => conv_std_logic_vector(7112, 16),
7423 => conv_std_logic_vector(7140, 16),
7424 => conv_std_logic_vector(0, 16),
7425 => conv_std_logic_vector(29, 16),
7426 => conv_std_logic_vector(58, 16),
7427 => conv_std_logic_vector(87, 16),
7428 => conv_std_logic_vector(116, 16),
7429 => conv_std_logic_vector(145, 16),
7430 => conv_std_logic_vector(174, 16),
7431 => conv_std_logic_vector(203, 16),
7432 => conv_std_logic_vector(232, 16),
7433 => conv_std_logic_vector(261, 16),
7434 => conv_std_logic_vector(290, 16),
7435 => conv_std_logic_vector(319, 16),
7436 => conv_std_logic_vector(348, 16),
7437 => conv_std_logic_vector(377, 16),
7438 => conv_std_logic_vector(406, 16),
7439 => conv_std_logic_vector(435, 16),
7440 => conv_std_logic_vector(464, 16),
7441 => conv_std_logic_vector(493, 16),
7442 => conv_std_logic_vector(522, 16),
7443 => conv_std_logic_vector(551, 16),
7444 => conv_std_logic_vector(580, 16),
7445 => conv_std_logic_vector(609, 16),
7446 => conv_std_logic_vector(638, 16),
7447 => conv_std_logic_vector(667, 16),
7448 => conv_std_logic_vector(696, 16),
7449 => conv_std_logic_vector(725, 16),
7450 => conv_std_logic_vector(754, 16),
7451 => conv_std_logic_vector(783, 16),
7452 => conv_std_logic_vector(812, 16),
7453 => conv_std_logic_vector(841, 16),
7454 => conv_std_logic_vector(870, 16),
7455 => conv_std_logic_vector(899, 16),
7456 => conv_std_logic_vector(928, 16),
7457 => conv_std_logic_vector(957, 16),
7458 => conv_std_logic_vector(986, 16),
7459 => conv_std_logic_vector(1015, 16),
7460 => conv_std_logic_vector(1044, 16),
7461 => conv_std_logic_vector(1073, 16),
7462 => conv_std_logic_vector(1102, 16),
7463 => conv_std_logic_vector(1131, 16),
7464 => conv_std_logic_vector(1160, 16),
7465 => conv_std_logic_vector(1189, 16),
7466 => conv_std_logic_vector(1218, 16),
7467 => conv_std_logic_vector(1247, 16),
7468 => conv_std_logic_vector(1276, 16),
7469 => conv_std_logic_vector(1305, 16),
7470 => conv_std_logic_vector(1334, 16),
7471 => conv_std_logic_vector(1363, 16),
7472 => conv_std_logic_vector(1392, 16),
7473 => conv_std_logic_vector(1421, 16),
7474 => conv_std_logic_vector(1450, 16),
7475 => conv_std_logic_vector(1479, 16),
7476 => conv_std_logic_vector(1508, 16),
7477 => conv_std_logic_vector(1537, 16),
7478 => conv_std_logic_vector(1566, 16),
7479 => conv_std_logic_vector(1595, 16),
7480 => conv_std_logic_vector(1624, 16),
7481 => conv_std_logic_vector(1653, 16),
7482 => conv_std_logic_vector(1682, 16),
7483 => conv_std_logic_vector(1711, 16),
7484 => conv_std_logic_vector(1740, 16),
7485 => conv_std_logic_vector(1769, 16),
7486 => conv_std_logic_vector(1798, 16),
7487 => conv_std_logic_vector(1827, 16),
7488 => conv_std_logic_vector(1856, 16),
7489 => conv_std_logic_vector(1885, 16),
7490 => conv_std_logic_vector(1914, 16),
7491 => conv_std_logic_vector(1943, 16),
7492 => conv_std_logic_vector(1972, 16),
7493 => conv_std_logic_vector(2001, 16),
7494 => conv_std_logic_vector(2030, 16),
7495 => conv_std_logic_vector(2059, 16),
7496 => conv_std_logic_vector(2088, 16),
7497 => conv_std_logic_vector(2117, 16),
7498 => conv_std_logic_vector(2146, 16),
7499 => conv_std_logic_vector(2175, 16),
7500 => conv_std_logic_vector(2204, 16),
7501 => conv_std_logic_vector(2233, 16),
7502 => conv_std_logic_vector(2262, 16),
7503 => conv_std_logic_vector(2291, 16),
7504 => conv_std_logic_vector(2320, 16),
7505 => conv_std_logic_vector(2349, 16),
7506 => conv_std_logic_vector(2378, 16),
7507 => conv_std_logic_vector(2407, 16),
7508 => conv_std_logic_vector(2436, 16),
7509 => conv_std_logic_vector(2465, 16),
7510 => conv_std_logic_vector(2494, 16),
7511 => conv_std_logic_vector(2523, 16),
7512 => conv_std_logic_vector(2552, 16),
7513 => conv_std_logic_vector(2581, 16),
7514 => conv_std_logic_vector(2610, 16),
7515 => conv_std_logic_vector(2639, 16),
7516 => conv_std_logic_vector(2668, 16),
7517 => conv_std_logic_vector(2697, 16),
7518 => conv_std_logic_vector(2726, 16),
7519 => conv_std_logic_vector(2755, 16),
7520 => conv_std_logic_vector(2784, 16),
7521 => conv_std_logic_vector(2813, 16),
7522 => conv_std_logic_vector(2842, 16),
7523 => conv_std_logic_vector(2871, 16),
7524 => conv_std_logic_vector(2900, 16),
7525 => conv_std_logic_vector(2929, 16),
7526 => conv_std_logic_vector(2958, 16),
7527 => conv_std_logic_vector(2987, 16),
7528 => conv_std_logic_vector(3016, 16),
7529 => conv_std_logic_vector(3045, 16),
7530 => conv_std_logic_vector(3074, 16),
7531 => conv_std_logic_vector(3103, 16),
7532 => conv_std_logic_vector(3132, 16),
7533 => conv_std_logic_vector(3161, 16),
7534 => conv_std_logic_vector(3190, 16),
7535 => conv_std_logic_vector(3219, 16),
7536 => conv_std_logic_vector(3248, 16),
7537 => conv_std_logic_vector(3277, 16),
7538 => conv_std_logic_vector(3306, 16),
7539 => conv_std_logic_vector(3335, 16),
7540 => conv_std_logic_vector(3364, 16),
7541 => conv_std_logic_vector(3393, 16),
7542 => conv_std_logic_vector(3422, 16),
7543 => conv_std_logic_vector(3451, 16),
7544 => conv_std_logic_vector(3480, 16),
7545 => conv_std_logic_vector(3509, 16),
7546 => conv_std_logic_vector(3538, 16),
7547 => conv_std_logic_vector(3567, 16),
7548 => conv_std_logic_vector(3596, 16),
7549 => conv_std_logic_vector(3625, 16),
7550 => conv_std_logic_vector(3654, 16),
7551 => conv_std_logic_vector(3683, 16),
7552 => conv_std_logic_vector(3712, 16),
7553 => conv_std_logic_vector(3741, 16),
7554 => conv_std_logic_vector(3770, 16),
7555 => conv_std_logic_vector(3799, 16),
7556 => conv_std_logic_vector(3828, 16),
7557 => conv_std_logic_vector(3857, 16),
7558 => conv_std_logic_vector(3886, 16),
7559 => conv_std_logic_vector(3915, 16),
7560 => conv_std_logic_vector(3944, 16),
7561 => conv_std_logic_vector(3973, 16),
7562 => conv_std_logic_vector(4002, 16),
7563 => conv_std_logic_vector(4031, 16),
7564 => conv_std_logic_vector(4060, 16),
7565 => conv_std_logic_vector(4089, 16),
7566 => conv_std_logic_vector(4118, 16),
7567 => conv_std_logic_vector(4147, 16),
7568 => conv_std_logic_vector(4176, 16),
7569 => conv_std_logic_vector(4205, 16),
7570 => conv_std_logic_vector(4234, 16),
7571 => conv_std_logic_vector(4263, 16),
7572 => conv_std_logic_vector(4292, 16),
7573 => conv_std_logic_vector(4321, 16),
7574 => conv_std_logic_vector(4350, 16),
7575 => conv_std_logic_vector(4379, 16),
7576 => conv_std_logic_vector(4408, 16),
7577 => conv_std_logic_vector(4437, 16),
7578 => conv_std_logic_vector(4466, 16),
7579 => conv_std_logic_vector(4495, 16),
7580 => conv_std_logic_vector(4524, 16),
7581 => conv_std_logic_vector(4553, 16),
7582 => conv_std_logic_vector(4582, 16),
7583 => conv_std_logic_vector(4611, 16),
7584 => conv_std_logic_vector(4640, 16),
7585 => conv_std_logic_vector(4669, 16),
7586 => conv_std_logic_vector(4698, 16),
7587 => conv_std_logic_vector(4727, 16),
7588 => conv_std_logic_vector(4756, 16),
7589 => conv_std_logic_vector(4785, 16),
7590 => conv_std_logic_vector(4814, 16),
7591 => conv_std_logic_vector(4843, 16),
7592 => conv_std_logic_vector(4872, 16),
7593 => conv_std_logic_vector(4901, 16),
7594 => conv_std_logic_vector(4930, 16),
7595 => conv_std_logic_vector(4959, 16),
7596 => conv_std_logic_vector(4988, 16),
7597 => conv_std_logic_vector(5017, 16),
7598 => conv_std_logic_vector(5046, 16),
7599 => conv_std_logic_vector(5075, 16),
7600 => conv_std_logic_vector(5104, 16),
7601 => conv_std_logic_vector(5133, 16),
7602 => conv_std_logic_vector(5162, 16),
7603 => conv_std_logic_vector(5191, 16),
7604 => conv_std_logic_vector(5220, 16),
7605 => conv_std_logic_vector(5249, 16),
7606 => conv_std_logic_vector(5278, 16),
7607 => conv_std_logic_vector(5307, 16),
7608 => conv_std_logic_vector(5336, 16),
7609 => conv_std_logic_vector(5365, 16),
7610 => conv_std_logic_vector(5394, 16),
7611 => conv_std_logic_vector(5423, 16),
7612 => conv_std_logic_vector(5452, 16),
7613 => conv_std_logic_vector(5481, 16),
7614 => conv_std_logic_vector(5510, 16),
7615 => conv_std_logic_vector(5539, 16),
7616 => conv_std_logic_vector(5568, 16),
7617 => conv_std_logic_vector(5597, 16),
7618 => conv_std_logic_vector(5626, 16),
7619 => conv_std_logic_vector(5655, 16),
7620 => conv_std_logic_vector(5684, 16),
7621 => conv_std_logic_vector(5713, 16),
7622 => conv_std_logic_vector(5742, 16),
7623 => conv_std_logic_vector(5771, 16),
7624 => conv_std_logic_vector(5800, 16),
7625 => conv_std_logic_vector(5829, 16),
7626 => conv_std_logic_vector(5858, 16),
7627 => conv_std_logic_vector(5887, 16),
7628 => conv_std_logic_vector(5916, 16),
7629 => conv_std_logic_vector(5945, 16),
7630 => conv_std_logic_vector(5974, 16),
7631 => conv_std_logic_vector(6003, 16),
7632 => conv_std_logic_vector(6032, 16),
7633 => conv_std_logic_vector(6061, 16),
7634 => conv_std_logic_vector(6090, 16),
7635 => conv_std_logic_vector(6119, 16),
7636 => conv_std_logic_vector(6148, 16),
7637 => conv_std_logic_vector(6177, 16),
7638 => conv_std_logic_vector(6206, 16),
7639 => conv_std_logic_vector(6235, 16),
7640 => conv_std_logic_vector(6264, 16),
7641 => conv_std_logic_vector(6293, 16),
7642 => conv_std_logic_vector(6322, 16),
7643 => conv_std_logic_vector(6351, 16),
7644 => conv_std_logic_vector(6380, 16),
7645 => conv_std_logic_vector(6409, 16),
7646 => conv_std_logic_vector(6438, 16),
7647 => conv_std_logic_vector(6467, 16),
7648 => conv_std_logic_vector(6496, 16),
7649 => conv_std_logic_vector(6525, 16),
7650 => conv_std_logic_vector(6554, 16),
7651 => conv_std_logic_vector(6583, 16),
7652 => conv_std_logic_vector(6612, 16),
7653 => conv_std_logic_vector(6641, 16),
7654 => conv_std_logic_vector(6670, 16),
7655 => conv_std_logic_vector(6699, 16),
7656 => conv_std_logic_vector(6728, 16),
7657 => conv_std_logic_vector(6757, 16),
7658 => conv_std_logic_vector(6786, 16),
7659 => conv_std_logic_vector(6815, 16),
7660 => conv_std_logic_vector(6844, 16),
7661 => conv_std_logic_vector(6873, 16),
7662 => conv_std_logic_vector(6902, 16),
7663 => conv_std_logic_vector(6931, 16),
7664 => conv_std_logic_vector(6960, 16),
7665 => conv_std_logic_vector(6989, 16),
7666 => conv_std_logic_vector(7018, 16),
7667 => conv_std_logic_vector(7047, 16),
7668 => conv_std_logic_vector(7076, 16),
7669 => conv_std_logic_vector(7105, 16),
7670 => conv_std_logic_vector(7134, 16),
7671 => conv_std_logic_vector(7163, 16),
7672 => conv_std_logic_vector(7192, 16),
7673 => conv_std_logic_vector(7221, 16),
7674 => conv_std_logic_vector(7250, 16),
7675 => conv_std_logic_vector(7279, 16),
7676 => conv_std_logic_vector(7308, 16),
7677 => conv_std_logic_vector(7337, 16),
7678 => conv_std_logic_vector(7366, 16),
7679 => conv_std_logic_vector(7395, 16),
7680 => conv_std_logic_vector(0, 16),
7681 => conv_std_logic_vector(30, 16),
7682 => conv_std_logic_vector(60, 16),
7683 => conv_std_logic_vector(90, 16),
7684 => conv_std_logic_vector(120, 16),
7685 => conv_std_logic_vector(150, 16),
7686 => conv_std_logic_vector(180, 16),
7687 => conv_std_logic_vector(210, 16),
7688 => conv_std_logic_vector(240, 16),
7689 => conv_std_logic_vector(270, 16),
7690 => conv_std_logic_vector(300, 16),
7691 => conv_std_logic_vector(330, 16),
7692 => conv_std_logic_vector(360, 16),
7693 => conv_std_logic_vector(390, 16),
7694 => conv_std_logic_vector(420, 16),
7695 => conv_std_logic_vector(450, 16),
7696 => conv_std_logic_vector(480, 16),
7697 => conv_std_logic_vector(510, 16),
7698 => conv_std_logic_vector(540, 16),
7699 => conv_std_logic_vector(570, 16),
7700 => conv_std_logic_vector(600, 16),
7701 => conv_std_logic_vector(630, 16),
7702 => conv_std_logic_vector(660, 16),
7703 => conv_std_logic_vector(690, 16),
7704 => conv_std_logic_vector(720, 16),
7705 => conv_std_logic_vector(750, 16),
7706 => conv_std_logic_vector(780, 16),
7707 => conv_std_logic_vector(810, 16),
7708 => conv_std_logic_vector(840, 16),
7709 => conv_std_logic_vector(870, 16),
7710 => conv_std_logic_vector(900, 16),
7711 => conv_std_logic_vector(930, 16),
7712 => conv_std_logic_vector(960, 16),
7713 => conv_std_logic_vector(990, 16),
7714 => conv_std_logic_vector(1020, 16),
7715 => conv_std_logic_vector(1050, 16),
7716 => conv_std_logic_vector(1080, 16),
7717 => conv_std_logic_vector(1110, 16),
7718 => conv_std_logic_vector(1140, 16),
7719 => conv_std_logic_vector(1170, 16),
7720 => conv_std_logic_vector(1200, 16),
7721 => conv_std_logic_vector(1230, 16),
7722 => conv_std_logic_vector(1260, 16),
7723 => conv_std_logic_vector(1290, 16),
7724 => conv_std_logic_vector(1320, 16),
7725 => conv_std_logic_vector(1350, 16),
7726 => conv_std_logic_vector(1380, 16),
7727 => conv_std_logic_vector(1410, 16),
7728 => conv_std_logic_vector(1440, 16),
7729 => conv_std_logic_vector(1470, 16),
7730 => conv_std_logic_vector(1500, 16),
7731 => conv_std_logic_vector(1530, 16),
7732 => conv_std_logic_vector(1560, 16),
7733 => conv_std_logic_vector(1590, 16),
7734 => conv_std_logic_vector(1620, 16),
7735 => conv_std_logic_vector(1650, 16),
7736 => conv_std_logic_vector(1680, 16),
7737 => conv_std_logic_vector(1710, 16),
7738 => conv_std_logic_vector(1740, 16),
7739 => conv_std_logic_vector(1770, 16),
7740 => conv_std_logic_vector(1800, 16),
7741 => conv_std_logic_vector(1830, 16),
7742 => conv_std_logic_vector(1860, 16),
7743 => conv_std_logic_vector(1890, 16),
7744 => conv_std_logic_vector(1920, 16),
7745 => conv_std_logic_vector(1950, 16),
7746 => conv_std_logic_vector(1980, 16),
7747 => conv_std_logic_vector(2010, 16),
7748 => conv_std_logic_vector(2040, 16),
7749 => conv_std_logic_vector(2070, 16),
7750 => conv_std_logic_vector(2100, 16),
7751 => conv_std_logic_vector(2130, 16),
7752 => conv_std_logic_vector(2160, 16),
7753 => conv_std_logic_vector(2190, 16),
7754 => conv_std_logic_vector(2220, 16),
7755 => conv_std_logic_vector(2250, 16),
7756 => conv_std_logic_vector(2280, 16),
7757 => conv_std_logic_vector(2310, 16),
7758 => conv_std_logic_vector(2340, 16),
7759 => conv_std_logic_vector(2370, 16),
7760 => conv_std_logic_vector(2400, 16),
7761 => conv_std_logic_vector(2430, 16),
7762 => conv_std_logic_vector(2460, 16),
7763 => conv_std_logic_vector(2490, 16),
7764 => conv_std_logic_vector(2520, 16),
7765 => conv_std_logic_vector(2550, 16),
7766 => conv_std_logic_vector(2580, 16),
7767 => conv_std_logic_vector(2610, 16),
7768 => conv_std_logic_vector(2640, 16),
7769 => conv_std_logic_vector(2670, 16),
7770 => conv_std_logic_vector(2700, 16),
7771 => conv_std_logic_vector(2730, 16),
7772 => conv_std_logic_vector(2760, 16),
7773 => conv_std_logic_vector(2790, 16),
7774 => conv_std_logic_vector(2820, 16),
7775 => conv_std_logic_vector(2850, 16),
7776 => conv_std_logic_vector(2880, 16),
7777 => conv_std_logic_vector(2910, 16),
7778 => conv_std_logic_vector(2940, 16),
7779 => conv_std_logic_vector(2970, 16),
7780 => conv_std_logic_vector(3000, 16),
7781 => conv_std_logic_vector(3030, 16),
7782 => conv_std_logic_vector(3060, 16),
7783 => conv_std_logic_vector(3090, 16),
7784 => conv_std_logic_vector(3120, 16),
7785 => conv_std_logic_vector(3150, 16),
7786 => conv_std_logic_vector(3180, 16),
7787 => conv_std_logic_vector(3210, 16),
7788 => conv_std_logic_vector(3240, 16),
7789 => conv_std_logic_vector(3270, 16),
7790 => conv_std_logic_vector(3300, 16),
7791 => conv_std_logic_vector(3330, 16),
7792 => conv_std_logic_vector(3360, 16),
7793 => conv_std_logic_vector(3390, 16),
7794 => conv_std_logic_vector(3420, 16),
7795 => conv_std_logic_vector(3450, 16),
7796 => conv_std_logic_vector(3480, 16),
7797 => conv_std_logic_vector(3510, 16),
7798 => conv_std_logic_vector(3540, 16),
7799 => conv_std_logic_vector(3570, 16),
7800 => conv_std_logic_vector(3600, 16),
7801 => conv_std_logic_vector(3630, 16),
7802 => conv_std_logic_vector(3660, 16),
7803 => conv_std_logic_vector(3690, 16),
7804 => conv_std_logic_vector(3720, 16),
7805 => conv_std_logic_vector(3750, 16),
7806 => conv_std_logic_vector(3780, 16),
7807 => conv_std_logic_vector(3810, 16),
7808 => conv_std_logic_vector(3840, 16),
7809 => conv_std_logic_vector(3870, 16),
7810 => conv_std_logic_vector(3900, 16),
7811 => conv_std_logic_vector(3930, 16),
7812 => conv_std_logic_vector(3960, 16),
7813 => conv_std_logic_vector(3990, 16),
7814 => conv_std_logic_vector(4020, 16),
7815 => conv_std_logic_vector(4050, 16),
7816 => conv_std_logic_vector(4080, 16),
7817 => conv_std_logic_vector(4110, 16),
7818 => conv_std_logic_vector(4140, 16),
7819 => conv_std_logic_vector(4170, 16),
7820 => conv_std_logic_vector(4200, 16),
7821 => conv_std_logic_vector(4230, 16),
7822 => conv_std_logic_vector(4260, 16),
7823 => conv_std_logic_vector(4290, 16),
7824 => conv_std_logic_vector(4320, 16),
7825 => conv_std_logic_vector(4350, 16),
7826 => conv_std_logic_vector(4380, 16),
7827 => conv_std_logic_vector(4410, 16),
7828 => conv_std_logic_vector(4440, 16),
7829 => conv_std_logic_vector(4470, 16),
7830 => conv_std_logic_vector(4500, 16),
7831 => conv_std_logic_vector(4530, 16),
7832 => conv_std_logic_vector(4560, 16),
7833 => conv_std_logic_vector(4590, 16),
7834 => conv_std_logic_vector(4620, 16),
7835 => conv_std_logic_vector(4650, 16),
7836 => conv_std_logic_vector(4680, 16),
7837 => conv_std_logic_vector(4710, 16),
7838 => conv_std_logic_vector(4740, 16),
7839 => conv_std_logic_vector(4770, 16),
7840 => conv_std_logic_vector(4800, 16),
7841 => conv_std_logic_vector(4830, 16),
7842 => conv_std_logic_vector(4860, 16),
7843 => conv_std_logic_vector(4890, 16),
7844 => conv_std_logic_vector(4920, 16),
7845 => conv_std_logic_vector(4950, 16),
7846 => conv_std_logic_vector(4980, 16),
7847 => conv_std_logic_vector(5010, 16),
7848 => conv_std_logic_vector(5040, 16),
7849 => conv_std_logic_vector(5070, 16),
7850 => conv_std_logic_vector(5100, 16),
7851 => conv_std_logic_vector(5130, 16),
7852 => conv_std_logic_vector(5160, 16),
7853 => conv_std_logic_vector(5190, 16),
7854 => conv_std_logic_vector(5220, 16),
7855 => conv_std_logic_vector(5250, 16),
7856 => conv_std_logic_vector(5280, 16),
7857 => conv_std_logic_vector(5310, 16),
7858 => conv_std_logic_vector(5340, 16),
7859 => conv_std_logic_vector(5370, 16),
7860 => conv_std_logic_vector(5400, 16),
7861 => conv_std_logic_vector(5430, 16),
7862 => conv_std_logic_vector(5460, 16),
7863 => conv_std_logic_vector(5490, 16),
7864 => conv_std_logic_vector(5520, 16),
7865 => conv_std_logic_vector(5550, 16),
7866 => conv_std_logic_vector(5580, 16),
7867 => conv_std_logic_vector(5610, 16),
7868 => conv_std_logic_vector(5640, 16),
7869 => conv_std_logic_vector(5670, 16),
7870 => conv_std_logic_vector(5700, 16),
7871 => conv_std_logic_vector(5730, 16),
7872 => conv_std_logic_vector(5760, 16),
7873 => conv_std_logic_vector(5790, 16),
7874 => conv_std_logic_vector(5820, 16),
7875 => conv_std_logic_vector(5850, 16),
7876 => conv_std_logic_vector(5880, 16),
7877 => conv_std_logic_vector(5910, 16),
7878 => conv_std_logic_vector(5940, 16),
7879 => conv_std_logic_vector(5970, 16),
7880 => conv_std_logic_vector(6000, 16),
7881 => conv_std_logic_vector(6030, 16),
7882 => conv_std_logic_vector(6060, 16),
7883 => conv_std_logic_vector(6090, 16),
7884 => conv_std_logic_vector(6120, 16),
7885 => conv_std_logic_vector(6150, 16),
7886 => conv_std_logic_vector(6180, 16),
7887 => conv_std_logic_vector(6210, 16),
7888 => conv_std_logic_vector(6240, 16),
7889 => conv_std_logic_vector(6270, 16),
7890 => conv_std_logic_vector(6300, 16),
7891 => conv_std_logic_vector(6330, 16),
7892 => conv_std_logic_vector(6360, 16),
7893 => conv_std_logic_vector(6390, 16),
7894 => conv_std_logic_vector(6420, 16),
7895 => conv_std_logic_vector(6450, 16),
7896 => conv_std_logic_vector(6480, 16),
7897 => conv_std_logic_vector(6510, 16),
7898 => conv_std_logic_vector(6540, 16),
7899 => conv_std_logic_vector(6570, 16),
7900 => conv_std_logic_vector(6600, 16),
7901 => conv_std_logic_vector(6630, 16),
7902 => conv_std_logic_vector(6660, 16),
7903 => conv_std_logic_vector(6690, 16),
7904 => conv_std_logic_vector(6720, 16),
7905 => conv_std_logic_vector(6750, 16),
7906 => conv_std_logic_vector(6780, 16),
7907 => conv_std_logic_vector(6810, 16),
7908 => conv_std_logic_vector(6840, 16),
7909 => conv_std_logic_vector(6870, 16),
7910 => conv_std_logic_vector(6900, 16),
7911 => conv_std_logic_vector(6930, 16),
7912 => conv_std_logic_vector(6960, 16),
7913 => conv_std_logic_vector(6990, 16),
7914 => conv_std_logic_vector(7020, 16),
7915 => conv_std_logic_vector(7050, 16),
7916 => conv_std_logic_vector(7080, 16),
7917 => conv_std_logic_vector(7110, 16),
7918 => conv_std_logic_vector(7140, 16),
7919 => conv_std_logic_vector(7170, 16),
7920 => conv_std_logic_vector(7200, 16),
7921 => conv_std_logic_vector(7230, 16),
7922 => conv_std_logic_vector(7260, 16),
7923 => conv_std_logic_vector(7290, 16),
7924 => conv_std_logic_vector(7320, 16),
7925 => conv_std_logic_vector(7350, 16),
7926 => conv_std_logic_vector(7380, 16),
7927 => conv_std_logic_vector(7410, 16),
7928 => conv_std_logic_vector(7440, 16),
7929 => conv_std_logic_vector(7470, 16),
7930 => conv_std_logic_vector(7500, 16),
7931 => conv_std_logic_vector(7530, 16),
7932 => conv_std_logic_vector(7560, 16),
7933 => conv_std_logic_vector(7590, 16),
7934 => conv_std_logic_vector(7620, 16),
7935 => conv_std_logic_vector(7650, 16),
7936 => conv_std_logic_vector(0, 16),
7937 => conv_std_logic_vector(31, 16),
7938 => conv_std_logic_vector(62, 16),
7939 => conv_std_logic_vector(93, 16),
7940 => conv_std_logic_vector(124, 16),
7941 => conv_std_logic_vector(155, 16),
7942 => conv_std_logic_vector(186, 16),
7943 => conv_std_logic_vector(217, 16),
7944 => conv_std_logic_vector(248, 16),
7945 => conv_std_logic_vector(279, 16),
7946 => conv_std_logic_vector(310, 16),
7947 => conv_std_logic_vector(341, 16),
7948 => conv_std_logic_vector(372, 16),
7949 => conv_std_logic_vector(403, 16),
7950 => conv_std_logic_vector(434, 16),
7951 => conv_std_logic_vector(465, 16),
7952 => conv_std_logic_vector(496, 16),
7953 => conv_std_logic_vector(527, 16),
7954 => conv_std_logic_vector(558, 16),
7955 => conv_std_logic_vector(589, 16),
7956 => conv_std_logic_vector(620, 16),
7957 => conv_std_logic_vector(651, 16),
7958 => conv_std_logic_vector(682, 16),
7959 => conv_std_logic_vector(713, 16),
7960 => conv_std_logic_vector(744, 16),
7961 => conv_std_logic_vector(775, 16),
7962 => conv_std_logic_vector(806, 16),
7963 => conv_std_logic_vector(837, 16),
7964 => conv_std_logic_vector(868, 16),
7965 => conv_std_logic_vector(899, 16),
7966 => conv_std_logic_vector(930, 16),
7967 => conv_std_logic_vector(961, 16),
7968 => conv_std_logic_vector(992, 16),
7969 => conv_std_logic_vector(1023, 16),
7970 => conv_std_logic_vector(1054, 16),
7971 => conv_std_logic_vector(1085, 16),
7972 => conv_std_logic_vector(1116, 16),
7973 => conv_std_logic_vector(1147, 16),
7974 => conv_std_logic_vector(1178, 16),
7975 => conv_std_logic_vector(1209, 16),
7976 => conv_std_logic_vector(1240, 16),
7977 => conv_std_logic_vector(1271, 16),
7978 => conv_std_logic_vector(1302, 16),
7979 => conv_std_logic_vector(1333, 16),
7980 => conv_std_logic_vector(1364, 16),
7981 => conv_std_logic_vector(1395, 16),
7982 => conv_std_logic_vector(1426, 16),
7983 => conv_std_logic_vector(1457, 16),
7984 => conv_std_logic_vector(1488, 16),
7985 => conv_std_logic_vector(1519, 16),
7986 => conv_std_logic_vector(1550, 16),
7987 => conv_std_logic_vector(1581, 16),
7988 => conv_std_logic_vector(1612, 16),
7989 => conv_std_logic_vector(1643, 16),
7990 => conv_std_logic_vector(1674, 16),
7991 => conv_std_logic_vector(1705, 16),
7992 => conv_std_logic_vector(1736, 16),
7993 => conv_std_logic_vector(1767, 16),
7994 => conv_std_logic_vector(1798, 16),
7995 => conv_std_logic_vector(1829, 16),
7996 => conv_std_logic_vector(1860, 16),
7997 => conv_std_logic_vector(1891, 16),
7998 => conv_std_logic_vector(1922, 16),
7999 => conv_std_logic_vector(1953, 16),
8000 => conv_std_logic_vector(1984, 16),
8001 => conv_std_logic_vector(2015, 16),
8002 => conv_std_logic_vector(2046, 16),
8003 => conv_std_logic_vector(2077, 16),
8004 => conv_std_logic_vector(2108, 16),
8005 => conv_std_logic_vector(2139, 16),
8006 => conv_std_logic_vector(2170, 16),
8007 => conv_std_logic_vector(2201, 16),
8008 => conv_std_logic_vector(2232, 16),
8009 => conv_std_logic_vector(2263, 16),
8010 => conv_std_logic_vector(2294, 16),
8011 => conv_std_logic_vector(2325, 16),
8012 => conv_std_logic_vector(2356, 16),
8013 => conv_std_logic_vector(2387, 16),
8014 => conv_std_logic_vector(2418, 16),
8015 => conv_std_logic_vector(2449, 16),
8016 => conv_std_logic_vector(2480, 16),
8017 => conv_std_logic_vector(2511, 16),
8018 => conv_std_logic_vector(2542, 16),
8019 => conv_std_logic_vector(2573, 16),
8020 => conv_std_logic_vector(2604, 16),
8021 => conv_std_logic_vector(2635, 16),
8022 => conv_std_logic_vector(2666, 16),
8023 => conv_std_logic_vector(2697, 16),
8024 => conv_std_logic_vector(2728, 16),
8025 => conv_std_logic_vector(2759, 16),
8026 => conv_std_logic_vector(2790, 16),
8027 => conv_std_logic_vector(2821, 16),
8028 => conv_std_logic_vector(2852, 16),
8029 => conv_std_logic_vector(2883, 16),
8030 => conv_std_logic_vector(2914, 16),
8031 => conv_std_logic_vector(2945, 16),
8032 => conv_std_logic_vector(2976, 16),
8033 => conv_std_logic_vector(3007, 16),
8034 => conv_std_logic_vector(3038, 16),
8035 => conv_std_logic_vector(3069, 16),
8036 => conv_std_logic_vector(3100, 16),
8037 => conv_std_logic_vector(3131, 16),
8038 => conv_std_logic_vector(3162, 16),
8039 => conv_std_logic_vector(3193, 16),
8040 => conv_std_logic_vector(3224, 16),
8041 => conv_std_logic_vector(3255, 16),
8042 => conv_std_logic_vector(3286, 16),
8043 => conv_std_logic_vector(3317, 16),
8044 => conv_std_logic_vector(3348, 16),
8045 => conv_std_logic_vector(3379, 16),
8046 => conv_std_logic_vector(3410, 16),
8047 => conv_std_logic_vector(3441, 16),
8048 => conv_std_logic_vector(3472, 16),
8049 => conv_std_logic_vector(3503, 16),
8050 => conv_std_logic_vector(3534, 16),
8051 => conv_std_logic_vector(3565, 16),
8052 => conv_std_logic_vector(3596, 16),
8053 => conv_std_logic_vector(3627, 16),
8054 => conv_std_logic_vector(3658, 16),
8055 => conv_std_logic_vector(3689, 16),
8056 => conv_std_logic_vector(3720, 16),
8057 => conv_std_logic_vector(3751, 16),
8058 => conv_std_logic_vector(3782, 16),
8059 => conv_std_logic_vector(3813, 16),
8060 => conv_std_logic_vector(3844, 16),
8061 => conv_std_logic_vector(3875, 16),
8062 => conv_std_logic_vector(3906, 16),
8063 => conv_std_logic_vector(3937, 16),
8064 => conv_std_logic_vector(3968, 16),
8065 => conv_std_logic_vector(3999, 16),
8066 => conv_std_logic_vector(4030, 16),
8067 => conv_std_logic_vector(4061, 16),
8068 => conv_std_logic_vector(4092, 16),
8069 => conv_std_logic_vector(4123, 16),
8070 => conv_std_logic_vector(4154, 16),
8071 => conv_std_logic_vector(4185, 16),
8072 => conv_std_logic_vector(4216, 16),
8073 => conv_std_logic_vector(4247, 16),
8074 => conv_std_logic_vector(4278, 16),
8075 => conv_std_logic_vector(4309, 16),
8076 => conv_std_logic_vector(4340, 16),
8077 => conv_std_logic_vector(4371, 16),
8078 => conv_std_logic_vector(4402, 16),
8079 => conv_std_logic_vector(4433, 16),
8080 => conv_std_logic_vector(4464, 16),
8081 => conv_std_logic_vector(4495, 16),
8082 => conv_std_logic_vector(4526, 16),
8083 => conv_std_logic_vector(4557, 16),
8084 => conv_std_logic_vector(4588, 16),
8085 => conv_std_logic_vector(4619, 16),
8086 => conv_std_logic_vector(4650, 16),
8087 => conv_std_logic_vector(4681, 16),
8088 => conv_std_logic_vector(4712, 16),
8089 => conv_std_logic_vector(4743, 16),
8090 => conv_std_logic_vector(4774, 16),
8091 => conv_std_logic_vector(4805, 16),
8092 => conv_std_logic_vector(4836, 16),
8093 => conv_std_logic_vector(4867, 16),
8094 => conv_std_logic_vector(4898, 16),
8095 => conv_std_logic_vector(4929, 16),
8096 => conv_std_logic_vector(4960, 16),
8097 => conv_std_logic_vector(4991, 16),
8098 => conv_std_logic_vector(5022, 16),
8099 => conv_std_logic_vector(5053, 16),
8100 => conv_std_logic_vector(5084, 16),
8101 => conv_std_logic_vector(5115, 16),
8102 => conv_std_logic_vector(5146, 16),
8103 => conv_std_logic_vector(5177, 16),
8104 => conv_std_logic_vector(5208, 16),
8105 => conv_std_logic_vector(5239, 16),
8106 => conv_std_logic_vector(5270, 16),
8107 => conv_std_logic_vector(5301, 16),
8108 => conv_std_logic_vector(5332, 16),
8109 => conv_std_logic_vector(5363, 16),
8110 => conv_std_logic_vector(5394, 16),
8111 => conv_std_logic_vector(5425, 16),
8112 => conv_std_logic_vector(5456, 16),
8113 => conv_std_logic_vector(5487, 16),
8114 => conv_std_logic_vector(5518, 16),
8115 => conv_std_logic_vector(5549, 16),
8116 => conv_std_logic_vector(5580, 16),
8117 => conv_std_logic_vector(5611, 16),
8118 => conv_std_logic_vector(5642, 16),
8119 => conv_std_logic_vector(5673, 16),
8120 => conv_std_logic_vector(5704, 16),
8121 => conv_std_logic_vector(5735, 16),
8122 => conv_std_logic_vector(5766, 16),
8123 => conv_std_logic_vector(5797, 16),
8124 => conv_std_logic_vector(5828, 16),
8125 => conv_std_logic_vector(5859, 16),
8126 => conv_std_logic_vector(5890, 16),
8127 => conv_std_logic_vector(5921, 16),
8128 => conv_std_logic_vector(5952, 16),
8129 => conv_std_logic_vector(5983, 16),
8130 => conv_std_logic_vector(6014, 16),
8131 => conv_std_logic_vector(6045, 16),
8132 => conv_std_logic_vector(6076, 16),
8133 => conv_std_logic_vector(6107, 16),
8134 => conv_std_logic_vector(6138, 16),
8135 => conv_std_logic_vector(6169, 16),
8136 => conv_std_logic_vector(6200, 16),
8137 => conv_std_logic_vector(6231, 16),
8138 => conv_std_logic_vector(6262, 16),
8139 => conv_std_logic_vector(6293, 16),
8140 => conv_std_logic_vector(6324, 16),
8141 => conv_std_logic_vector(6355, 16),
8142 => conv_std_logic_vector(6386, 16),
8143 => conv_std_logic_vector(6417, 16),
8144 => conv_std_logic_vector(6448, 16),
8145 => conv_std_logic_vector(6479, 16),
8146 => conv_std_logic_vector(6510, 16),
8147 => conv_std_logic_vector(6541, 16),
8148 => conv_std_logic_vector(6572, 16),
8149 => conv_std_logic_vector(6603, 16),
8150 => conv_std_logic_vector(6634, 16),
8151 => conv_std_logic_vector(6665, 16),
8152 => conv_std_logic_vector(6696, 16),
8153 => conv_std_logic_vector(6727, 16),
8154 => conv_std_logic_vector(6758, 16),
8155 => conv_std_logic_vector(6789, 16),
8156 => conv_std_logic_vector(6820, 16),
8157 => conv_std_logic_vector(6851, 16),
8158 => conv_std_logic_vector(6882, 16),
8159 => conv_std_logic_vector(6913, 16),
8160 => conv_std_logic_vector(6944, 16),
8161 => conv_std_logic_vector(6975, 16),
8162 => conv_std_logic_vector(7006, 16),
8163 => conv_std_logic_vector(7037, 16),
8164 => conv_std_logic_vector(7068, 16),
8165 => conv_std_logic_vector(7099, 16),
8166 => conv_std_logic_vector(7130, 16),
8167 => conv_std_logic_vector(7161, 16),
8168 => conv_std_logic_vector(7192, 16),
8169 => conv_std_logic_vector(7223, 16),
8170 => conv_std_logic_vector(7254, 16),
8171 => conv_std_logic_vector(7285, 16),
8172 => conv_std_logic_vector(7316, 16),
8173 => conv_std_logic_vector(7347, 16),
8174 => conv_std_logic_vector(7378, 16),
8175 => conv_std_logic_vector(7409, 16),
8176 => conv_std_logic_vector(7440, 16),
8177 => conv_std_logic_vector(7471, 16),
8178 => conv_std_logic_vector(7502, 16),
8179 => conv_std_logic_vector(7533, 16),
8180 => conv_std_logic_vector(7564, 16),
8181 => conv_std_logic_vector(7595, 16),
8182 => conv_std_logic_vector(7626, 16),
8183 => conv_std_logic_vector(7657, 16),
8184 => conv_std_logic_vector(7688, 16),
8185 => conv_std_logic_vector(7719, 16),
8186 => conv_std_logic_vector(7750, 16),
8187 => conv_std_logic_vector(7781, 16),
8188 => conv_std_logic_vector(7812, 16),
8189 => conv_std_logic_vector(7843, 16),
8190 => conv_std_logic_vector(7874, 16),
8191 => conv_std_logic_vector(7905, 16),
8192 => conv_std_logic_vector(0, 16),
8193 => conv_std_logic_vector(32, 16),
8194 => conv_std_logic_vector(64, 16),
8195 => conv_std_logic_vector(96, 16),
8196 => conv_std_logic_vector(128, 16),
8197 => conv_std_logic_vector(160, 16),
8198 => conv_std_logic_vector(192, 16),
8199 => conv_std_logic_vector(224, 16),
8200 => conv_std_logic_vector(256, 16),
8201 => conv_std_logic_vector(288, 16),
8202 => conv_std_logic_vector(320, 16),
8203 => conv_std_logic_vector(352, 16),
8204 => conv_std_logic_vector(384, 16),
8205 => conv_std_logic_vector(416, 16),
8206 => conv_std_logic_vector(448, 16),
8207 => conv_std_logic_vector(480, 16),
8208 => conv_std_logic_vector(512, 16),
8209 => conv_std_logic_vector(544, 16),
8210 => conv_std_logic_vector(576, 16),
8211 => conv_std_logic_vector(608, 16),
8212 => conv_std_logic_vector(640, 16),
8213 => conv_std_logic_vector(672, 16),
8214 => conv_std_logic_vector(704, 16),
8215 => conv_std_logic_vector(736, 16),
8216 => conv_std_logic_vector(768, 16),
8217 => conv_std_logic_vector(800, 16),
8218 => conv_std_logic_vector(832, 16),
8219 => conv_std_logic_vector(864, 16),
8220 => conv_std_logic_vector(896, 16),
8221 => conv_std_logic_vector(928, 16),
8222 => conv_std_logic_vector(960, 16),
8223 => conv_std_logic_vector(992, 16),
8224 => conv_std_logic_vector(1024, 16),
8225 => conv_std_logic_vector(1056, 16),
8226 => conv_std_logic_vector(1088, 16),
8227 => conv_std_logic_vector(1120, 16),
8228 => conv_std_logic_vector(1152, 16),
8229 => conv_std_logic_vector(1184, 16),
8230 => conv_std_logic_vector(1216, 16),
8231 => conv_std_logic_vector(1248, 16),
8232 => conv_std_logic_vector(1280, 16),
8233 => conv_std_logic_vector(1312, 16),
8234 => conv_std_logic_vector(1344, 16),
8235 => conv_std_logic_vector(1376, 16),
8236 => conv_std_logic_vector(1408, 16),
8237 => conv_std_logic_vector(1440, 16),
8238 => conv_std_logic_vector(1472, 16),
8239 => conv_std_logic_vector(1504, 16),
8240 => conv_std_logic_vector(1536, 16),
8241 => conv_std_logic_vector(1568, 16),
8242 => conv_std_logic_vector(1600, 16),
8243 => conv_std_logic_vector(1632, 16),
8244 => conv_std_logic_vector(1664, 16),
8245 => conv_std_logic_vector(1696, 16),
8246 => conv_std_logic_vector(1728, 16),
8247 => conv_std_logic_vector(1760, 16),
8248 => conv_std_logic_vector(1792, 16),
8249 => conv_std_logic_vector(1824, 16),
8250 => conv_std_logic_vector(1856, 16),
8251 => conv_std_logic_vector(1888, 16),
8252 => conv_std_logic_vector(1920, 16),
8253 => conv_std_logic_vector(1952, 16),
8254 => conv_std_logic_vector(1984, 16),
8255 => conv_std_logic_vector(2016, 16),
8256 => conv_std_logic_vector(2048, 16),
8257 => conv_std_logic_vector(2080, 16),
8258 => conv_std_logic_vector(2112, 16),
8259 => conv_std_logic_vector(2144, 16),
8260 => conv_std_logic_vector(2176, 16),
8261 => conv_std_logic_vector(2208, 16),
8262 => conv_std_logic_vector(2240, 16),
8263 => conv_std_logic_vector(2272, 16),
8264 => conv_std_logic_vector(2304, 16),
8265 => conv_std_logic_vector(2336, 16),
8266 => conv_std_logic_vector(2368, 16),
8267 => conv_std_logic_vector(2400, 16),
8268 => conv_std_logic_vector(2432, 16),
8269 => conv_std_logic_vector(2464, 16),
8270 => conv_std_logic_vector(2496, 16),
8271 => conv_std_logic_vector(2528, 16),
8272 => conv_std_logic_vector(2560, 16),
8273 => conv_std_logic_vector(2592, 16),
8274 => conv_std_logic_vector(2624, 16),
8275 => conv_std_logic_vector(2656, 16),
8276 => conv_std_logic_vector(2688, 16),
8277 => conv_std_logic_vector(2720, 16),
8278 => conv_std_logic_vector(2752, 16),
8279 => conv_std_logic_vector(2784, 16),
8280 => conv_std_logic_vector(2816, 16),
8281 => conv_std_logic_vector(2848, 16),
8282 => conv_std_logic_vector(2880, 16),
8283 => conv_std_logic_vector(2912, 16),
8284 => conv_std_logic_vector(2944, 16),
8285 => conv_std_logic_vector(2976, 16),
8286 => conv_std_logic_vector(3008, 16),
8287 => conv_std_logic_vector(3040, 16),
8288 => conv_std_logic_vector(3072, 16),
8289 => conv_std_logic_vector(3104, 16),
8290 => conv_std_logic_vector(3136, 16),
8291 => conv_std_logic_vector(3168, 16),
8292 => conv_std_logic_vector(3200, 16),
8293 => conv_std_logic_vector(3232, 16),
8294 => conv_std_logic_vector(3264, 16),
8295 => conv_std_logic_vector(3296, 16),
8296 => conv_std_logic_vector(3328, 16),
8297 => conv_std_logic_vector(3360, 16),
8298 => conv_std_logic_vector(3392, 16),
8299 => conv_std_logic_vector(3424, 16),
8300 => conv_std_logic_vector(3456, 16),
8301 => conv_std_logic_vector(3488, 16),
8302 => conv_std_logic_vector(3520, 16),
8303 => conv_std_logic_vector(3552, 16),
8304 => conv_std_logic_vector(3584, 16),
8305 => conv_std_logic_vector(3616, 16),
8306 => conv_std_logic_vector(3648, 16),
8307 => conv_std_logic_vector(3680, 16),
8308 => conv_std_logic_vector(3712, 16),
8309 => conv_std_logic_vector(3744, 16),
8310 => conv_std_logic_vector(3776, 16),
8311 => conv_std_logic_vector(3808, 16),
8312 => conv_std_logic_vector(3840, 16),
8313 => conv_std_logic_vector(3872, 16),
8314 => conv_std_logic_vector(3904, 16),
8315 => conv_std_logic_vector(3936, 16),
8316 => conv_std_logic_vector(3968, 16),
8317 => conv_std_logic_vector(4000, 16),
8318 => conv_std_logic_vector(4032, 16),
8319 => conv_std_logic_vector(4064, 16),
8320 => conv_std_logic_vector(4096, 16),
8321 => conv_std_logic_vector(4128, 16),
8322 => conv_std_logic_vector(4160, 16),
8323 => conv_std_logic_vector(4192, 16),
8324 => conv_std_logic_vector(4224, 16),
8325 => conv_std_logic_vector(4256, 16),
8326 => conv_std_logic_vector(4288, 16),
8327 => conv_std_logic_vector(4320, 16),
8328 => conv_std_logic_vector(4352, 16),
8329 => conv_std_logic_vector(4384, 16),
8330 => conv_std_logic_vector(4416, 16),
8331 => conv_std_logic_vector(4448, 16),
8332 => conv_std_logic_vector(4480, 16),
8333 => conv_std_logic_vector(4512, 16),
8334 => conv_std_logic_vector(4544, 16),
8335 => conv_std_logic_vector(4576, 16),
8336 => conv_std_logic_vector(4608, 16),
8337 => conv_std_logic_vector(4640, 16),
8338 => conv_std_logic_vector(4672, 16),
8339 => conv_std_logic_vector(4704, 16),
8340 => conv_std_logic_vector(4736, 16),
8341 => conv_std_logic_vector(4768, 16),
8342 => conv_std_logic_vector(4800, 16),
8343 => conv_std_logic_vector(4832, 16),
8344 => conv_std_logic_vector(4864, 16),
8345 => conv_std_logic_vector(4896, 16),
8346 => conv_std_logic_vector(4928, 16),
8347 => conv_std_logic_vector(4960, 16),
8348 => conv_std_logic_vector(4992, 16),
8349 => conv_std_logic_vector(5024, 16),
8350 => conv_std_logic_vector(5056, 16),
8351 => conv_std_logic_vector(5088, 16),
8352 => conv_std_logic_vector(5120, 16),
8353 => conv_std_logic_vector(5152, 16),
8354 => conv_std_logic_vector(5184, 16),
8355 => conv_std_logic_vector(5216, 16),
8356 => conv_std_logic_vector(5248, 16),
8357 => conv_std_logic_vector(5280, 16),
8358 => conv_std_logic_vector(5312, 16),
8359 => conv_std_logic_vector(5344, 16),
8360 => conv_std_logic_vector(5376, 16),
8361 => conv_std_logic_vector(5408, 16),
8362 => conv_std_logic_vector(5440, 16),
8363 => conv_std_logic_vector(5472, 16),
8364 => conv_std_logic_vector(5504, 16),
8365 => conv_std_logic_vector(5536, 16),
8366 => conv_std_logic_vector(5568, 16),
8367 => conv_std_logic_vector(5600, 16),
8368 => conv_std_logic_vector(5632, 16),
8369 => conv_std_logic_vector(5664, 16),
8370 => conv_std_logic_vector(5696, 16),
8371 => conv_std_logic_vector(5728, 16),
8372 => conv_std_logic_vector(5760, 16),
8373 => conv_std_logic_vector(5792, 16),
8374 => conv_std_logic_vector(5824, 16),
8375 => conv_std_logic_vector(5856, 16),
8376 => conv_std_logic_vector(5888, 16),
8377 => conv_std_logic_vector(5920, 16),
8378 => conv_std_logic_vector(5952, 16),
8379 => conv_std_logic_vector(5984, 16),
8380 => conv_std_logic_vector(6016, 16),
8381 => conv_std_logic_vector(6048, 16),
8382 => conv_std_logic_vector(6080, 16),
8383 => conv_std_logic_vector(6112, 16),
8384 => conv_std_logic_vector(6144, 16),
8385 => conv_std_logic_vector(6176, 16),
8386 => conv_std_logic_vector(6208, 16),
8387 => conv_std_logic_vector(6240, 16),
8388 => conv_std_logic_vector(6272, 16),
8389 => conv_std_logic_vector(6304, 16),
8390 => conv_std_logic_vector(6336, 16),
8391 => conv_std_logic_vector(6368, 16),
8392 => conv_std_logic_vector(6400, 16),
8393 => conv_std_logic_vector(6432, 16),
8394 => conv_std_logic_vector(6464, 16),
8395 => conv_std_logic_vector(6496, 16),
8396 => conv_std_logic_vector(6528, 16),
8397 => conv_std_logic_vector(6560, 16),
8398 => conv_std_logic_vector(6592, 16),
8399 => conv_std_logic_vector(6624, 16),
8400 => conv_std_logic_vector(6656, 16),
8401 => conv_std_logic_vector(6688, 16),
8402 => conv_std_logic_vector(6720, 16),
8403 => conv_std_logic_vector(6752, 16),
8404 => conv_std_logic_vector(6784, 16),
8405 => conv_std_logic_vector(6816, 16),
8406 => conv_std_logic_vector(6848, 16),
8407 => conv_std_logic_vector(6880, 16),
8408 => conv_std_logic_vector(6912, 16),
8409 => conv_std_logic_vector(6944, 16),
8410 => conv_std_logic_vector(6976, 16),
8411 => conv_std_logic_vector(7008, 16),
8412 => conv_std_logic_vector(7040, 16),
8413 => conv_std_logic_vector(7072, 16),
8414 => conv_std_logic_vector(7104, 16),
8415 => conv_std_logic_vector(7136, 16),
8416 => conv_std_logic_vector(7168, 16),
8417 => conv_std_logic_vector(7200, 16),
8418 => conv_std_logic_vector(7232, 16),
8419 => conv_std_logic_vector(7264, 16),
8420 => conv_std_logic_vector(7296, 16),
8421 => conv_std_logic_vector(7328, 16),
8422 => conv_std_logic_vector(7360, 16),
8423 => conv_std_logic_vector(7392, 16),
8424 => conv_std_logic_vector(7424, 16),
8425 => conv_std_logic_vector(7456, 16),
8426 => conv_std_logic_vector(7488, 16),
8427 => conv_std_logic_vector(7520, 16),
8428 => conv_std_logic_vector(7552, 16),
8429 => conv_std_logic_vector(7584, 16),
8430 => conv_std_logic_vector(7616, 16),
8431 => conv_std_logic_vector(7648, 16),
8432 => conv_std_logic_vector(7680, 16),
8433 => conv_std_logic_vector(7712, 16),
8434 => conv_std_logic_vector(7744, 16),
8435 => conv_std_logic_vector(7776, 16),
8436 => conv_std_logic_vector(7808, 16),
8437 => conv_std_logic_vector(7840, 16),
8438 => conv_std_logic_vector(7872, 16),
8439 => conv_std_logic_vector(7904, 16),
8440 => conv_std_logic_vector(7936, 16),
8441 => conv_std_logic_vector(7968, 16),
8442 => conv_std_logic_vector(8000, 16),
8443 => conv_std_logic_vector(8032, 16),
8444 => conv_std_logic_vector(8064, 16),
8445 => conv_std_logic_vector(8096, 16),
8446 => conv_std_logic_vector(8128, 16),
8447 => conv_std_logic_vector(8160, 16),
8448 => conv_std_logic_vector(0, 16),
8449 => conv_std_logic_vector(33, 16),
8450 => conv_std_logic_vector(66, 16),
8451 => conv_std_logic_vector(99, 16),
8452 => conv_std_logic_vector(132, 16),
8453 => conv_std_logic_vector(165, 16),
8454 => conv_std_logic_vector(198, 16),
8455 => conv_std_logic_vector(231, 16),
8456 => conv_std_logic_vector(264, 16),
8457 => conv_std_logic_vector(297, 16),
8458 => conv_std_logic_vector(330, 16),
8459 => conv_std_logic_vector(363, 16),
8460 => conv_std_logic_vector(396, 16),
8461 => conv_std_logic_vector(429, 16),
8462 => conv_std_logic_vector(462, 16),
8463 => conv_std_logic_vector(495, 16),
8464 => conv_std_logic_vector(528, 16),
8465 => conv_std_logic_vector(561, 16),
8466 => conv_std_logic_vector(594, 16),
8467 => conv_std_logic_vector(627, 16),
8468 => conv_std_logic_vector(660, 16),
8469 => conv_std_logic_vector(693, 16),
8470 => conv_std_logic_vector(726, 16),
8471 => conv_std_logic_vector(759, 16),
8472 => conv_std_logic_vector(792, 16),
8473 => conv_std_logic_vector(825, 16),
8474 => conv_std_logic_vector(858, 16),
8475 => conv_std_logic_vector(891, 16),
8476 => conv_std_logic_vector(924, 16),
8477 => conv_std_logic_vector(957, 16),
8478 => conv_std_logic_vector(990, 16),
8479 => conv_std_logic_vector(1023, 16),
8480 => conv_std_logic_vector(1056, 16),
8481 => conv_std_logic_vector(1089, 16),
8482 => conv_std_logic_vector(1122, 16),
8483 => conv_std_logic_vector(1155, 16),
8484 => conv_std_logic_vector(1188, 16),
8485 => conv_std_logic_vector(1221, 16),
8486 => conv_std_logic_vector(1254, 16),
8487 => conv_std_logic_vector(1287, 16),
8488 => conv_std_logic_vector(1320, 16),
8489 => conv_std_logic_vector(1353, 16),
8490 => conv_std_logic_vector(1386, 16),
8491 => conv_std_logic_vector(1419, 16),
8492 => conv_std_logic_vector(1452, 16),
8493 => conv_std_logic_vector(1485, 16),
8494 => conv_std_logic_vector(1518, 16),
8495 => conv_std_logic_vector(1551, 16),
8496 => conv_std_logic_vector(1584, 16),
8497 => conv_std_logic_vector(1617, 16),
8498 => conv_std_logic_vector(1650, 16),
8499 => conv_std_logic_vector(1683, 16),
8500 => conv_std_logic_vector(1716, 16),
8501 => conv_std_logic_vector(1749, 16),
8502 => conv_std_logic_vector(1782, 16),
8503 => conv_std_logic_vector(1815, 16),
8504 => conv_std_logic_vector(1848, 16),
8505 => conv_std_logic_vector(1881, 16),
8506 => conv_std_logic_vector(1914, 16),
8507 => conv_std_logic_vector(1947, 16),
8508 => conv_std_logic_vector(1980, 16),
8509 => conv_std_logic_vector(2013, 16),
8510 => conv_std_logic_vector(2046, 16),
8511 => conv_std_logic_vector(2079, 16),
8512 => conv_std_logic_vector(2112, 16),
8513 => conv_std_logic_vector(2145, 16),
8514 => conv_std_logic_vector(2178, 16),
8515 => conv_std_logic_vector(2211, 16),
8516 => conv_std_logic_vector(2244, 16),
8517 => conv_std_logic_vector(2277, 16),
8518 => conv_std_logic_vector(2310, 16),
8519 => conv_std_logic_vector(2343, 16),
8520 => conv_std_logic_vector(2376, 16),
8521 => conv_std_logic_vector(2409, 16),
8522 => conv_std_logic_vector(2442, 16),
8523 => conv_std_logic_vector(2475, 16),
8524 => conv_std_logic_vector(2508, 16),
8525 => conv_std_logic_vector(2541, 16),
8526 => conv_std_logic_vector(2574, 16),
8527 => conv_std_logic_vector(2607, 16),
8528 => conv_std_logic_vector(2640, 16),
8529 => conv_std_logic_vector(2673, 16),
8530 => conv_std_logic_vector(2706, 16),
8531 => conv_std_logic_vector(2739, 16),
8532 => conv_std_logic_vector(2772, 16),
8533 => conv_std_logic_vector(2805, 16),
8534 => conv_std_logic_vector(2838, 16),
8535 => conv_std_logic_vector(2871, 16),
8536 => conv_std_logic_vector(2904, 16),
8537 => conv_std_logic_vector(2937, 16),
8538 => conv_std_logic_vector(2970, 16),
8539 => conv_std_logic_vector(3003, 16),
8540 => conv_std_logic_vector(3036, 16),
8541 => conv_std_logic_vector(3069, 16),
8542 => conv_std_logic_vector(3102, 16),
8543 => conv_std_logic_vector(3135, 16),
8544 => conv_std_logic_vector(3168, 16),
8545 => conv_std_logic_vector(3201, 16),
8546 => conv_std_logic_vector(3234, 16),
8547 => conv_std_logic_vector(3267, 16),
8548 => conv_std_logic_vector(3300, 16),
8549 => conv_std_logic_vector(3333, 16),
8550 => conv_std_logic_vector(3366, 16),
8551 => conv_std_logic_vector(3399, 16),
8552 => conv_std_logic_vector(3432, 16),
8553 => conv_std_logic_vector(3465, 16),
8554 => conv_std_logic_vector(3498, 16),
8555 => conv_std_logic_vector(3531, 16),
8556 => conv_std_logic_vector(3564, 16),
8557 => conv_std_logic_vector(3597, 16),
8558 => conv_std_logic_vector(3630, 16),
8559 => conv_std_logic_vector(3663, 16),
8560 => conv_std_logic_vector(3696, 16),
8561 => conv_std_logic_vector(3729, 16),
8562 => conv_std_logic_vector(3762, 16),
8563 => conv_std_logic_vector(3795, 16),
8564 => conv_std_logic_vector(3828, 16),
8565 => conv_std_logic_vector(3861, 16),
8566 => conv_std_logic_vector(3894, 16),
8567 => conv_std_logic_vector(3927, 16),
8568 => conv_std_logic_vector(3960, 16),
8569 => conv_std_logic_vector(3993, 16),
8570 => conv_std_logic_vector(4026, 16),
8571 => conv_std_logic_vector(4059, 16),
8572 => conv_std_logic_vector(4092, 16),
8573 => conv_std_logic_vector(4125, 16),
8574 => conv_std_logic_vector(4158, 16),
8575 => conv_std_logic_vector(4191, 16),
8576 => conv_std_logic_vector(4224, 16),
8577 => conv_std_logic_vector(4257, 16),
8578 => conv_std_logic_vector(4290, 16),
8579 => conv_std_logic_vector(4323, 16),
8580 => conv_std_logic_vector(4356, 16),
8581 => conv_std_logic_vector(4389, 16),
8582 => conv_std_logic_vector(4422, 16),
8583 => conv_std_logic_vector(4455, 16),
8584 => conv_std_logic_vector(4488, 16),
8585 => conv_std_logic_vector(4521, 16),
8586 => conv_std_logic_vector(4554, 16),
8587 => conv_std_logic_vector(4587, 16),
8588 => conv_std_logic_vector(4620, 16),
8589 => conv_std_logic_vector(4653, 16),
8590 => conv_std_logic_vector(4686, 16),
8591 => conv_std_logic_vector(4719, 16),
8592 => conv_std_logic_vector(4752, 16),
8593 => conv_std_logic_vector(4785, 16),
8594 => conv_std_logic_vector(4818, 16),
8595 => conv_std_logic_vector(4851, 16),
8596 => conv_std_logic_vector(4884, 16),
8597 => conv_std_logic_vector(4917, 16),
8598 => conv_std_logic_vector(4950, 16),
8599 => conv_std_logic_vector(4983, 16),
8600 => conv_std_logic_vector(5016, 16),
8601 => conv_std_logic_vector(5049, 16),
8602 => conv_std_logic_vector(5082, 16),
8603 => conv_std_logic_vector(5115, 16),
8604 => conv_std_logic_vector(5148, 16),
8605 => conv_std_logic_vector(5181, 16),
8606 => conv_std_logic_vector(5214, 16),
8607 => conv_std_logic_vector(5247, 16),
8608 => conv_std_logic_vector(5280, 16),
8609 => conv_std_logic_vector(5313, 16),
8610 => conv_std_logic_vector(5346, 16),
8611 => conv_std_logic_vector(5379, 16),
8612 => conv_std_logic_vector(5412, 16),
8613 => conv_std_logic_vector(5445, 16),
8614 => conv_std_logic_vector(5478, 16),
8615 => conv_std_logic_vector(5511, 16),
8616 => conv_std_logic_vector(5544, 16),
8617 => conv_std_logic_vector(5577, 16),
8618 => conv_std_logic_vector(5610, 16),
8619 => conv_std_logic_vector(5643, 16),
8620 => conv_std_logic_vector(5676, 16),
8621 => conv_std_logic_vector(5709, 16),
8622 => conv_std_logic_vector(5742, 16),
8623 => conv_std_logic_vector(5775, 16),
8624 => conv_std_logic_vector(5808, 16),
8625 => conv_std_logic_vector(5841, 16),
8626 => conv_std_logic_vector(5874, 16),
8627 => conv_std_logic_vector(5907, 16),
8628 => conv_std_logic_vector(5940, 16),
8629 => conv_std_logic_vector(5973, 16),
8630 => conv_std_logic_vector(6006, 16),
8631 => conv_std_logic_vector(6039, 16),
8632 => conv_std_logic_vector(6072, 16),
8633 => conv_std_logic_vector(6105, 16),
8634 => conv_std_logic_vector(6138, 16),
8635 => conv_std_logic_vector(6171, 16),
8636 => conv_std_logic_vector(6204, 16),
8637 => conv_std_logic_vector(6237, 16),
8638 => conv_std_logic_vector(6270, 16),
8639 => conv_std_logic_vector(6303, 16),
8640 => conv_std_logic_vector(6336, 16),
8641 => conv_std_logic_vector(6369, 16),
8642 => conv_std_logic_vector(6402, 16),
8643 => conv_std_logic_vector(6435, 16),
8644 => conv_std_logic_vector(6468, 16),
8645 => conv_std_logic_vector(6501, 16),
8646 => conv_std_logic_vector(6534, 16),
8647 => conv_std_logic_vector(6567, 16),
8648 => conv_std_logic_vector(6600, 16),
8649 => conv_std_logic_vector(6633, 16),
8650 => conv_std_logic_vector(6666, 16),
8651 => conv_std_logic_vector(6699, 16),
8652 => conv_std_logic_vector(6732, 16),
8653 => conv_std_logic_vector(6765, 16),
8654 => conv_std_logic_vector(6798, 16),
8655 => conv_std_logic_vector(6831, 16),
8656 => conv_std_logic_vector(6864, 16),
8657 => conv_std_logic_vector(6897, 16),
8658 => conv_std_logic_vector(6930, 16),
8659 => conv_std_logic_vector(6963, 16),
8660 => conv_std_logic_vector(6996, 16),
8661 => conv_std_logic_vector(7029, 16),
8662 => conv_std_logic_vector(7062, 16),
8663 => conv_std_logic_vector(7095, 16),
8664 => conv_std_logic_vector(7128, 16),
8665 => conv_std_logic_vector(7161, 16),
8666 => conv_std_logic_vector(7194, 16),
8667 => conv_std_logic_vector(7227, 16),
8668 => conv_std_logic_vector(7260, 16),
8669 => conv_std_logic_vector(7293, 16),
8670 => conv_std_logic_vector(7326, 16),
8671 => conv_std_logic_vector(7359, 16),
8672 => conv_std_logic_vector(7392, 16),
8673 => conv_std_logic_vector(7425, 16),
8674 => conv_std_logic_vector(7458, 16),
8675 => conv_std_logic_vector(7491, 16),
8676 => conv_std_logic_vector(7524, 16),
8677 => conv_std_logic_vector(7557, 16),
8678 => conv_std_logic_vector(7590, 16),
8679 => conv_std_logic_vector(7623, 16),
8680 => conv_std_logic_vector(7656, 16),
8681 => conv_std_logic_vector(7689, 16),
8682 => conv_std_logic_vector(7722, 16),
8683 => conv_std_logic_vector(7755, 16),
8684 => conv_std_logic_vector(7788, 16),
8685 => conv_std_logic_vector(7821, 16),
8686 => conv_std_logic_vector(7854, 16),
8687 => conv_std_logic_vector(7887, 16),
8688 => conv_std_logic_vector(7920, 16),
8689 => conv_std_logic_vector(7953, 16),
8690 => conv_std_logic_vector(7986, 16),
8691 => conv_std_logic_vector(8019, 16),
8692 => conv_std_logic_vector(8052, 16),
8693 => conv_std_logic_vector(8085, 16),
8694 => conv_std_logic_vector(8118, 16),
8695 => conv_std_logic_vector(8151, 16),
8696 => conv_std_logic_vector(8184, 16),
8697 => conv_std_logic_vector(8217, 16),
8698 => conv_std_logic_vector(8250, 16),
8699 => conv_std_logic_vector(8283, 16),
8700 => conv_std_logic_vector(8316, 16),
8701 => conv_std_logic_vector(8349, 16),
8702 => conv_std_logic_vector(8382, 16),
8703 => conv_std_logic_vector(8415, 16),
8704 => conv_std_logic_vector(0, 16),
8705 => conv_std_logic_vector(34, 16),
8706 => conv_std_logic_vector(68, 16),
8707 => conv_std_logic_vector(102, 16),
8708 => conv_std_logic_vector(136, 16),
8709 => conv_std_logic_vector(170, 16),
8710 => conv_std_logic_vector(204, 16),
8711 => conv_std_logic_vector(238, 16),
8712 => conv_std_logic_vector(272, 16),
8713 => conv_std_logic_vector(306, 16),
8714 => conv_std_logic_vector(340, 16),
8715 => conv_std_logic_vector(374, 16),
8716 => conv_std_logic_vector(408, 16),
8717 => conv_std_logic_vector(442, 16),
8718 => conv_std_logic_vector(476, 16),
8719 => conv_std_logic_vector(510, 16),
8720 => conv_std_logic_vector(544, 16),
8721 => conv_std_logic_vector(578, 16),
8722 => conv_std_logic_vector(612, 16),
8723 => conv_std_logic_vector(646, 16),
8724 => conv_std_logic_vector(680, 16),
8725 => conv_std_logic_vector(714, 16),
8726 => conv_std_logic_vector(748, 16),
8727 => conv_std_logic_vector(782, 16),
8728 => conv_std_logic_vector(816, 16),
8729 => conv_std_logic_vector(850, 16),
8730 => conv_std_logic_vector(884, 16),
8731 => conv_std_logic_vector(918, 16),
8732 => conv_std_logic_vector(952, 16),
8733 => conv_std_logic_vector(986, 16),
8734 => conv_std_logic_vector(1020, 16),
8735 => conv_std_logic_vector(1054, 16),
8736 => conv_std_logic_vector(1088, 16),
8737 => conv_std_logic_vector(1122, 16),
8738 => conv_std_logic_vector(1156, 16),
8739 => conv_std_logic_vector(1190, 16),
8740 => conv_std_logic_vector(1224, 16),
8741 => conv_std_logic_vector(1258, 16),
8742 => conv_std_logic_vector(1292, 16),
8743 => conv_std_logic_vector(1326, 16),
8744 => conv_std_logic_vector(1360, 16),
8745 => conv_std_logic_vector(1394, 16),
8746 => conv_std_logic_vector(1428, 16),
8747 => conv_std_logic_vector(1462, 16),
8748 => conv_std_logic_vector(1496, 16),
8749 => conv_std_logic_vector(1530, 16),
8750 => conv_std_logic_vector(1564, 16),
8751 => conv_std_logic_vector(1598, 16),
8752 => conv_std_logic_vector(1632, 16),
8753 => conv_std_logic_vector(1666, 16),
8754 => conv_std_logic_vector(1700, 16),
8755 => conv_std_logic_vector(1734, 16),
8756 => conv_std_logic_vector(1768, 16),
8757 => conv_std_logic_vector(1802, 16),
8758 => conv_std_logic_vector(1836, 16),
8759 => conv_std_logic_vector(1870, 16),
8760 => conv_std_logic_vector(1904, 16),
8761 => conv_std_logic_vector(1938, 16),
8762 => conv_std_logic_vector(1972, 16),
8763 => conv_std_logic_vector(2006, 16),
8764 => conv_std_logic_vector(2040, 16),
8765 => conv_std_logic_vector(2074, 16),
8766 => conv_std_logic_vector(2108, 16),
8767 => conv_std_logic_vector(2142, 16),
8768 => conv_std_logic_vector(2176, 16),
8769 => conv_std_logic_vector(2210, 16),
8770 => conv_std_logic_vector(2244, 16),
8771 => conv_std_logic_vector(2278, 16),
8772 => conv_std_logic_vector(2312, 16),
8773 => conv_std_logic_vector(2346, 16),
8774 => conv_std_logic_vector(2380, 16),
8775 => conv_std_logic_vector(2414, 16),
8776 => conv_std_logic_vector(2448, 16),
8777 => conv_std_logic_vector(2482, 16),
8778 => conv_std_logic_vector(2516, 16),
8779 => conv_std_logic_vector(2550, 16),
8780 => conv_std_logic_vector(2584, 16),
8781 => conv_std_logic_vector(2618, 16),
8782 => conv_std_logic_vector(2652, 16),
8783 => conv_std_logic_vector(2686, 16),
8784 => conv_std_logic_vector(2720, 16),
8785 => conv_std_logic_vector(2754, 16),
8786 => conv_std_logic_vector(2788, 16),
8787 => conv_std_logic_vector(2822, 16),
8788 => conv_std_logic_vector(2856, 16),
8789 => conv_std_logic_vector(2890, 16),
8790 => conv_std_logic_vector(2924, 16),
8791 => conv_std_logic_vector(2958, 16),
8792 => conv_std_logic_vector(2992, 16),
8793 => conv_std_logic_vector(3026, 16),
8794 => conv_std_logic_vector(3060, 16),
8795 => conv_std_logic_vector(3094, 16),
8796 => conv_std_logic_vector(3128, 16),
8797 => conv_std_logic_vector(3162, 16),
8798 => conv_std_logic_vector(3196, 16),
8799 => conv_std_logic_vector(3230, 16),
8800 => conv_std_logic_vector(3264, 16),
8801 => conv_std_logic_vector(3298, 16),
8802 => conv_std_logic_vector(3332, 16),
8803 => conv_std_logic_vector(3366, 16),
8804 => conv_std_logic_vector(3400, 16),
8805 => conv_std_logic_vector(3434, 16),
8806 => conv_std_logic_vector(3468, 16),
8807 => conv_std_logic_vector(3502, 16),
8808 => conv_std_logic_vector(3536, 16),
8809 => conv_std_logic_vector(3570, 16),
8810 => conv_std_logic_vector(3604, 16),
8811 => conv_std_logic_vector(3638, 16),
8812 => conv_std_logic_vector(3672, 16),
8813 => conv_std_logic_vector(3706, 16),
8814 => conv_std_logic_vector(3740, 16),
8815 => conv_std_logic_vector(3774, 16),
8816 => conv_std_logic_vector(3808, 16),
8817 => conv_std_logic_vector(3842, 16),
8818 => conv_std_logic_vector(3876, 16),
8819 => conv_std_logic_vector(3910, 16),
8820 => conv_std_logic_vector(3944, 16),
8821 => conv_std_logic_vector(3978, 16),
8822 => conv_std_logic_vector(4012, 16),
8823 => conv_std_logic_vector(4046, 16),
8824 => conv_std_logic_vector(4080, 16),
8825 => conv_std_logic_vector(4114, 16),
8826 => conv_std_logic_vector(4148, 16),
8827 => conv_std_logic_vector(4182, 16),
8828 => conv_std_logic_vector(4216, 16),
8829 => conv_std_logic_vector(4250, 16),
8830 => conv_std_logic_vector(4284, 16),
8831 => conv_std_logic_vector(4318, 16),
8832 => conv_std_logic_vector(4352, 16),
8833 => conv_std_logic_vector(4386, 16),
8834 => conv_std_logic_vector(4420, 16),
8835 => conv_std_logic_vector(4454, 16),
8836 => conv_std_logic_vector(4488, 16),
8837 => conv_std_logic_vector(4522, 16),
8838 => conv_std_logic_vector(4556, 16),
8839 => conv_std_logic_vector(4590, 16),
8840 => conv_std_logic_vector(4624, 16),
8841 => conv_std_logic_vector(4658, 16),
8842 => conv_std_logic_vector(4692, 16),
8843 => conv_std_logic_vector(4726, 16),
8844 => conv_std_logic_vector(4760, 16),
8845 => conv_std_logic_vector(4794, 16),
8846 => conv_std_logic_vector(4828, 16),
8847 => conv_std_logic_vector(4862, 16),
8848 => conv_std_logic_vector(4896, 16),
8849 => conv_std_logic_vector(4930, 16),
8850 => conv_std_logic_vector(4964, 16),
8851 => conv_std_logic_vector(4998, 16),
8852 => conv_std_logic_vector(5032, 16),
8853 => conv_std_logic_vector(5066, 16),
8854 => conv_std_logic_vector(5100, 16),
8855 => conv_std_logic_vector(5134, 16),
8856 => conv_std_logic_vector(5168, 16),
8857 => conv_std_logic_vector(5202, 16),
8858 => conv_std_logic_vector(5236, 16),
8859 => conv_std_logic_vector(5270, 16),
8860 => conv_std_logic_vector(5304, 16),
8861 => conv_std_logic_vector(5338, 16),
8862 => conv_std_logic_vector(5372, 16),
8863 => conv_std_logic_vector(5406, 16),
8864 => conv_std_logic_vector(5440, 16),
8865 => conv_std_logic_vector(5474, 16),
8866 => conv_std_logic_vector(5508, 16),
8867 => conv_std_logic_vector(5542, 16),
8868 => conv_std_logic_vector(5576, 16),
8869 => conv_std_logic_vector(5610, 16),
8870 => conv_std_logic_vector(5644, 16),
8871 => conv_std_logic_vector(5678, 16),
8872 => conv_std_logic_vector(5712, 16),
8873 => conv_std_logic_vector(5746, 16),
8874 => conv_std_logic_vector(5780, 16),
8875 => conv_std_logic_vector(5814, 16),
8876 => conv_std_logic_vector(5848, 16),
8877 => conv_std_logic_vector(5882, 16),
8878 => conv_std_logic_vector(5916, 16),
8879 => conv_std_logic_vector(5950, 16),
8880 => conv_std_logic_vector(5984, 16),
8881 => conv_std_logic_vector(6018, 16),
8882 => conv_std_logic_vector(6052, 16),
8883 => conv_std_logic_vector(6086, 16),
8884 => conv_std_logic_vector(6120, 16),
8885 => conv_std_logic_vector(6154, 16),
8886 => conv_std_logic_vector(6188, 16),
8887 => conv_std_logic_vector(6222, 16),
8888 => conv_std_logic_vector(6256, 16),
8889 => conv_std_logic_vector(6290, 16),
8890 => conv_std_logic_vector(6324, 16),
8891 => conv_std_logic_vector(6358, 16),
8892 => conv_std_logic_vector(6392, 16),
8893 => conv_std_logic_vector(6426, 16),
8894 => conv_std_logic_vector(6460, 16),
8895 => conv_std_logic_vector(6494, 16),
8896 => conv_std_logic_vector(6528, 16),
8897 => conv_std_logic_vector(6562, 16),
8898 => conv_std_logic_vector(6596, 16),
8899 => conv_std_logic_vector(6630, 16),
8900 => conv_std_logic_vector(6664, 16),
8901 => conv_std_logic_vector(6698, 16),
8902 => conv_std_logic_vector(6732, 16),
8903 => conv_std_logic_vector(6766, 16),
8904 => conv_std_logic_vector(6800, 16),
8905 => conv_std_logic_vector(6834, 16),
8906 => conv_std_logic_vector(6868, 16),
8907 => conv_std_logic_vector(6902, 16),
8908 => conv_std_logic_vector(6936, 16),
8909 => conv_std_logic_vector(6970, 16),
8910 => conv_std_logic_vector(7004, 16),
8911 => conv_std_logic_vector(7038, 16),
8912 => conv_std_logic_vector(7072, 16),
8913 => conv_std_logic_vector(7106, 16),
8914 => conv_std_logic_vector(7140, 16),
8915 => conv_std_logic_vector(7174, 16),
8916 => conv_std_logic_vector(7208, 16),
8917 => conv_std_logic_vector(7242, 16),
8918 => conv_std_logic_vector(7276, 16),
8919 => conv_std_logic_vector(7310, 16),
8920 => conv_std_logic_vector(7344, 16),
8921 => conv_std_logic_vector(7378, 16),
8922 => conv_std_logic_vector(7412, 16),
8923 => conv_std_logic_vector(7446, 16),
8924 => conv_std_logic_vector(7480, 16),
8925 => conv_std_logic_vector(7514, 16),
8926 => conv_std_logic_vector(7548, 16),
8927 => conv_std_logic_vector(7582, 16),
8928 => conv_std_logic_vector(7616, 16),
8929 => conv_std_logic_vector(7650, 16),
8930 => conv_std_logic_vector(7684, 16),
8931 => conv_std_logic_vector(7718, 16),
8932 => conv_std_logic_vector(7752, 16),
8933 => conv_std_logic_vector(7786, 16),
8934 => conv_std_logic_vector(7820, 16),
8935 => conv_std_logic_vector(7854, 16),
8936 => conv_std_logic_vector(7888, 16),
8937 => conv_std_logic_vector(7922, 16),
8938 => conv_std_logic_vector(7956, 16),
8939 => conv_std_logic_vector(7990, 16),
8940 => conv_std_logic_vector(8024, 16),
8941 => conv_std_logic_vector(8058, 16),
8942 => conv_std_logic_vector(8092, 16),
8943 => conv_std_logic_vector(8126, 16),
8944 => conv_std_logic_vector(8160, 16),
8945 => conv_std_logic_vector(8194, 16),
8946 => conv_std_logic_vector(8228, 16),
8947 => conv_std_logic_vector(8262, 16),
8948 => conv_std_logic_vector(8296, 16),
8949 => conv_std_logic_vector(8330, 16),
8950 => conv_std_logic_vector(8364, 16),
8951 => conv_std_logic_vector(8398, 16),
8952 => conv_std_logic_vector(8432, 16),
8953 => conv_std_logic_vector(8466, 16),
8954 => conv_std_logic_vector(8500, 16),
8955 => conv_std_logic_vector(8534, 16),
8956 => conv_std_logic_vector(8568, 16),
8957 => conv_std_logic_vector(8602, 16),
8958 => conv_std_logic_vector(8636, 16),
8959 => conv_std_logic_vector(8670, 16),
8960 => conv_std_logic_vector(0, 16),
8961 => conv_std_logic_vector(35, 16),
8962 => conv_std_logic_vector(70, 16),
8963 => conv_std_logic_vector(105, 16),
8964 => conv_std_logic_vector(140, 16),
8965 => conv_std_logic_vector(175, 16),
8966 => conv_std_logic_vector(210, 16),
8967 => conv_std_logic_vector(245, 16),
8968 => conv_std_logic_vector(280, 16),
8969 => conv_std_logic_vector(315, 16),
8970 => conv_std_logic_vector(350, 16),
8971 => conv_std_logic_vector(385, 16),
8972 => conv_std_logic_vector(420, 16),
8973 => conv_std_logic_vector(455, 16),
8974 => conv_std_logic_vector(490, 16),
8975 => conv_std_logic_vector(525, 16),
8976 => conv_std_logic_vector(560, 16),
8977 => conv_std_logic_vector(595, 16),
8978 => conv_std_logic_vector(630, 16),
8979 => conv_std_logic_vector(665, 16),
8980 => conv_std_logic_vector(700, 16),
8981 => conv_std_logic_vector(735, 16),
8982 => conv_std_logic_vector(770, 16),
8983 => conv_std_logic_vector(805, 16),
8984 => conv_std_logic_vector(840, 16),
8985 => conv_std_logic_vector(875, 16),
8986 => conv_std_logic_vector(910, 16),
8987 => conv_std_logic_vector(945, 16),
8988 => conv_std_logic_vector(980, 16),
8989 => conv_std_logic_vector(1015, 16),
8990 => conv_std_logic_vector(1050, 16),
8991 => conv_std_logic_vector(1085, 16),
8992 => conv_std_logic_vector(1120, 16),
8993 => conv_std_logic_vector(1155, 16),
8994 => conv_std_logic_vector(1190, 16),
8995 => conv_std_logic_vector(1225, 16),
8996 => conv_std_logic_vector(1260, 16),
8997 => conv_std_logic_vector(1295, 16),
8998 => conv_std_logic_vector(1330, 16),
8999 => conv_std_logic_vector(1365, 16),
9000 => conv_std_logic_vector(1400, 16),
9001 => conv_std_logic_vector(1435, 16),
9002 => conv_std_logic_vector(1470, 16),
9003 => conv_std_logic_vector(1505, 16),
9004 => conv_std_logic_vector(1540, 16),
9005 => conv_std_logic_vector(1575, 16),
9006 => conv_std_logic_vector(1610, 16),
9007 => conv_std_logic_vector(1645, 16),
9008 => conv_std_logic_vector(1680, 16),
9009 => conv_std_logic_vector(1715, 16),
9010 => conv_std_logic_vector(1750, 16),
9011 => conv_std_logic_vector(1785, 16),
9012 => conv_std_logic_vector(1820, 16),
9013 => conv_std_logic_vector(1855, 16),
9014 => conv_std_logic_vector(1890, 16),
9015 => conv_std_logic_vector(1925, 16),
9016 => conv_std_logic_vector(1960, 16),
9017 => conv_std_logic_vector(1995, 16),
9018 => conv_std_logic_vector(2030, 16),
9019 => conv_std_logic_vector(2065, 16),
9020 => conv_std_logic_vector(2100, 16),
9021 => conv_std_logic_vector(2135, 16),
9022 => conv_std_logic_vector(2170, 16),
9023 => conv_std_logic_vector(2205, 16),
9024 => conv_std_logic_vector(2240, 16),
9025 => conv_std_logic_vector(2275, 16),
9026 => conv_std_logic_vector(2310, 16),
9027 => conv_std_logic_vector(2345, 16),
9028 => conv_std_logic_vector(2380, 16),
9029 => conv_std_logic_vector(2415, 16),
9030 => conv_std_logic_vector(2450, 16),
9031 => conv_std_logic_vector(2485, 16),
9032 => conv_std_logic_vector(2520, 16),
9033 => conv_std_logic_vector(2555, 16),
9034 => conv_std_logic_vector(2590, 16),
9035 => conv_std_logic_vector(2625, 16),
9036 => conv_std_logic_vector(2660, 16),
9037 => conv_std_logic_vector(2695, 16),
9038 => conv_std_logic_vector(2730, 16),
9039 => conv_std_logic_vector(2765, 16),
9040 => conv_std_logic_vector(2800, 16),
9041 => conv_std_logic_vector(2835, 16),
9042 => conv_std_logic_vector(2870, 16),
9043 => conv_std_logic_vector(2905, 16),
9044 => conv_std_logic_vector(2940, 16),
9045 => conv_std_logic_vector(2975, 16),
9046 => conv_std_logic_vector(3010, 16),
9047 => conv_std_logic_vector(3045, 16),
9048 => conv_std_logic_vector(3080, 16),
9049 => conv_std_logic_vector(3115, 16),
9050 => conv_std_logic_vector(3150, 16),
9051 => conv_std_logic_vector(3185, 16),
9052 => conv_std_logic_vector(3220, 16),
9053 => conv_std_logic_vector(3255, 16),
9054 => conv_std_logic_vector(3290, 16),
9055 => conv_std_logic_vector(3325, 16),
9056 => conv_std_logic_vector(3360, 16),
9057 => conv_std_logic_vector(3395, 16),
9058 => conv_std_logic_vector(3430, 16),
9059 => conv_std_logic_vector(3465, 16),
9060 => conv_std_logic_vector(3500, 16),
9061 => conv_std_logic_vector(3535, 16),
9062 => conv_std_logic_vector(3570, 16),
9063 => conv_std_logic_vector(3605, 16),
9064 => conv_std_logic_vector(3640, 16),
9065 => conv_std_logic_vector(3675, 16),
9066 => conv_std_logic_vector(3710, 16),
9067 => conv_std_logic_vector(3745, 16),
9068 => conv_std_logic_vector(3780, 16),
9069 => conv_std_logic_vector(3815, 16),
9070 => conv_std_logic_vector(3850, 16),
9071 => conv_std_logic_vector(3885, 16),
9072 => conv_std_logic_vector(3920, 16),
9073 => conv_std_logic_vector(3955, 16),
9074 => conv_std_logic_vector(3990, 16),
9075 => conv_std_logic_vector(4025, 16),
9076 => conv_std_logic_vector(4060, 16),
9077 => conv_std_logic_vector(4095, 16),
9078 => conv_std_logic_vector(4130, 16),
9079 => conv_std_logic_vector(4165, 16),
9080 => conv_std_logic_vector(4200, 16),
9081 => conv_std_logic_vector(4235, 16),
9082 => conv_std_logic_vector(4270, 16),
9083 => conv_std_logic_vector(4305, 16),
9084 => conv_std_logic_vector(4340, 16),
9085 => conv_std_logic_vector(4375, 16),
9086 => conv_std_logic_vector(4410, 16),
9087 => conv_std_logic_vector(4445, 16),
9088 => conv_std_logic_vector(4480, 16),
9089 => conv_std_logic_vector(4515, 16),
9090 => conv_std_logic_vector(4550, 16),
9091 => conv_std_logic_vector(4585, 16),
9092 => conv_std_logic_vector(4620, 16),
9093 => conv_std_logic_vector(4655, 16),
9094 => conv_std_logic_vector(4690, 16),
9095 => conv_std_logic_vector(4725, 16),
9096 => conv_std_logic_vector(4760, 16),
9097 => conv_std_logic_vector(4795, 16),
9098 => conv_std_logic_vector(4830, 16),
9099 => conv_std_logic_vector(4865, 16),
9100 => conv_std_logic_vector(4900, 16),
9101 => conv_std_logic_vector(4935, 16),
9102 => conv_std_logic_vector(4970, 16),
9103 => conv_std_logic_vector(5005, 16),
9104 => conv_std_logic_vector(5040, 16),
9105 => conv_std_logic_vector(5075, 16),
9106 => conv_std_logic_vector(5110, 16),
9107 => conv_std_logic_vector(5145, 16),
9108 => conv_std_logic_vector(5180, 16),
9109 => conv_std_logic_vector(5215, 16),
9110 => conv_std_logic_vector(5250, 16),
9111 => conv_std_logic_vector(5285, 16),
9112 => conv_std_logic_vector(5320, 16),
9113 => conv_std_logic_vector(5355, 16),
9114 => conv_std_logic_vector(5390, 16),
9115 => conv_std_logic_vector(5425, 16),
9116 => conv_std_logic_vector(5460, 16),
9117 => conv_std_logic_vector(5495, 16),
9118 => conv_std_logic_vector(5530, 16),
9119 => conv_std_logic_vector(5565, 16),
9120 => conv_std_logic_vector(5600, 16),
9121 => conv_std_logic_vector(5635, 16),
9122 => conv_std_logic_vector(5670, 16),
9123 => conv_std_logic_vector(5705, 16),
9124 => conv_std_logic_vector(5740, 16),
9125 => conv_std_logic_vector(5775, 16),
9126 => conv_std_logic_vector(5810, 16),
9127 => conv_std_logic_vector(5845, 16),
9128 => conv_std_logic_vector(5880, 16),
9129 => conv_std_logic_vector(5915, 16),
9130 => conv_std_logic_vector(5950, 16),
9131 => conv_std_logic_vector(5985, 16),
9132 => conv_std_logic_vector(6020, 16),
9133 => conv_std_logic_vector(6055, 16),
9134 => conv_std_logic_vector(6090, 16),
9135 => conv_std_logic_vector(6125, 16),
9136 => conv_std_logic_vector(6160, 16),
9137 => conv_std_logic_vector(6195, 16),
9138 => conv_std_logic_vector(6230, 16),
9139 => conv_std_logic_vector(6265, 16),
9140 => conv_std_logic_vector(6300, 16),
9141 => conv_std_logic_vector(6335, 16),
9142 => conv_std_logic_vector(6370, 16),
9143 => conv_std_logic_vector(6405, 16),
9144 => conv_std_logic_vector(6440, 16),
9145 => conv_std_logic_vector(6475, 16),
9146 => conv_std_logic_vector(6510, 16),
9147 => conv_std_logic_vector(6545, 16),
9148 => conv_std_logic_vector(6580, 16),
9149 => conv_std_logic_vector(6615, 16),
9150 => conv_std_logic_vector(6650, 16),
9151 => conv_std_logic_vector(6685, 16),
9152 => conv_std_logic_vector(6720, 16),
9153 => conv_std_logic_vector(6755, 16),
9154 => conv_std_logic_vector(6790, 16),
9155 => conv_std_logic_vector(6825, 16),
9156 => conv_std_logic_vector(6860, 16),
9157 => conv_std_logic_vector(6895, 16),
9158 => conv_std_logic_vector(6930, 16),
9159 => conv_std_logic_vector(6965, 16),
9160 => conv_std_logic_vector(7000, 16),
9161 => conv_std_logic_vector(7035, 16),
9162 => conv_std_logic_vector(7070, 16),
9163 => conv_std_logic_vector(7105, 16),
9164 => conv_std_logic_vector(7140, 16),
9165 => conv_std_logic_vector(7175, 16),
9166 => conv_std_logic_vector(7210, 16),
9167 => conv_std_logic_vector(7245, 16),
9168 => conv_std_logic_vector(7280, 16),
9169 => conv_std_logic_vector(7315, 16),
9170 => conv_std_logic_vector(7350, 16),
9171 => conv_std_logic_vector(7385, 16),
9172 => conv_std_logic_vector(7420, 16),
9173 => conv_std_logic_vector(7455, 16),
9174 => conv_std_logic_vector(7490, 16),
9175 => conv_std_logic_vector(7525, 16),
9176 => conv_std_logic_vector(7560, 16),
9177 => conv_std_logic_vector(7595, 16),
9178 => conv_std_logic_vector(7630, 16),
9179 => conv_std_logic_vector(7665, 16),
9180 => conv_std_logic_vector(7700, 16),
9181 => conv_std_logic_vector(7735, 16),
9182 => conv_std_logic_vector(7770, 16),
9183 => conv_std_logic_vector(7805, 16),
9184 => conv_std_logic_vector(7840, 16),
9185 => conv_std_logic_vector(7875, 16),
9186 => conv_std_logic_vector(7910, 16),
9187 => conv_std_logic_vector(7945, 16),
9188 => conv_std_logic_vector(7980, 16),
9189 => conv_std_logic_vector(8015, 16),
9190 => conv_std_logic_vector(8050, 16),
9191 => conv_std_logic_vector(8085, 16),
9192 => conv_std_logic_vector(8120, 16),
9193 => conv_std_logic_vector(8155, 16),
9194 => conv_std_logic_vector(8190, 16),
9195 => conv_std_logic_vector(8225, 16),
9196 => conv_std_logic_vector(8260, 16),
9197 => conv_std_logic_vector(8295, 16),
9198 => conv_std_logic_vector(8330, 16),
9199 => conv_std_logic_vector(8365, 16),
9200 => conv_std_logic_vector(8400, 16),
9201 => conv_std_logic_vector(8435, 16),
9202 => conv_std_logic_vector(8470, 16),
9203 => conv_std_logic_vector(8505, 16),
9204 => conv_std_logic_vector(8540, 16),
9205 => conv_std_logic_vector(8575, 16),
9206 => conv_std_logic_vector(8610, 16),
9207 => conv_std_logic_vector(8645, 16),
9208 => conv_std_logic_vector(8680, 16),
9209 => conv_std_logic_vector(8715, 16),
9210 => conv_std_logic_vector(8750, 16),
9211 => conv_std_logic_vector(8785, 16),
9212 => conv_std_logic_vector(8820, 16),
9213 => conv_std_logic_vector(8855, 16),
9214 => conv_std_logic_vector(8890, 16),
9215 => conv_std_logic_vector(8925, 16),
9216 => conv_std_logic_vector(0, 16),
9217 => conv_std_logic_vector(36, 16),
9218 => conv_std_logic_vector(72, 16),
9219 => conv_std_logic_vector(108, 16),
9220 => conv_std_logic_vector(144, 16),
9221 => conv_std_logic_vector(180, 16),
9222 => conv_std_logic_vector(216, 16),
9223 => conv_std_logic_vector(252, 16),
9224 => conv_std_logic_vector(288, 16),
9225 => conv_std_logic_vector(324, 16),
9226 => conv_std_logic_vector(360, 16),
9227 => conv_std_logic_vector(396, 16),
9228 => conv_std_logic_vector(432, 16),
9229 => conv_std_logic_vector(468, 16),
9230 => conv_std_logic_vector(504, 16),
9231 => conv_std_logic_vector(540, 16),
9232 => conv_std_logic_vector(576, 16),
9233 => conv_std_logic_vector(612, 16),
9234 => conv_std_logic_vector(648, 16),
9235 => conv_std_logic_vector(684, 16),
9236 => conv_std_logic_vector(720, 16),
9237 => conv_std_logic_vector(756, 16),
9238 => conv_std_logic_vector(792, 16),
9239 => conv_std_logic_vector(828, 16),
9240 => conv_std_logic_vector(864, 16),
9241 => conv_std_logic_vector(900, 16),
9242 => conv_std_logic_vector(936, 16),
9243 => conv_std_logic_vector(972, 16),
9244 => conv_std_logic_vector(1008, 16),
9245 => conv_std_logic_vector(1044, 16),
9246 => conv_std_logic_vector(1080, 16),
9247 => conv_std_logic_vector(1116, 16),
9248 => conv_std_logic_vector(1152, 16),
9249 => conv_std_logic_vector(1188, 16),
9250 => conv_std_logic_vector(1224, 16),
9251 => conv_std_logic_vector(1260, 16),
9252 => conv_std_logic_vector(1296, 16),
9253 => conv_std_logic_vector(1332, 16),
9254 => conv_std_logic_vector(1368, 16),
9255 => conv_std_logic_vector(1404, 16),
9256 => conv_std_logic_vector(1440, 16),
9257 => conv_std_logic_vector(1476, 16),
9258 => conv_std_logic_vector(1512, 16),
9259 => conv_std_logic_vector(1548, 16),
9260 => conv_std_logic_vector(1584, 16),
9261 => conv_std_logic_vector(1620, 16),
9262 => conv_std_logic_vector(1656, 16),
9263 => conv_std_logic_vector(1692, 16),
9264 => conv_std_logic_vector(1728, 16),
9265 => conv_std_logic_vector(1764, 16),
9266 => conv_std_logic_vector(1800, 16),
9267 => conv_std_logic_vector(1836, 16),
9268 => conv_std_logic_vector(1872, 16),
9269 => conv_std_logic_vector(1908, 16),
9270 => conv_std_logic_vector(1944, 16),
9271 => conv_std_logic_vector(1980, 16),
9272 => conv_std_logic_vector(2016, 16),
9273 => conv_std_logic_vector(2052, 16),
9274 => conv_std_logic_vector(2088, 16),
9275 => conv_std_logic_vector(2124, 16),
9276 => conv_std_logic_vector(2160, 16),
9277 => conv_std_logic_vector(2196, 16),
9278 => conv_std_logic_vector(2232, 16),
9279 => conv_std_logic_vector(2268, 16),
9280 => conv_std_logic_vector(2304, 16),
9281 => conv_std_logic_vector(2340, 16),
9282 => conv_std_logic_vector(2376, 16),
9283 => conv_std_logic_vector(2412, 16),
9284 => conv_std_logic_vector(2448, 16),
9285 => conv_std_logic_vector(2484, 16),
9286 => conv_std_logic_vector(2520, 16),
9287 => conv_std_logic_vector(2556, 16),
9288 => conv_std_logic_vector(2592, 16),
9289 => conv_std_logic_vector(2628, 16),
9290 => conv_std_logic_vector(2664, 16),
9291 => conv_std_logic_vector(2700, 16),
9292 => conv_std_logic_vector(2736, 16),
9293 => conv_std_logic_vector(2772, 16),
9294 => conv_std_logic_vector(2808, 16),
9295 => conv_std_logic_vector(2844, 16),
9296 => conv_std_logic_vector(2880, 16),
9297 => conv_std_logic_vector(2916, 16),
9298 => conv_std_logic_vector(2952, 16),
9299 => conv_std_logic_vector(2988, 16),
9300 => conv_std_logic_vector(3024, 16),
9301 => conv_std_logic_vector(3060, 16),
9302 => conv_std_logic_vector(3096, 16),
9303 => conv_std_logic_vector(3132, 16),
9304 => conv_std_logic_vector(3168, 16),
9305 => conv_std_logic_vector(3204, 16),
9306 => conv_std_logic_vector(3240, 16),
9307 => conv_std_logic_vector(3276, 16),
9308 => conv_std_logic_vector(3312, 16),
9309 => conv_std_logic_vector(3348, 16),
9310 => conv_std_logic_vector(3384, 16),
9311 => conv_std_logic_vector(3420, 16),
9312 => conv_std_logic_vector(3456, 16),
9313 => conv_std_logic_vector(3492, 16),
9314 => conv_std_logic_vector(3528, 16),
9315 => conv_std_logic_vector(3564, 16),
9316 => conv_std_logic_vector(3600, 16),
9317 => conv_std_logic_vector(3636, 16),
9318 => conv_std_logic_vector(3672, 16),
9319 => conv_std_logic_vector(3708, 16),
9320 => conv_std_logic_vector(3744, 16),
9321 => conv_std_logic_vector(3780, 16),
9322 => conv_std_logic_vector(3816, 16),
9323 => conv_std_logic_vector(3852, 16),
9324 => conv_std_logic_vector(3888, 16),
9325 => conv_std_logic_vector(3924, 16),
9326 => conv_std_logic_vector(3960, 16),
9327 => conv_std_logic_vector(3996, 16),
9328 => conv_std_logic_vector(4032, 16),
9329 => conv_std_logic_vector(4068, 16),
9330 => conv_std_logic_vector(4104, 16),
9331 => conv_std_logic_vector(4140, 16),
9332 => conv_std_logic_vector(4176, 16),
9333 => conv_std_logic_vector(4212, 16),
9334 => conv_std_logic_vector(4248, 16),
9335 => conv_std_logic_vector(4284, 16),
9336 => conv_std_logic_vector(4320, 16),
9337 => conv_std_logic_vector(4356, 16),
9338 => conv_std_logic_vector(4392, 16),
9339 => conv_std_logic_vector(4428, 16),
9340 => conv_std_logic_vector(4464, 16),
9341 => conv_std_logic_vector(4500, 16),
9342 => conv_std_logic_vector(4536, 16),
9343 => conv_std_logic_vector(4572, 16),
9344 => conv_std_logic_vector(4608, 16),
9345 => conv_std_logic_vector(4644, 16),
9346 => conv_std_logic_vector(4680, 16),
9347 => conv_std_logic_vector(4716, 16),
9348 => conv_std_logic_vector(4752, 16),
9349 => conv_std_logic_vector(4788, 16),
9350 => conv_std_logic_vector(4824, 16),
9351 => conv_std_logic_vector(4860, 16),
9352 => conv_std_logic_vector(4896, 16),
9353 => conv_std_logic_vector(4932, 16),
9354 => conv_std_logic_vector(4968, 16),
9355 => conv_std_logic_vector(5004, 16),
9356 => conv_std_logic_vector(5040, 16),
9357 => conv_std_logic_vector(5076, 16),
9358 => conv_std_logic_vector(5112, 16),
9359 => conv_std_logic_vector(5148, 16),
9360 => conv_std_logic_vector(5184, 16),
9361 => conv_std_logic_vector(5220, 16),
9362 => conv_std_logic_vector(5256, 16),
9363 => conv_std_logic_vector(5292, 16),
9364 => conv_std_logic_vector(5328, 16),
9365 => conv_std_logic_vector(5364, 16),
9366 => conv_std_logic_vector(5400, 16),
9367 => conv_std_logic_vector(5436, 16),
9368 => conv_std_logic_vector(5472, 16),
9369 => conv_std_logic_vector(5508, 16),
9370 => conv_std_logic_vector(5544, 16),
9371 => conv_std_logic_vector(5580, 16),
9372 => conv_std_logic_vector(5616, 16),
9373 => conv_std_logic_vector(5652, 16),
9374 => conv_std_logic_vector(5688, 16),
9375 => conv_std_logic_vector(5724, 16),
9376 => conv_std_logic_vector(5760, 16),
9377 => conv_std_logic_vector(5796, 16),
9378 => conv_std_logic_vector(5832, 16),
9379 => conv_std_logic_vector(5868, 16),
9380 => conv_std_logic_vector(5904, 16),
9381 => conv_std_logic_vector(5940, 16),
9382 => conv_std_logic_vector(5976, 16),
9383 => conv_std_logic_vector(6012, 16),
9384 => conv_std_logic_vector(6048, 16),
9385 => conv_std_logic_vector(6084, 16),
9386 => conv_std_logic_vector(6120, 16),
9387 => conv_std_logic_vector(6156, 16),
9388 => conv_std_logic_vector(6192, 16),
9389 => conv_std_logic_vector(6228, 16),
9390 => conv_std_logic_vector(6264, 16),
9391 => conv_std_logic_vector(6300, 16),
9392 => conv_std_logic_vector(6336, 16),
9393 => conv_std_logic_vector(6372, 16),
9394 => conv_std_logic_vector(6408, 16),
9395 => conv_std_logic_vector(6444, 16),
9396 => conv_std_logic_vector(6480, 16),
9397 => conv_std_logic_vector(6516, 16),
9398 => conv_std_logic_vector(6552, 16),
9399 => conv_std_logic_vector(6588, 16),
9400 => conv_std_logic_vector(6624, 16),
9401 => conv_std_logic_vector(6660, 16),
9402 => conv_std_logic_vector(6696, 16),
9403 => conv_std_logic_vector(6732, 16),
9404 => conv_std_logic_vector(6768, 16),
9405 => conv_std_logic_vector(6804, 16),
9406 => conv_std_logic_vector(6840, 16),
9407 => conv_std_logic_vector(6876, 16),
9408 => conv_std_logic_vector(6912, 16),
9409 => conv_std_logic_vector(6948, 16),
9410 => conv_std_logic_vector(6984, 16),
9411 => conv_std_logic_vector(7020, 16),
9412 => conv_std_logic_vector(7056, 16),
9413 => conv_std_logic_vector(7092, 16),
9414 => conv_std_logic_vector(7128, 16),
9415 => conv_std_logic_vector(7164, 16),
9416 => conv_std_logic_vector(7200, 16),
9417 => conv_std_logic_vector(7236, 16),
9418 => conv_std_logic_vector(7272, 16),
9419 => conv_std_logic_vector(7308, 16),
9420 => conv_std_logic_vector(7344, 16),
9421 => conv_std_logic_vector(7380, 16),
9422 => conv_std_logic_vector(7416, 16),
9423 => conv_std_logic_vector(7452, 16),
9424 => conv_std_logic_vector(7488, 16),
9425 => conv_std_logic_vector(7524, 16),
9426 => conv_std_logic_vector(7560, 16),
9427 => conv_std_logic_vector(7596, 16),
9428 => conv_std_logic_vector(7632, 16),
9429 => conv_std_logic_vector(7668, 16),
9430 => conv_std_logic_vector(7704, 16),
9431 => conv_std_logic_vector(7740, 16),
9432 => conv_std_logic_vector(7776, 16),
9433 => conv_std_logic_vector(7812, 16),
9434 => conv_std_logic_vector(7848, 16),
9435 => conv_std_logic_vector(7884, 16),
9436 => conv_std_logic_vector(7920, 16),
9437 => conv_std_logic_vector(7956, 16),
9438 => conv_std_logic_vector(7992, 16),
9439 => conv_std_logic_vector(8028, 16),
9440 => conv_std_logic_vector(8064, 16),
9441 => conv_std_logic_vector(8100, 16),
9442 => conv_std_logic_vector(8136, 16),
9443 => conv_std_logic_vector(8172, 16),
9444 => conv_std_logic_vector(8208, 16),
9445 => conv_std_logic_vector(8244, 16),
9446 => conv_std_logic_vector(8280, 16),
9447 => conv_std_logic_vector(8316, 16),
9448 => conv_std_logic_vector(8352, 16),
9449 => conv_std_logic_vector(8388, 16),
9450 => conv_std_logic_vector(8424, 16),
9451 => conv_std_logic_vector(8460, 16),
9452 => conv_std_logic_vector(8496, 16),
9453 => conv_std_logic_vector(8532, 16),
9454 => conv_std_logic_vector(8568, 16),
9455 => conv_std_logic_vector(8604, 16),
9456 => conv_std_logic_vector(8640, 16),
9457 => conv_std_logic_vector(8676, 16),
9458 => conv_std_logic_vector(8712, 16),
9459 => conv_std_logic_vector(8748, 16),
9460 => conv_std_logic_vector(8784, 16),
9461 => conv_std_logic_vector(8820, 16),
9462 => conv_std_logic_vector(8856, 16),
9463 => conv_std_logic_vector(8892, 16),
9464 => conv_std_logic_vector(8928, 16),
9465 => conv_std_logic_vector(8964, 16),
9466 => conv_std_logic_vector(9000, 16),
9467 => conv_std_logic_vector(9036, 16),
9468 => conv_std_logic_vector(9072, 16),
9469 => conv_std_logic_vector(9108, 16),
9470 => conv_std_logic_vector(9144, 16),
9471 => conv_std_logic_vector(9180, 16),
9472 => conv_std_logic_vector(0, 16),
9473 => conv_std_logic_vector(37, 16),
9474 => conv_std_logic_vector(74, 16),
9475 => conv_std_logic_vector(111, 16),
9476 => conv_std_logic_vector(148, 16),
9477 => conv_std_logic_vector(185, 16),
9478 => conv_std_logic_vector(222, 16),
9479 => conv_std_logic_vector(259, 16),
9480 => conv_std_logic_vector(296, 16),
9481 => conv_std_logic_vector(333, 16),
9482 => conv_std_logic_vector(370, 16),
9483 => conv_std_logic_vector(407, 16),
9484 => conv_std_logic_vector(444, 16),
9485 => conv_std_logic_vector(481, 16),
9486 => conv_std_logic_vector(518, 16),
9487 => conv_std_logic_vector(555, 16),
9488 => conv_std_logic_vector(592, 16),
9489 => conv_std_logic_vector(629, 16),
9490 => conv_std_logic_vector(666, 16),
9491 => conv_std_logic_vector(703, 16),
9492 => conv_std_logic_vector(740, 16),
9493 => conv_std_logic_vector(777, 16),
9494 => conv_std_logic_vector(814, 16),
9495 => conv_std_logic_vector(851, 16),
9496 => conv_std_logic_vector(888, 16),
9497 => conv_std_logic_vector(925, 16),
9498 => conv_std_logic_vector(962, 16),
9499 => conv_std_logic_vector(999, 16),
9500 => conv_std_logic_vector(1036, 16),
9501 => conv_std_logic_vector(1073, 16),
9502 => conv_std_logic_vector(1110, 16),
9503 => conv_std_logic_vector(1147, 16),
9504 => conv_std_logic_vector(1184, 16),
9505 => conv_std_logic_vector(1221, 16),
9506 => conv_std_logic_vector(1258, 16),
9507 => conv_std_logic_vector(1295, 16),
9508 => conv_std_logic_vector(1332, 16),
9509 => conv_std_logic_vector(1369, 16),
9510 => conv_std_logic_vector(1406, 16),
9511 => conv_std_logic_vector(1443, 16),
9512 => conv_std_logic_vector(1480, 16),
9513 => conv_std_logic_vector(1517, 16),
9514 => conv_std_logic_vector(1554, 16),
9515 => conv_std_logic_vector(1591, 16),
9516 => conv_std_logic_vector(1628, 16),
9517 => conv_std_logic_vector(1665, 16),
9518 => conv_std_logic_vector(1702, 16),
9519 => conv_std_logic_vector(1739, 16),
9520 => conv_std_logic_vector(1776, 16),
9521 => conv_std_logic_vector(1813, 16),
9522 => conv_std_logic_vector(1850, 16),
9523 => conv_std_logic_vector(1887, 16),
9524 => conv_std_logic_vector(1924, 16),
9525 => conv_std_logic_vector(1961, 16),
9526 => conv_std_logic_vector(1998, 16),
9527 => conv_std_logic_vector(2035, 16),
9528 => conv_std_logic_vector(2072, 16),
9529 => conv_std_logic_vector(2109, 16),
9530 => conv_std_logic_vector(2146, 16),
9531 => conv_std_logic_vector(2183, 16),
9532 => conv_std_logic_vector(2220, 16),
9533 => conv_std_logic_vector(2257, 16),
9534 => conv_std_logic_vector(2294, 16),
9535 => conv_std_logic_vector(2331, 16),
9536 => conv_std_logic_vector(2368, 16),
9537 => conv_std_logic_vector(2405, 16),
9538 => conv_std_logic_vector(2442, 16),
9539 => conv_std_logic_vector(2479, 16),
9540 => conv_std_logic_vector(2516, 16),
9541 => conv_std_logic_vector(2553, 16),
9542 => conv_std_logic_vector(2590, 16),
9543 => conv_std_logic_vector(2627, 16),
9544 => conv_std_logic_vector(2664, 16),
9545 => conv_std_logic_vector(2701, 16),
9546 => conv_std_logic_vector(2738, 16),
9547 => conv_std_logic_vector(2775, 16),
9548 => conv_std_logic_vector(2812, 16),
9549 => conv_std_logic_vector(2849, 16),
9550 => conv_std_logic_vector(2886, 16),
9551 => conv_std_logic_vector(2923, 16),
9552 => conv_std_logic_vector(2960, 16),
9553 => conv_std_logic_vector(2997, 16),
9554 => conv_std_logic_vector(3034, 16),
9555 => conv_std_logic_vector(3071, 16),
9556 => conv_std_logic_vector(3108, 16),
9557 => conv_std_logic_vector(3145, 16),
9558 => conv_std_logic_vector(3182, 16),
9559 => conv_std_logic_vector(3219, 16),
9560 => conv_std_logic_vector(3256, 16),
9561 => conv_std_logic_vector(3293, 16),
9562 => conv_std_logic_vector(3330, 16),
9563 => conv_std_logic_vector(3367, 16),
9564 => conv_std_logic_vector(3404, 16),
9565 => conv_std_logic_vector(3441, 16),
9566 => conv_std_logic_vector(3478, 16),
9567 => conv_std_logic_vector(3515, 16),
9568 => conv_std_logic_vector(3552, 16),
9569 => conv_std_logic_vector(3589, 16),
9570 => conv_std_logic_vector(3626, 16),
9571 => conv_std_logic_vector(3663, 16),
9572 => conv_std_logic_vector(3700, 16),
9573 => conv_std_logic_vector(3737, 16),
9574 => conv_std_logic_vector(3774, 16),
9575 => conv_std_logic_vector(3811, 16),
9576 => conv_std_logic_vector(3848, 16),
9577 => conv_std_logic_vector(3885, 16),
9578 => conv_std_logic_vector(3922, 16),
9579 => conv_std_logic_vector(3959, 16),
9580 => conv_std_logic_vector(3996, 16),
9581 => conv_std_logic_vector(4033, 16),
9582 => conv_std_logic_vector(4070, 16),
9583 => conv_std_logic_vector(4107, 16),
9584 => conv_std_logic_vector(4144, 16),
9585 => conv_std_logic_vector(4181, 16),
9586 => conv_std_logic_vector(4218, 16),
9587 => conv_std_logic_vector(4255, 16),
9588 => conv_std_logic_vector(4292, 16),
9589 => conv_std_logic_vector(4329, 16),
9590 => conv_std_logic_vector(4366, 16),
9591 => conv_std_logic_vector(4403, 16),
9592 => conv_std_logic_vector(4440, 16),
9593 => conv_std_logic_vector(4477, 16),
9594 => conv_std_logic_vector(4514, 16),
9595 => conv_std_logic_vector(4551, 16),
9596 => conv_std_logic_vector(4588, 16),
9597 => conv_std_logic_vector(4625, 16),
9598 => conv_std_logic_vector(4662, 16),
9599 => conv_std_logic_vector(4699, 16),
9600 => conv_std_logic_vector(4736, 16),
9601 => conv_std_logic_vector(4773, 16),
9602 => conv_std_logic_vector(4810, 16),
9603 => conv_std_logic_vector(4847, 16),
9604 => conv_std_logic_vector(4884, 16),
9605 => conv_std_logic_vector(4921, 16),
9606 => conv_std_logic_vector(4958, 16),
9607 => conv_std_logic_vector(4995, 16),
9608 => conv_std_logic_vector(5032, 16),
9609 => conv_std_logic_vector(5069, 16),
9610 => conv_std_logic_vector(5106, 16),
9611 => conv_std_logic_vector(5143, 16),
9612 => conv_std_logic_vector(5180, 16),
9613 => conv_std_logic_vector(5217, 16),
9614 => conv_std_logic_vector(5254, 16),
9615 => conv_std_logic_vector(5291, 16),
9616 => conv_std_logic_vector(5328, 16),
9617 => conv_std_logic_vector(5365, 16),
9618 => conv_std_logic_vector(5402, 16),
9619 => conv_std_logic_vector(5439, 16),
9620 => conv_std_logic_vector(5476, 16),
9621 => conv_std_logic_vector(5513, 16),
9622 => conv_std_logic_vector(5550, 16),
9623 => conv_std_logic_vector(5587, 16),
9624 => conv_std_logic_vector(5624, 16),
9625 => conv_std_logic_vector(5661, 16),
9626 => conv_std_logic_vector(5698, 16),
9627 => conv_std_logic_vector(5735, 16),
9628 => conv_std_logic_vector(5772, 16),
9629 => conv_std_logic_vector(5809, 16),
9630 => conv_std_logic_vector(5846, 16),
9631 => conv_std_logic_vector(5883, 16),
9632 => conv_std_logic_vector(5920, 16),
9633 => conv_std_logic_vector(5957, 16),
9634 => conv_std_logic_vector(5994, 16),
9635 => conv_std_logic_vector(6031, 16),
9636 => conv_std_logic_vector(6068, 16),
9637 => conv_std_logic_vector(6105, 16),
9638 => conv_std_logic_vector(6142, 16),
9639 => conv_std_logic_vector(6179, 16),
9640 => conv_std_logic_vector(6216, 16),
9641 => conv_std_logic_vector(6253, 16),
9642 => conv_std_logic_vector(6290, 16),
9643 => conv_std_logic_vector(6327, 16),
9644 => conv_std_logic_vector(6364, 16),
9645 => conv_std_logic_vector(6401, 16),
9646 => conv_std_logic_vector(6438, 16),
9647 => conv_std_logic_vector(6475, 16),
9648 => conv_std_logic_vector(6512, 16),
9649 => conv_std_logic_vector(6549, 16),
9650 => conv_std_logic_vector(6586, 16),
9651 => conv_std_logic_vector(6623, 16),
9652 => conv_std_logic_vector(6660, 16),
9653 => conv_std_logic_vector(6697, 16),
9654 => conv_std_logic_vector(6734, 16),
9655 => conv_std_logic_vector(6771, 16),
9656 => conv_std_logic_vector(6808, 16),
9657 => conv_std_logic_vector(6845, 16),
9658 => conv_std_logic_vector(6882, 16),
9659 => conv_std_logic_vector(6919, 16),
9660 => conv_std_logic_vector(6956, 16),
9661 => conv_std_logic_vector(6993, 16),
9662 => conv_std_logic_vector(7030, 16),
9663 => conv_std_logic_vector(7067, 16),
9664 => conv_std_logic_vector(7104, 16),
9665 => conv_std_logic_vector(7141, 16),
9666 => conv_std_logic_vector(7178, 16),
9667 => conv_std_logic_vector(7215, 16),
9668 => conv_std_logic_vector(7252, 16),
9669 => conv_std_logic_vector(7289, 16),
9670 => conv_std_logic_vector(7326, 16),
9671 => conv_std_logic_vector(7363, 16),
9672 => conv_std_logic_vector(7400, 16),
9673 => conv_std_logic_vector(7437, 16),
9674 => conv_std_logic_vector(7474, 16),
9675 => conv_std_logic_vector(7511, 16),
9676 => conv_std_logic_vector(7548, 16),
9677 => conv_std_logic_vector(7585, 16),
9678 => conv_std_logic_vector(7622, 16),
9679 => conv_std_logic_vector(7659, 16),
9680 => conv_std_logic_vector(7696, 16),
9681 => conv_std_logic_vector(7733, 16),
9682 => conv_std_logic_vector(7770, 16),
9683 => conv_std_logic_vector(7807, 16),
9684 => conv_std_logic_vector(7844, 16),
9685 => conv_std_logic_vector(7881, 16),
9686 => conv_std_logic_vector(7918, 16),
9687 => conv_std_logic_vector(7955, 16),
9688 => conv_std_logic_vector(7992, 16),
9689 => conv_std_logic_vector(8029, 16),
9690 => conv_std_logic_vector(8066, 16),
9691 => conv_std_logic_vector(8103, 16),
9692 => conv_std_logic_vector(8140, 16),
9693 => conv_std_logic_vector(8177, 16),
9694 => conv_std_logic_vector(8214, 16),
9695 => conv_std_logic_vector(8251, 16),
9696 => conv_std_logic_vector(8288, 16),
9697 => conv_std_logic_vector(8325, 16),
9698 => conv_std_logic_vector(8362, 16),
9699 => conv_std_logic_vector(8399, 16),
9700 => conv_std_logic_vector(8436, 16),
9701 => conv_std_logic_vector(8473, 16),
9702 => conv_std_logic_vector(8510, 16),
9703 => conv_std_logic_vector(8547, 16),
9704 => conv_std_logic_vector(8584, 16),
9705 => conv_std_logic_vector(8621, 16),
9706 => conv_std_logic_vector(8658, 16),
9707 => conv_std_logic_vector(8695, 16),
9708 => conv_std_logic_vector(8732, 16),
9709 => conv_std_logic_vector(8769, 16),
9710 => conv_std_logic_vector(8806, 16),
9711 => conv_std_logic_vector(8843, 16),
9712 => conv_std_logic_vector(8880, 16),
9713 => conv_std_logic_vector(8917, 16),
9714 => conv_std_logic_vector(8954, 16),
9715 => conv_std_logic_vector(8991, 16),
9716 => conv_std_logic_vector(9028, 16),
9717 => conv_std_logic_vector(9065, 16),
9718 => conv_std_logic_vector(9102, 16),
9719 => conv_std_logic_vector(9139, 16),
9720 => conv_std_logic_vector(9176, 16),
9721 => conv_std_logic_vector(9213, 16),
9722 => conv_std_logic_vector(9250, 16),
9723 => conv_std_logic_vector(9287, 16),
9724 => conv_std_logic_vector(9324, 16),
9725 => conv_std_logic_vector(9361, 16),
9726 => conv_std_logic_vector(9398, 16),
9727 => conv_std_logic_vector(9435, 16),
9728 => conv_std_logic_vector(0, 16),
9729 => conv_std_logic_vector(38, 16),
9730 => conv_std_logic_vector(76, 16),
9731 => conv_std_logic_vector(114, 16),
9732 => conv_std_logic_vector(152, 16),
9733 => conv_std_logic_vector(190, 16),
9734 => conv_std_logic_vector(228, 16),
9735 => conv_std_logic_vector(266, 16),
9736 => conv_std_logic_vector(304, 16),
9737 => conv_std_logic_vector(342, 16),
9738 => conv_std_logic_vector(380, 16),
9739 => conv_std_logic_vector(418, 16),
9740 => conv_std_logic_vector(456, 16),
9741 => conv_std_logic_vector(494, 16),
9742 => conv_std_logic_vector(532, 16),
9743 => conv_std_logic_vector(570, 16),
9744 => conv_std_logic_vector(608, 16),
9745 => conv_std_logic_vector(646, 16),
9746 => conv_std_logic_vector(684, 16),
9747 => conv_std_logic_vector(722, 16),
9748 => conv_std_logic_vector(760, 16),
9749 => conv_std_logic_vector(798, 16),
9750 => conv_std_logic_vector(836, 16),
9751 => conv_std_logic_vector(874, 16),
9752 => conv_std_logic_vector(912, 16),
9753 => conv_std_logic_vector(950, 16),
9754 => conv_std_logic_vector(988, 16),
9755 => conv_std_logic_vector(1026, 16),
9756 => conv_std_logic_vector(1064, 16),
9757 => conv_std_logic_vector(1102, 16),
9758 => conv_std_logic_vector(1140, 16),
9759 => conv_std_logic_vector(1178, 16),
9760 => conv_std_logic_vector(1216, 16),
9761 => conv_std_logic_vector(1254, 16),
9762 => conv_std_logic_vector(1292, 16),
9763 => conv_std_logic_vector(1330, 16),
9764 => conv_std_logic_vector(1368, 16),
9765 => conv_std_logic_vector(1406, 16),
9766 => conv_std_logic_vector(1444, 16),
9767 => conv_std_logic_vector(1482, 16),
9768 => conv_std_logic_vector(1520, 16),
9769 => conv_std_logic_vector(1558, 16),
9770 => conv_std_logic_vector(1596, 16),
9771 => conv_std_logic_vector(1634, 16),
9772 => conv_std_logic_vector(1672, 16),
9773 => conv_std_logic_vector(1710, 16),
9774 => conv_std_logic_vector(1748, 16),
9775 => conv_std_logic_vector(1786, 16),
9776 => conv_std_logic_vector(1824, 16),
9777 => conv_std_logic_vector(1862, 16),
9778 => conv_std_logic_vector(1900, 16),
9779 => conv_std_logic_vector(1938, 16),
9780 => conv_std_logic_vector(1976, 16),
9781 => conv_std_logic_vector(2014, 16),
9782 => conv_std_logic_vector(2052, 16),
9783 => conv_std_logic_vector(2090, 16),
9784 => conv_std_logic_vector(2128, 16),
9785 => conv_std_logic_vector(2166, 16),
9786 => conv_std_logic_vector(2204, 16),
9787 => conv_std_logic_vector(2242, 16),
9788 => conv_std_logic_vector(2280, 16),
9789 => conv_std_logic_vector(2318, 16),
9790 => conv_std_logic_vector(2356, 16),
9791 => conv_std_logic_vector(2394, 16),
9792 => conv_std_logic_vector(2432, 16),
9793 => conv_std_logic_vector(2470, 16),
9794 => conv_std_logic_vector(2508, 16),
9795 => conv_std_logic_vector(2546, 16),
9796 => conv_std_logic_vector(2584, 16),
9797 => conv_std_logic_vector(2622, 16),
9798 => conv_std_logic_vector(2660, 16),
9799 => conv_std_logic_vector(2698, 16),
9800 => conv_std_logic_vector(2736, 16),
9801 => conv_std_logic_vector(2774, 16),
9802 => conv_std_logic_vector(2812, 16),
9803 => conv_std_logic_vector(2850, 16),
9804 => conv_std_logic_vector(2888, 16),
9805 => conv_std_logic_vector(2926, 16),
9806 => conv_std_logic_vector(2964, 16),
9807 => conv_std_logic_vector(3002, 16),
9808 => conv_std_logic_vector(3040, 16),
9809 => conv_std_logic_vector(3078, 16),
9810 => conv_std_logic_vector(3116, 16),
9811 => conv_std_logic_vector(3154, 16),
9812 => conv_std_logic_vector(3192, 16),
9813 => conv_std_logic_vector(3230, 16),
9814 => conv_std_logic_vector(3268, 16),
9815 => conv_std_logic_vector(3306, 16),
9816 => conv_std_logic_vector(3344, 16),
9817 => conv_std_logic_vector(3382, 16),
9818 => conv_std_logic_vector(3420, 16),
9819 => conv_std_logic_vector(3458, 16),
9820 => conv_std_logic_vector(3496, 16),
9821 => conv_std_logic_vector(3534, 16),
9822 => conv_std_logic_vector(3572, 16),
9823 => conv_std_logic_vector(3610, 16),
9824 => conv_std_logic_vector(3648, 16),
9825 => conv_std_logic_vector(3686, 16),
9826 => conv_std_logic_vector(3724, 16),
9827 => conv_std_logic_vector(3762, 16),
9828 => conv_std_logic_vector(3800, 16),
9829 => conv_std_logic_vector(3838, 16),
9830 => conv_std_logic_vector(3876, 16),
9831 => conv_std_logic_vector(3914, 16),
9832 => conv_std_logic_vector(3952, 16),
9833 => conv_std_logic_vector(3990, 16),
9834 => conv_std_logic_vector(4028, 16),
9835 => conv_std_logic_vector(4066, 16),
9836 => conv_std_logic_vector(4104, 16),
9837 => conv_std_logic_vector(4142, 16),
9838 => conv_std_logic_vector(4180, 16),
9839 => conv_std_logic_vector(4218, 16),
9840 => conv_std_logic_vector(4256, 16),
9841 => conv_std_logic_vector(4294, 16),
9842 => conv_std_logic_vector(4332, 16),
9843 => conv_std_logic_vector(4370, 16),
9844 => conv_std_logic_vector(4408, 16),
9845 => conv_std_logic_vector(4446, 16),
9846 => conv_std_logic_vector(4484, 16),
9847 => conv_std_logic_vector(4522, 16),
9848 => conv_std_logic_vector(4560, 16),
9849 => conv_std_logic_vector(4598, 16),
9850 => conv_std_logic_vector(4636, 16),
9851 => conv_std_logic_vector(4674, 16),
9852 => conv_std_logic_vector(4712, 16),
9853 => conv_std_logic_vector(4750, 16),
9854 => conv_std_logic_vector(4788, 16),
9855 => conv_std_logic_vector(4826, 16),
9856 => conv_std_logic_vector(4864, 16),
9857 => conv_std_logic_vector(4902, 16),
9858 => conv_std_logic_vector(4940, 16),
9859 => conv_std_logic_vector(4978, 16),
9860 => conv_std_logic_vector(5016, 16),
9861 => conv_std_logic_vector(5054, 16),
9862 => conv_std_logic_vector(5092, 16),
9863 => conv_std_logic_vector(5130, 16),
9864 => conv_std_logic_vector(5168, 16),
9865 => conv_std_logic_vector(5206, 16),
9866 => conv_std_logic_vector(5244, 16),
9867 => conv_std_logic_vector(5282, 16),
9868 => conv_std_logic_vector(5320, 16),
9869 => conv_std_logic_vector(5358, 16),
9870 => conv_std_logic_vector(5396, 16),
9871 => conv_std_logic_vector(5434, 16),
9872 => conv_std_logic_vector(5472, 16),
9873 => conv_std_logic_vector(5510, 16),
9874 => conv_std_logic_vector(5548, 16),
9875 => conv_std_logic_vector(5586, 16),
9876 => conv_std_logic_vector(5624, 16),
9877 => conv_std_logic_vector(5662, 16),
9878 => conv_std_logic_vector(5700, 16),
9879 => conv_std_logic_vector(5738, 16),
9880 => conv_std_logic_vector(5776, 16),
9881 => conv_std_logic_vector(5814, 16),
9882 => conv_std_logic_vector(5852, 16),
9883 => conv_std_logic_vector(5890, 16),
9884 => conv_std_logic_vector(5928, 16),
9885 => conv_std_logic_vector(5966, 16),
9886 => conv_std_logic_vector(6004, 16),
9887 => conv_std_logic_vector(6042, 16),
9888 => conv_std_logic_vector(6080, 16),
9889 => conv_std_logic_vector(6118, 16),
9890 => conv_std_logic_vector(6156, 16),
9891 => conv_std_logic_vector(6194, 16),
9892 => conv_std_logic_vector(6232, 16),
9893 => conv_std_logic_vector(6270, 16),
9894 => conv_std_logic_vector(6308, 16),
9895 => conv_std_logic_vector(6346, 16),
9896 => conv_std_logic_vector(6384, 16),
9897 => conv_std_logic_vector(6422, 16),
9898 => conv_std_logic_vector(6460, 16),
9899 => conv_std_logic_vector(6498, 16),
9900 => conv_std_logic_vector(6536, 16),
9901 => conv_std_logic_vector(6574, 16),
9902 => conv_std_logic_vector(6612, 16),
9903 => conv_std_logic_vector(6650, 16),
9904 => conv_std_logic_vector(6688, 16),
9905 => conv_std_logic_vector(6726, 16),
9906 => conv_std_logic_vector(6764, 16),
9907 => conv_std_logic_vector(6802, 16),
9908 => conv_std_logic_vector(6840, 16),
9909 => conv_std_logic_vector(6878, 16),
9910 => conv_std_logic_vector(6916, 16),
9911 => conv_std_logic_vector(6954, 16),
9912 => conv_std_logic_vector(6992, 16),
9913 => conv_std_logic_vector(7030, 16),
9914 => conv_std_logic_vector(7068, 16),
9915 => conv_std_logic_vector(7106, 16),
9916 => conv_std_logic_vector(7144, 16),
9917 => conv_std_logic_vector(7182, 16),
9918 => conv_std_logic_vector(7220, 16),
9919 => conv_std_logic_vector(7258, 16),
9920 => conv_std_logic_vector(7296, 16),
9921 => conv_std_logic_vector(7334, 16),
9922 => conv_std_logic_vector(7372, 16),
9923 => conv_std_logic_vector(7410, 16),
9924 => conv_std_logic_vector(7448, 16),
9925 => conv_std_logic_vector(7486, 16),
9926 => conv_std_logic_vector(7524, 16),
9927 => conv_std_logic_vector(7562, 16),
9928 => conv_std_logic_vector(7600, 16),
9929 => conv_std_logic_vector(7638, 16),
9930 => conv_std_logic_vector(7676, 16),
9931 => conv_std_logic_vector(7714, 16),
9932 => conv_std_logic_vector(7752, 16),
9933 => conv_std_logic_vector(7790, 16),
9934 => conv_std_logic_vector(7828, 16),
9935 => conv_std_logic_vector(7866, 16),
9936 => conv_std_logic_vector(7904, 16),
9937 => conv_std_logic_vector(7942, 16),
9938 => conv_std_logic_vector(7980, 16),
9939 => conv_std_logic_vector(8018, 16),
9940 => conv_std_logic_vector(8056, 16),
9941 => conv_std_logic_vector(8094, 16),
9942 => conv_std_logic_vector(8132, 16),
9943 => conv_std_logic_vector(8170, 16),
9944 => conv_std_logic_vector(8208, 16),
9945 => conv_std_logic_vector(8246, 16),
9946 => conv_std_logic_vector(8284, 16),
9947 => conv_std_logic_vector(8322, 16),
9948 => conv_std_logic_vector(8360, 16),
9949 => conv_std_logic_vector(8398, 16),
9950 => conv_std_logic_vector(8436, 16),
9951 => conv_std_logic_vector(8474, 16),
9952 => conv_std_logic_vector(8512, 16),
9953 => conv_std_logic_vector(8550, 16),
9954 => conv_std_logic_vector(8588, 16),
9955 => conv_std_logic_vector(8626, 16),
9956 => conv_std_logic_vector(8664, 16),
9957 => conv_std_logic_vector(8702, 16),
9958 => conv_std_logic_vector(8740, 16),
9959 => conv_std_logic_vector(8778, 16),
9960 => conv_std_logic_vector(8816, 16),
9961 => conv_std_logic_vector(8854, 16),
9962 => conv_std_logic_vector(8892, 16),
9963 => conv_std_logic_vector(8930, 16),
9964 => conv_std_logic_vector(8968, 16),
9965 => conv_std_logic_vector(9006, 16),
9966 => conv_std_logic_vector(9044, 16),
9967 => conv_std_logic_vector(9082, 16),
9968 => conv_std_logic_vector(9120, 16),
9969 => conv_std_logic_vector(9158, 16),
9970 => conv_std_logic_vector(9196, 16),
9971 => conv_std_logic_vector(9234, 16),
9972 => conv_std_logic_vector(9272, 16),
9973 => conv_std_logic_vector(9310, 16),
9974 => conv_std_logic_vector(9348, 16),
9975 => conv_std_logic_vector(9386, 16),
9976 => conv_std_logic_vector(9424, 16),
9977 => conv_std_logic_vector(9462, 16),
9978 => conv_std_logic_vector(9500, 16),
9979 => conv_std_logic_vector(9538, 16),
9980 => conv_std_logic_vector(9576, 16),
9981 => conv_std_logic_vector(9614, 16),
9982 => conv_std_logic_vector(9652, 16),
9983 => conv_std_logic_vector(9690, 16),
9984 => conv_std_logic_vector(0, 16),
9985 => conv_std_logic_vector(39, 16),
9986 => conv_std_logic_vector(78, 16),
9987 => conv_std_logic_vector(117, 16),
9988 => conv_std_logic_vector(156, 16),
9989 => conv_std_logic_vector(195, 16),
9990 => conv_std_logic_vector(234, 16),
9991 => conv_std_logic_vector(273, 16),
9992 => conv_std_logic_vector(312, 16),
9993 => conv_std_logic_vector(351, 16),
9994 => conv_std_logic_vector(390, 16),
9995 => conv_std_logic_vector(429, 16),
9996 => conv_std_logic_vector(468, 16),
9997 => conv_std_logic_vector(507, 16),
9998 => conv_std_logic_vector(546, 16),
9999 => conv_std_logic_vector(585, 16),
10000 => conv_std_logic_vector(624, 16),
10001 => conv_std_logic_vector(663, 16),
10002 => conv_std_logic_vector(702, 16),
10003 => conv_std_logic_vector(741, 16),
10004 => conv_std_logic_vector(780, 16),
10005 => conv_std_logic_vector(819, 16),
10006 => conv_std_logic_vector(858, 16),
10007 => conv_std_logic_vector(897, 16),
10008 => conv_std_logic_vector(936, 16),
10009 => conv_std_logic_vector(975, 16),
10010 => conv_std_logic_vector(1014, 16),
10011 => conv_std_logic_vector(1053, 16),
10012 => conv_std_logic_vector(1092, 16),
10013 => conv_std_logic_vector(1131, 16),
10014 => conv_std_logic_vector(1170, 16),
10015 => conv_std_logic_vector(1209, 16),
10016 => conv_std_logic_vector(1248, 16),
10017 => conv_std_logic_vector(1287, 16),
10018 => conv_std_logic_vector(1326, 16),
10019 => conv_std_logic_vector(1365, 16),
10020 => conv_std_logic_vector(1404, 16),
10021 => conv_std_logic_vector(1443, 16),
10022 => conv_std_logic_vector(1482, 16),
10023 => conv_std_logic_vector(1521, 16),
10024 => conv_std_logic_vector(1560, 16),
10025 => conv_std_logic_vector(1599, 16),
10026 => conv_std_logic_vector(1638, 16),
10027 => conv_std_logic_vector(1677, 16),
10028 => conv_std_logic_vector(1716, 16),
10029 => conv_std_logic_vector(1755, 16),
10030 => conv_std_logic_vector(1794, 16),
10031 => conv_std_logic_vector(1833, 16),
10032 => conv_std_logic_vector(1872, 16),
10033 => conv_std_logic_vector(1911, 16),
10034 => conv_std_logic_vector(1950, 16),
10035 => conv_std_logic_vector(1989, 16),
10036 => conv_std_logic_vector(2028, 16),
10037 => conv_std_logic_vector(2067, 16),
10038 => conv_std_logic_vector(2106, 16),
10039 => conv_std_logic_vector(2145, 16),
10040 => conv_std_logic_vector(2184, 16),
10041 => conv_std_logic_vector(2223, 16),
10042 => conv_std_logic_vector(2262, 16),
10043 => conv_std_logic_vector(2301, 16),
10044 => conv_std_logic_vector(2340, 16),
10045 => conv_std_logic_vector(2379, 16),
10046 => conv_std_logic_vector(2418, 16),
10047 => conv_std_logic_vector(2457, 16),
10048 => conv_std_logic_vector(2496, 16),
10049 => conv_std_logic_vector(2535, 16),
10050 => conv_std_logic_vector(2574, 16),
10051 => conv_std_logic_vector(2613, 16),
10052 => conv_std_logic_vector(2652, 16),
10053 => conv_std_logic_vector(2691, 16),
10054 => conv_std_logic_vector(2730, 16),
10055 => conv_std_logic_vector(2769, 16),
10056 => conv_std_logic_vector(2808, 16),
10057 => conv_std_logic_vector(2847, 16),
10058 => conv_std_logic_vector(2886, 16),
10059 => conv_std_logic_vector(2925, 16),
10060 => conv_std_logic_vector(2964, 16),
10061 => conv_std_logic_vector(3003, 16),
10062 => conv_std_logic_vector(3042, 16),
10063 => conv_std_logic_vector(3081, 16),
10064 => conv_std_logic_vector(3120, 16),
10065 => conv_std_logic_vector(3159, 16),
10066 => conv_std_logic_vector(3198, 16),
10067 => conv_std_logic_vector(3237, 16),
10068 => conv_std_logic_vector(3276, 16),
10069 => conv_std_logic_vector(3315, 16),
10070 => conv_std_logic_vector(3354, 16),
10071 => conv_std_logic_vector(3393, 16),
10072 => conv_std_logic_vector(3432, 16),
10073 => conv_std_logic_vector(3471, 16),
10074 => conv_std_logic_vector(3510, 16),
10075 => conv_std_logic_vector(3549, 16),
10076 => conv_std_logic_vector(3588, 16),
10077 => conv_std_logic_vector(3627, 16),
10078 => conv_std_logic_vector(3666, 16),
10079 => conv_std_logic_vector(3705, 16),
10080 => conv_std_logic_vector(3744, 16),
10081 => conv_std_logic_vector(3783, 16),
10082 => conv_std_logic_vector(3822, 16),
10083 => conv_std_logic_vector(3861, 16),
10084 => conv_std_logic_vector(3900, 16),
10085 => conv_std_logic_vector(3939, 16),
10086 => conv_std_logic_vector(3978, 16),
10087 => conv_std_logic_vector(4017, 16),
10088 => conv_std_logic_vector(4056, 16),
10089 => conv_std_logic_vector(4095, 16),
10090 => conv_std_logic_vector(4134, 16),
10091 => conv_std_logic_vector(4173, 16),
10092 => conv_std_logic_vector(4212, 16),
10093 => conv_std_logic_vector(4251, 16),
10094 => conv_std_logic_vector(4290, 16),
10095 => conv_std_logic_vector(4329, 16),
10096 => conv_std_logic_vector(4368, 16),
10097 => conv_std_logic_vector(4407, 16),
10098 => conv_std_logic_vector(4446, 16),
10099 => conv_std_logic_vector(4485, 16),
10100 => conv_std_logic_vector(4524, 16),
10101 => conv_std_logic_vector(4563, 16),
10102 => conv_std_logic_vector(4602, 16),
10103 => conv_std_logic_vector(4641, 16),
10104 => conv_std_logic_vector(4680, 16),
10105 => conv_std_logic_vector(4719, 16),
10106 => conv_std_logic_vector(4758, 16),
10107 => conv_std_logic_vector(4797, 16),
10108 => conv_std_logic_vector(4836, 16),
10109 => conv_std_logic_vector(4875, 16),
10110 => conv_std_logic_vector(4914, 16),
10111 => conv_std_logic_vector(4953, 16),
10112 => conv_std_logic_vector(4992, 16),
10113 => conv_std_logic_vector(5031, 16),
10114 => conv_std_logic_vector(5070, 16),
10115 => conv_std_logic_vector(5109, 16),
10116 => conv_std_logic_vector(5148, 16),
10117 => conv_std_logic_vector(5187, 16),
10118 => conv_std_logic_vector(5226, 16),
10119 => conv_std_logic_vector(5265, 16),
10120 => conv_std_logic_vector(5304, 16),
10121 => conv_std_logic_vector(5343, 16),
10122 => conv_std_logic_vector(5382, 16),
10123 => conv_std_logic_vector(5421, 16),
10124 => conv_std_logic_vector(5460, 16),
10125 => conv_std_logic_vector(5499, 16),
10126 => conv_std_logic_vector(5538, 16),
10127 => conv_std_logic_vector(5577, 16),
10128 => conv_std_logic_vector(5616, 16),
10129 => conv_std_logic_vector(5655, 16),
10130 => conv_std_logic_vector(5694, 16),
10131 => conv_std_logic_vector(5733, 16),
10132 => conv_std_logic_vector(5772, 16),
10133 => conv_std_logic_vector(5811, 16),
10134 => conv_std_logic_vector(5850, 16),
10135 => conv_std_logic_vector(5889, 16),
10136 => conv_std_logic_vector(5928, 16),
10137 => conv_std_logic_vector(5967, 16),
10138 => conv_std_logic_vector(6006, 16),
10139 => conv_std_logic_vector(6045, 16),
10140 => conv_std_logic_vector(6084, 16),
10141 => conv_std_logic_vector(6123, 16),
10142 => conv_std_logic_vector(6162, 16),
10143 => conv_std_logic_vector(6201, 16),
10144 => conv_std_logic_vector(6240, 16),
10145 => conv_std_logic_vector(6279, 16),
10146 => conv_std_logic_vector(6318, 16),
10147 => conv_std_logic_vector(6357, 16),
10148 => conv_std_logic_vector(6396, 16),
10149 => conv_std_logic_vector(6435, 16),
10150 => conv_std_logic_vector(6474, 16),
10151 => conv_std_logic_vector(6513, 16),
10152 => conv_std_logic_vector(6552, 16),
10153 => conv_std_logic_vector(6591, 16),
10154 => conv_std_logic_vector(6630, 16),
10155 => conv_std_logic_vector(6669, 16),
10156 => conv_std_logic_vector(6708, 16),
10157 => conv_std_logic_vector(6747, 16),
10158 => conv_std_logic_vector(6786, 16),
10159 => conv_std_logic_vector(6825, 16),
10160 => conv_std_logic_vector(6864, 16),
10161 => conv_std_logic_vector(6903, 16),
10162 => conv_std_logic_vector(6942, 16),
10163 => conv_std_logic_vector(6981, 16),
10164 => conv_std_logic_vector(7020, 16),
10165 => conv_std_logic_vector(7059, 16),
10166 => conv_std_logic_vector(7098, 16),
10167 => conv_std_logic_vector(7137, 16),
10168 => conv_std_logic_vector(7176, 16),
10169 => conv_std_logic_vector(7215, 16),
10170 => conv_std_logic_vector(7254, 16),
10171 => conv_std_logic_vector(7293, 16),
10172 => conv_std_logic_vector(7332, 16),
10173 => conv_std_logic_vector(7371, 16),
10174 => conv_std_logic_vector(7410, 16),
10175 => conv_std_logic_vector(7449, 16),
10176 => conv_std_logic_vector(7488, 16),
10177 => conv_std_logic_vector(7527, 16),
10178 => conv_std_logic_vector(7566, 16),
10179 => conv_std_logic_vector(7605, 16),
10180 => conv_std_logic_vector(7644, 16),
10181 => conv_std_logic_vector(7683, 16),
10182 => conv_std_logic_vector(7722, 16),
10183 => conv_std_logic_vector(7761, 16),
10184 => conv_std_logic_vector(7800, 16),
10185 => conv_std_logic_vector(7839, 16),
10186 => conv_std_logic_vector(7878, 16),
10187 => conv_std_logic_vector(7917, 16),
10188 => conv_std_logic_vector(7956, 16),
10189 => conv_std_logic_vector(7995, 16),
10190 => conv_std_logic_vector(8034, 16),
10191 => conv_std_logic_vector(8073, 16),
10192 => conv_std_logic_vector(8112, 16),
10193 => conv_std_logic_vector(8151, 16),
10194 => conv_std_logic_vector(8190, 16),
10195 => conv_std_logic_vector(8229, 16),
10196 => conv_std_logic_vector(8268, 16),
10197 => conv_std_logic_vector(8307, 16),
10198 => conv_std_logic_vector(8346, 16),
10199 => conv_std_logic_vector(8385, 16),
10200 => conv_std_logic_vector(8424, 16),
10201 => conv_std_logic_vector(8463, 16),
10202 => conv_std_logic_vector(8502, 16),
10203 => conv_std_logic_vector(8541, 16),
10204 => conv_std_logic_vector(8580, 16),
10205 => conv_std_logic_vector(8619, 16),
10206 => conv_std_logic_vector(8658, 16),
10207 => conv_std_logic_vector(8697, 16),
10208 => conv_std_logic_vector(8736, 16),
10209 => conv_std_logic_vector(8775, 16),
10210 => conv_std_logic_vector(8814, 16),
10211 => conv_std_logic_vector(8853, 16),
10212 => conv_std_logic_vector(8892, 16),
10213 => conv_std_logic_vector(8931, 16),
10214 => conv_std_logic_vector(8970, 16),
10215 => conv_std_logic_vector(9009, 16),
10216 => conv_std_logic_vector(9048, 16),
10217 => conv_std_logic_vector(9087, 16),
10218 => conv_std_logic_vector(9126, 16),
10219 => conv_std_logic_vector(9165, 16),
10220 => conv_std_logic_vector(9204, 16),
10221 => conv_std_logic_vector(9243, 16),
10222 => conv_std_logic_vector(9282, 16),
10223 => conv_std_logic_vector(9321, 16),
10224 => conv_std_logic_vector(9360, 16),
10225 => conv_std_logic_vector(9399, 16),
10226 => conv_std_logic_vector(9438, 16),
10227 => conv_std_logic_vector(9477, 16),
10228 => conv_std_logic_vector(9516, 16),
10229 => conv_std_logic_vector(9555, 16),
10230 => conv_std_logic_vector(9594, 16),
10231 => conv_std_logic_vector(9633, 16),
10232 => conv_std_logic_vector(9672, 16),
10233 => conv_std_logic_vector(9711, 16),
10234 => conv_std_logic_vector(9750, 16),
10235 => conv_std_logic_vector(9789, 16),
10236 => conv_std_logic_vector(9828, 16),
10237 => conv_std_logic_vector(9867, 16),
10238 => conv_std_logic_vector(9906, 16),
10239 => conv_std_logic_vector(9945, 16),
10240 => conv_std_logic_vector(0, 16),
10241 => conv_std_logic_vector(40, 16),
10242 => conv_std_logic_vector(80, 16),
10243 => conv_std_logic_vector(120, 16),
10244 => conv_std_logic_vector(160, 16),
10245 => conv_std_logic_vector(200, 16),
10246 => conv_std_logic_vector(240, 16),
10247 => conv_std_logic_vector(280, 16),
10248 => conv_std_logic_vector(320, 16),
10249 => conv_std_logic_vector(360, 16),
10250 => conv_std_logic_vector(400, 16),
10251 => conv_std_logic_vector(440, 16),
10252 => conv_std_logic_vector(480, 16),
10253 => conv_std_logic_vector(520, 16),
10254 => conv_std_logic_vector(560, 16),
10255 => conv_std_logic_vector(600, 16),
10256 => conv_std_logic_vector(640, 16),
10257 => conv_std_logic_vector(680, 16),
10258 => conv_std_logic_vector(720, 16),
10259 => conv_std_logic_vector(760, 16),
10260 => conv_std_logic_vector(800, 16),
10261 => conv_std_logic_vector(840, 16),
10262 => conv_std_logic_vector(880, 16),
10263 => conv_std_logic_vector(920, 16),
10264 => conv_std_logic_vector(960, 16),
10265 => conv_std_logic_vector(1000, 16),
10266 => conv_std_logic_vector(1040, 16),
10267 => conv_std_logic_vector(1080, 16),
10268 => conv_std_logic_vector(1120, 16),
10269 => conv_std_logic_vector(1160, 16),
10270 => conv_std_logic_vector(1200, 16),
10271 => conv_std_logic_vector(1240, 16),
10272 => conv_std_logic_vector(1280, 16),
10273 => conv_std_logic_vector(1320, 16),
10274 => conv_std_logic_vector(1360, 16),
10275 => conv_std_logic_vector(1400, 16),
10276 => conv_std_logic_vector(1440, 16),
10277 => conv_std_logic_vector(1480, 16),
10278 => conv_std_logic_vector(1520, 16),
10279 => conv_std_logic_vector(1560, 16),
10280 => conv_std_logic_vector(1600, 16),
10281 => conv_std_logic_vector(1640, 16),
10282 => conv_std_logic_vector(1680, 16),
10283 => conv_std_logic_vector(1720, 16),
10284 => conv_std_logic_vector(1760, 16),
10285 => conv_std_logic_vector(1800, 16),
10286 => conv_std_logic_vector(1840, 16),
10287 => conv_std_logic_vector(1880, 16),
10288 => conv_std_logic_vector(1920, 16),
10289 => conv_std_logic_vector(1960, 16),
10290 => conv_std_logic_vector(2000, 16),
10291 => conv_std_logic_vector(2040, 16),
10292 => conv_std_logic_vector(2080, 16),
10293 => conv_std_logic_vector(2120, 16),
10294 => conv_std_logic_vector(2160, 16),
10295 => conv_std_logic_vector(2200, 16),
10296 => conv_std_logic_vector(2240, 16),
10297 => conv_std_logic_vector(2280, 16),
10298 => conv_std_logic_vector(2320, 16),
10299 => conv_std_logic_vector(2360, 16),
10300 => conv_std_logic_vector(2400, 16),
10301 => conv_std_logic_vector(2440, 16),
10302 => conv_std_logic_vector(2480, 16),
10303 => conv_std_logic_vector(2520, 16),
10304 => conv_std_logic_vector(2560, 16),
10305 => conv_std_logic_vector(2600, 16),
10306 => conv_std_logic_vector(2640, 16),
10307 => conv_std_logic_vector(2680, 16),
10308 => conv_std_logic_vector(2720, 16),
10309 => conv_std_logic_vector(2760, 16),
10310 => conv_std_logic_vector(2800, 16),
10311 => conv_std_logic_vector(2840, 16),
10312 => conv_std_logic_vector(2880, 16),
10313 => conv_std_logic_vector(2920, 16),
10314 => conv_std_logic_vector(2960, 16),
10315 => conv_std_logic_vector(3000, 16),
10316 => conv_std_logic_vector(3040, 16),
10317 => conv_std_logic_vector(3080, 16),
10318 => conv_std_logic_vector(3120, 16),
10319 => conv_std_logic_vector(3160, 16),
10320 => conv_std_logic_vector(3200, 16),
10321 => conv_std_logic_vector(3240, 16),
10322 => conv_std_logic_vector(3280, 16),
10323 => conv_std_logic_vector(3320, 16),
10324 => conv_std_logic_vector(3360, 16),
10325 => conv_std_logic_vector(3400, 16),
10326 => conv_std_logic_vector(3440, 16),
10327 => conv_std_logic_vector(3480, 16),
10328 => conv_std_logic_vector(3520, 16),
10329 => conv_std_logic_vector(3560, 16),
10330 => conv_std_logic_vector(3600, 16),
10331 => conv_std_logic_vector(3640, 16),
10332 => conv_std_logic_vector(3680, 16),
10333 => conv_std_logic_vector(3720, 16),
10334 => conv_std_logic_vector(3760, 16),
10335 => conv_std_logic_vector(3800, 16),
10336 => conv_std_logic_vector(3840, 16),
10337 => conv_std_logic_vector(3880, 16),
10338 => conv_std_logic_vector(3920, 16),
10339 => conv_std_logic_vector(3960, 16),
10340 => conv_std_logic_vector(4000, 16),
10341 => conv_std_logic_vector(4040, 16),
10342 => conv_std_logic_vector(4080, 16),
10343 => conv_std_logic_vector(4120, 16),
10344 => conv_std_logic_vector(4160, 16),
10345 => conv_std_logic_vector(4200, 16),
10346 => conv_std_logic_vector(4240, 16),
10347 => conv_std_logic_vector(4280, 16),
10348 => conv_std_logic_vector(4320, 16),
10349 => conv_std_logic_vector(4360, 16),
10350 => conv_std_logic_vector(4400, 16),
10351 => conv_std_logic_vector(4440, 16),
10352 => conv_std_logic_vector(4480, 16),
10353 => conv_std_logic_vector(4520, 16),
10354 => conv_std_logic_vector(4560, 16),
10355 => conv_std_logic_vector(4600, 16),
10356 => conv_std_logic_vector(4640, 16),
10357 => conv_std_logic_vector(4680, 16),
10358 => conv_std_logic_vector(4720, 16),
10359 => conv_std_logic_vector(4760, 16),
10360 => conv_std_logic_vector(4800, 16),
10361 => conv_std_logic_vector(4840, 16),
10362 => conv_std_logic_vector(4880, 16),
10363 => conv_std_logic_vector(4920, 16),
10364 => conv_std_logic_vector(4960, 16),
10365 => conv_std_logic_vector(5000, 16),
10366 => conv_std_logic_vector(5040, 16),
10367 => conv_std_logic_vector(5080, 16),
10368 => conv_std_logic_vector(5120, 16),
10369 => conv_std_logic_vector(5160, 16),
10370 => conv_std_logic_vector(5200, 16),
10371 => conv_std_logic_vector(5240, 16),
10372 => conv_std_logic_vector(5280, 16),
10373 => conv_std_logic_vector(5320, 16),
10374 => conv_std_logic_vector(5360, 16),
10375 => conv_std_logic_vector(5400, 16),
10376 => conv_std_logic_vector(5440, 16),
10377 => conv_std_logic_vector(5480, 16),
10378 => conv_std_logic_vector(5520, 16),
10379 => conv_std_logic_vector(5560, 16),
10380 => conv_std_logic_vector(5600, 16),
10381 => conv_std_logic_vector(5640, 16),
10382 => conv_std_logic_vector(5680, 16),
10383 => conv_std_logic_vector(5720, 16),
10384 => conv_std_logic_vector(5760, 16),
10385 => conv_std_logic_vector(5800, 16),
10386 => conv_std_logic_vector(5840, 16),
10387 => conv_std_logic_vector(5880, 16),
10388 => conv_std_logic_vector(5920, 16),
10389 => conv_std_logic_vector(5960, 16),
10390 => conv_std_logic_vector(6000, 16),
10391 => conv_std_logic_vector(6040, 16),
10392 => conv_std_logic_vector(6080, 16),
10393 => conv_std_logic_vector(6120, 16),
10394 => conv_std_logic_vector(6160, 16),
10395 => conv_std_logic_vector(6200, 16),
10396 => conv_std_logic_vector(6240, 16),
10397 => conv_std_logic_vector(6280, 16),
10398 => conv_std_logic_vector(6320, 16),
10399 => conv_std_logic_vector(6360, 16),
10400 => conv_std_logic_vector(6400, 16),
10401 => conv_std_logic_vector(6440, 16),
10402 => conv_std_logic_vector(6480, 16),
10403 => conv_std_logic_vector(6520, 16),
10404 => conv_std_logic_vector(6560, 16),
10405 => conv_std_logic_vector(6600, 16),
10406 => conv_std_logic_vector(6640, 16),
10407 => conv_std_logic_vector(6680, 16),
10408 => conv_std_logic_vector(6720, 16),
10409 => conv_std_logic_vector(6760, 16),
10410 => conv_std_logic_vector(6800, 16),
10411 => conv_std_logic_vector(6840, 16),
10412 => conv_std_logic_vector(6880, 16),
10413 => conv_std_logic_vector(6920, 16),
10414 => conv_std_logic_vector(6960, 16),
10415 => conv_std_logic_vector(7000, 16),
10416 => conv_std_logic_vector(7040, 16),
10417 => conv_std_logic_vector(7080, 16),
10418 => conv_std_logic_vector(7120, 16),
10419 => conv_std_logic_vector(7160, 16),
10420 => conv_std_logic_vector(7200, 16),
10421 => conv_std_logic_vector(7240, 16),
10422 => conv_std_logic_vector(7280, 16),
10423 => conv_std_logic_vector(7320, 16),
10424 => conv_std_logic_vector(7360, 16),
10425 => conv_std_logic_vector(7400, 16),
10426 => conv_std_logic_vector(7440, 16),
10427 => conv_std_logic_vector(7480, 16),
10428 => conv_std_logic_vector(7520, 16),
10429 => conv_std_logic_vector(7560, 16),
10430 => conv_std_logic_vector(7600, 16),
10431 => conv_std_logic_vector(7640, 16),
10432 => conv_std_logic_vector(7680, 16),
10433 => conv_std_logic_vector(7720, 16),
10434 => conv_std_logic_vector(7760, 16),
10435 => conv_std_logic_vector(7800, 16),
10436 => conv_std_logic_vector(7840, 16),
10437 => conv_std_logic_vector(7880, 16),
10438 => conv_std_logic_vector(7920, 16),
10439 => conv_std_logic_vector(7960, 16),
10440 => conv_std_logic_vector(8000, 16),
10441 => conv_std_logic_vector(8040, 16),
10442 => conv_std_logic_vector(8080, 16),
10443 => conv_std_logic_vector(8120, 16),
10444 => conv_std_logic_vector(8160, 16),
10445 => conv_std_logic_vector(8200, 16),
10446 => conv_std_logic_vector(8240, 16),
10447 => conv_std_logic_vector(8280, 16),
10448 => conv_std_logic_vector(8320, 16),
10449 => conv_std_logic_vector(8360, 16),
10450 => conv_std_logic_vector(8400, 16),
10451 => conv_std_logic_vector(8440, 16),
10452 => conv_std_logic_vector(8480, 16),
10453 => conv_std_logic_vector(8520, 16),
10454 => conv_std_logic_vector(8560, 16),
10455 => conv_std_logic_vector(8600, 16),
10456 => conv_std_logic_vector(8640, 16),
10457 => conv_std_logic_vector(8680, 16),
10458 => conv_std_logic_vector(8720, 16),
10459 => conv_std_logic_vector(8760, 16),
10460 => conv_std_logic_vector(8800, 16),
10461 => conv_std_logic_vector(8840, 16),
10462 => conv_std_logic_vector(8880, 16),
10463 => conv_std_logic_vector(8920, 16),
10464 => conv_std_logic_vector(8960, 16),
10465 => conv_std_logic_vector(9000, 16),
10466 => conv_std_logic_vector(9040, 16),
10467 => conv_std_logic_vector(9080, 16),
10468 => conv_std_logic_vector(9120, 16),
10469 => conv_std_logic_vector(9160, 16),
10470 => conv_std_logic_vector(9200, 16),
10471 => conv_std_logic_vector(9240, 16),
10472 => conv_std_logic_vector(9280, 16),
10473 => conv_std_logic_vector(9320, 16),
10474 => conv_std_logic_vector(9360, 16),
10475 => conv_std_logic_vector(9400, 16),
10476 => conv_std_logic_vector(9440, 16),
10477 => conv_std_logic_vector(9480, 16),
10478 => conv_std_logic_vector(9520, 16),
10479 => conv_std_logic_vector(9560, 16),
10480 => conv_std_logic_vector(9600, 16),
10481 => conv_std_logic_vector(9640, 16),
10482 => conv_std_logic_vector(9680, 16),
10483 => conv_std_logic_vector(9720, 16),
10484 => conv_std_logic_vector(9760, 16),
10485 => conv_std_logic_vector(9800, 16),
10486 => conv_std_logic_vector(9840, 16),
10487 => conv_std_logic_vector(9880, 16),
10488 => conv_std_logic_vector(9920, 16),
10489 => conv_std_logic_vector(9960, 16),
10490 => conv_std_logic_vector(10000, 16),
10491 => conv_std_logic_vector(10040, 16),
10492 => conv_std_logic_vector(10080, 16),
10493 => conv_std_logic_vector(10120, 16),
10494 => conv_std_logic_vector(10160, 16),
10495 => conv_std_logic_vector(10200, 16),
10496 => conv_std_logic_vector(0, 16),
10497 => conv_std_logic_vector(41, 16),
10498 => conv_std_logic_vector(82, 16),
10499 => conv_std_logic_vector(123, 16),
10500 => conv_std_logic_vector(164, 16),
10501 => conv_std_logic_vector(205, 16),
10502 => conv_std_logic_vector(246, 16),
10503 => conv_std_logic_vector(287, 16),
10504 => conv_std_logic_vector(328, 16),
10505 => conv_std_logic_vector(369, 16),
10506 => conv_std_logic_vector(410, 16),
10507 => conv_std_logic_vector(451, 16),
10508 => conv_std_logic_vector(492, 16),
10509 => conv_std_logic_vector(533, 16),
10510 => conv_std_logic_vector(574, 16),
10511 => conv_std_logic_vector(615, 16),
10512 => conv_std_logic_vector(656, 16),
10513 => conv_std_logic_vector(697, 16),
10514 => conv_std_logic_vector(738, 16),
10515 => conv_std_logic_vector(779, 16),
10516 => conv_std_logic_vector(820, 16),
10517 => conv_std_logic_vector(861, 16),
10518 => conv_std_logic_vector(902, 16),
10519 => conv_std_logic_vector(943, 16),
10520 => conv_std_logic_vector(984, 16),
10521 => conv_std_logic_vector(1025, 16),
10522 => conv_std_logic_vector(1066, 16),
10523 => conv_std_logic_vector(1107, 16),
10524 => conv_std_logic_vector(1148, 16),
10525 => conv_std_logic_vector(1189, 16),
10526 => conv_std_logic_vector(1230, 16),
10527 => conv_std_logic_vector(1271, 16),
10528 => conv_std_logic_vector(1312, 16),
10529 => conv_std_logic_vector(1353, 16),
10530 => conv_std_logic_vector(1394, 16),
10531 => conv_std_logic_vector(1435, 16),
10532 => conv_std_logic_vector(1476, 16),
10533 => conv_std_logic_vector(1517, 16),
10534 => conv_std_logic_vector(1558, 16),
10535 => conv_std_logic_vector(1599, 16),
10536 => conv_std_logic_vector(1640, 16),
10537 => conv_std_logic_vector(1681, 16),
10538 => conv_std_logic_vector(1722, 16),
10539 => conv_std_logic_vector(1763, 16),
10540 => conv_std_logic_vector(1804, 16),
10541 => conv_std_logic_vector(1845, 16),
10542 => conv_std_logic_vector(1886, 16),
10543 => conv_std_logic_vector(1927, 16),
10544 => conv_std_logic_vector(1968, 16),
10545 => conv_std_logic_vector(2009, 16),
10546 => conv_std_logic_vector(2050, 16),
10547 => conv_std_logic_vector(2091, 16),
10548 => conv_std_logic_vector(2132, 16),
10549 => conv_std_logic_vector(2173, 16),
10550 => conv_std_logic_vector(2214, 16),
10551 => conv_std_logic_vector(2255, 16),
10552 => conv_std_logic_vector(2296, 16),
10553 => conv_std_logic_vector(2337, 16),
10554 => conv_std_logic_vector(2378, 16),
10555 => conv_std_logic_vector(2419, 16),
10556 => conv_std_logic_vector(2460, 16),
10557 => conv_std_logic_vector(2501, 16),
10558 => conv_std_logic_vector(2542, 16),
10559 => conv_std_logic_vector(2583, 16),
10560 => conv_std_logic_vector(2624, 16),
10561 => conv_std_logic_vector(2665, 16),
10562 => conv_std_logic_vector(2706, 16),
10563 => conv_std_logic_vector(2747, 16),
10564 => conv_std_logic_vector(2788, 16),
10565 => conv_std_logic_vector(2829, 16),
10566 => conv_std_logic_vector(2870, 16),
10567 => conv_std_logic_vector(2911, 16),
10568 => conv_std_logic_vector(2952, 16),
10569 => conv_std_logic_vector(2993, 16),
10570 => conv_std_logic_vector(3034, 16),
10571 => conv_std_logic_vector(3075, 16),
10572 => conv_std_logic_vector(3116, 16),
10573 => conv_std_logic_vector(3157, 16),
10574 => conv_std_logic_vector(3198, 16),
10575 => conv_std_logic_vector(3239, 16),
10576 => conv_std_logic_vector(3280, 16),
10577 => conv_std_logic_vector(3321, 16),
10578 => conv_std_logic_vector(3362, 16),
10579 => conv_std_logic_vector(3403, 16),
10580 => conv_std_logic_vector(3444, 16),
10581 => conv_std_logic_vector(3485, 16),
10582 => conv_std_logic_vector(3526, 16),
10583 => conv_std_logic_vector(3567, 16),
10584 => conv_std_logic_vector(3608, 16),
10585 => conv_std_logic_vector(3649, 16),
10586 => conv_std_logic_vector(3690, 16),
10587 => conv_std_logic_vector(3731, 16),
10588 => conv_std_logic_vector(3772, 16),
10589 => conv_std_logic_vector(3813, 16),
10590 => conv_std_logic_vector(3854, 16),
10591 => conv_std_logic_vector(3895, 16),
10592 => conv_std_logic_vector(3936, 16),
10593 => conv_std_logic_vector(3977, 16),
10594 => conv_std_logic_vector(4018, 16),
10595 => conv_std_logic_vector(4059, 16),
10596 => conv_std_logic_vector(4100, 16),
10597 => conv_std_logic_vector(4141, 16),
10598 => conv_std_logic_vector(4182, 16),
10599 => conv_std_logic_vector(4223, 16),
10600 => conv_std_logic_vector(4264, 16),
10601 => conv_std_logic_vector(4305, 16),
10602 => conv_std_logic_vector(4346, 16),
10603 => conv_std_logic_vector(4387, 16),
10604 => conv_std_logic_vector(4428, 16),
10605 => conv_std_logic_vector(4469, 16),
10606 => conv_std_logic_vector(4510, 16),
10607 => conv_std_logic_vector(4551, 16),
10608 => conv_std_logic_vector(4592, 16),
10609 => conv_std_logic_vector(4633, 16),
10610 => conv_std_logic_vector(4674, 16),
10611 => conv_std_logic_vector(4715, 16),
10612 => conv_std_logic_vector(4756, 16),
10613 => conv_std_logic_vector(4797, 16),
10614 => conv_std_logic_vector(4838, 16),
10615 => conv_std_logic_vector(4879, 16),
10616 => conv_std_logic_vector(4920, 16),
10617 => conv_std_logic_vector(4961, 16),
10618 => conv_std_logic_vector(5002, 16),
10619 => conv_std_logic_vector(5043, 16),
10620 => conv_std_logic_vector(5084, 16),
10621 => conv_std_logic_vector(5125, 16),
10622 => conv_std_logic_vector(5166, 16),
10623 => conv_std_logic_vector(5207, 16),
10624 => conv_std_logic_vector(5248, 16),
10625 => conv_std_logic_vector(5289, 16),
10626 => conv_std_logic_vector(5330, 16),
10627 => conv_std_logic_vector(5371, 16),
10628 => conv_std_logic_vector(5412, 16),
10629 => conv_std_logic_vector(5453, 16),
10630 => conv_std_logic_vector(5494, 16),
10631 => conv_std_logic_vector(5535, 16),
10632 => conv_std_logic_vector(5576, 16),
10633 => conv_std_logic_vector(5617, 16),
10634 => conv_std_logic_vector(5658, 16),
10635 => conv_std_logic_vector(5699, 16),
10636 => conv_std_logic_vector(5740, 16),
10637 => conv_std_logic_vector(5781, 16),
10638 => conv_std_logic_vector(5822, 16),
10639 => conv_std_logic_vector(5863, 16),
10640 => conv_std_logic_vector(5904, 16),
10641 => conv_std_logic_vector(5945, 16),
10642 => conv_std_logic_vector(5986, 16),
10643 => conv_std_logic_vector(6027, 16),
10644 => conv_std_logic_vector(6068, 16),
10645 => conv_std_logic_vector(6109, 16),
10646 => conv_std_logic_vector(6150, 16),
10647 => conv_std_logic_vector(6191, 16),
10648 => conv_std_logic_vector(6232, 16),
10649 => conv_std_logic_vector(6273, 16),
10650 => conv_std_logic_vector(6314, 16),
10651 => conv_std_logic_vector(6355, 16),
10652 => conv_std_logic_vector(6396, 16),
10653 => conv_std_logic_vector(6437, 16),
10654 => conv_std_logic_vector(6478, 16),
10655 => conv_std_logic_vector(6519, 16),
10656 => conv_std_logic_vector(6560, 16),
10657 => conv_std_logic_vector(6601, 16),
10658 => conv_std_logic_vector(6642, 16),
10659 => conv_std_logic_vector(6683, 16),
10660 => conv_std_logic_vector(6724, 16),
10661 => conv_std_logic_vector(6765, 16),
10662 => conv_std_logic_vector(6806, 16),
10663 => conv_std_logic_vector(6847, 16),
10664 => conv_std_logic_vector(6888, 16),
10665 => conv_std_logic_vector(6929, 16),
10666 => conv_std_logic_vector(6970, 16),
10667 => conv_std_logic_vector(7011, 16),
10668 => conv_std_logic_vector(7052, 16),
10669 => conv_std_logic_vector(7093, 16),
10670 => conv_std_logic_vector(7134, 16),
10671 => conv_std_logic_vector(7175, 16),
10672 => conv_std_logic_vector(7216, 16),
10673 => conv_std_logic_vector(7257, 16),
10674 => conv_std_logic_vector(7298, 16),
10675 => conv_std_logic_vector(7339, 16),
10676 => conv_std_logic_vector(7380, 16),
10677 => conv_std_logic_vector(7421, 16),
10678 => conv_std_logic_vector(7462, 16),
10679 => conv_std_logic_vector(7503, 16),
10680 => conv_std_logic_vector(7544, 16),
10681 => conv_std_logic_vector(7585, 16),
10682 => conv_std_logic_vector(7626, 16),
10683 => conv_std_logic_vector(7667, 16),
10684 => conv_std_logic_vector(7708, 16),
10685 => conv_std_logic_vector(7749, 16),
10686 => conv_std_logic_vector(7790, 16),
10687 => conv_std_logic_vector(7831, 16),
10688 => conv_std_logic_vector(7872, 16),
10689 => conv_std_logic_vector(7913, 16),
10690 => conv_std_logic_vector(7954, 16),
10691 => conv_std_logic_vector(7995, 16),
10692 => conv_std_logic_vector(8036, 16),
10693 => conv_std_logic_vector(8077, 16),
10694 => conv_std_logic_vector(8118, 16),
10695 => conv_std_logic_vector(8159, 16),
10696 => conv_std_logic_vector(8200, 16),
10697 => conv_std_logic_vector(8241, 16),
10698 => conv_std_logic_vector(8282, 16),
10699 => conv_std_logic_vector(8323, 16),
10700 => conv_std_logic_vector(8364, 16),
10701 => conv_std_logic_vector(8405, 16),
10702 => conv_std_logic_vector(8446, 16),
10703 => conv_std_logic_vector(8487, 16),
10704 => conv_std_logic_vector(8528, 16),
10705 => conv_std_logic_vector(8569, 16),
10706 => conv_std_logic_vector(8610, 16),
10707 => conv_std_logic_vector(8651, 16),
10708 => conv_std_logic_vector(8692, 16),
10709 => conv_std_logic_vector(8733, 16),
10710 => conv_std_logic_vector(8774, 16),
10711 => conv_std_logic_vector(8815, 16),
10712 => conv_std_logic_vector(8856, 16),
10713 => conv_std_logic_vector(8897, 16),
10714 => conv_std_logic_vector(8938, 16),
10715 => conv_std_logic_vector(8979, 16),
10716 => conv_std_logic_vector(9020, 16),
10717 => conv_std_logic_vector(9061, 16),
10718 => conv_std_logic_vector(9102, 16),
10719 => conv_std_logic_vector(9143, 16),
10720 => conv_std_logic_vector(9184, 16),
10721 => conv_std_logic_vector(9225, 16),
10722 => conv_std_logic_vector(9266, 16),
10723 => conv_std_logic_vector(9307, 16),
10724 => conv_std_logic_vector(9348, 16),
10725 => conv_std_logic_vector(9389, 16),
10726 => conv_std_logic_vector(9430, 16),
10727 => conv_std_logic_vector(9471, 16),
10728 => conv_std_logic_vector(9512, 16),
10729 => conv_std_logic_vector(9553, 16),
10730 => conv_std_logic_vector(9594, 16),
10731 => conv_std_logic_vector(9635, 16),
10732 => conv_std_logic_vector(9676, 16),
10733 => conv_std_logic_vector(9717, 16),
10734 => conv_std_logic_vector(9758, 16),
10735 => conv_std_logic_vector(9799, 16),
10736 => conv_std_logic_vector(9840, 16),
10737 => conv_std_logic_vector(9881, 16),
10738 => conv_std_logic_vector(9922, 16),
10739 => conv_std_logic_vector(9963, 16),
10740 => conv_std_logic_vector(10004, 16),
10741 => conv_std_logic_vector(10045, 16),
10742 => conv_std_logic_vector(10086, 16),
10743 => conv_std_logic_vector(10127, 16),
10744 => conv_std_logic_vector(10168, 16),
10745 => conv_std_logic_vector(10209, 16),
10746 => conv_std_logic_vector(10250, 16),
10747 => conv_std_logic_vector(10291, 16),
10748 => conv_std_logic_vector(10332, 16),
10749 => conv_std_logic_vector(10373, 16),
10750 => conv_std_logic_vector(10414, 16),
10751 => conv_std_logic_vector(10455, 16),
10752 => conv_std_logic_vector(0, 16),
10753 => conv_std_logic_vector(42, 16),
10754 => conv_std_logic_vector(84, 16),
10755 => conv_std_logic_vector(126, 16),
10756 => conv_std_logic_vector(168, 16),
10757 => conv_std_logic_vector(210, 16),
10758 => conv_std_logic_vector(252, 16),
10759 => conv_std_logic_vector(294, 16),
10760 => conv_std_logic_vector(336, 16),
10761 => conv_std_logic_vector(378, 16),
10762 => conv_std_logic_vector(420, 16),
10763 => conv_std_logic_vector(462, 16),
10764 => conv_std_logic_vector(504, 16),
10765 => conv_std_logic_vector(546, 16),
10766 => conv_std_logic_vector(588, 16),
10767 => conv_std_logic_vector(630, 16),
10768 => conv_std_logic_vector(672, 16),
10769 => conv_std_logic_vector(714, 16),
10770 => conv_std_logic_vector(756, 16),
10771 => conv_std_logic_vector(798, 16),
10772 => conv_std_logic_vector(840, 16),
10773 => conv_std_logic_vector(882, 16),
10774 => conv_std_logic_vector(924, 16),
10775 => conv_std_logic_vector(966, 16),
10776 => conv_std_logic_vector(1008, 16),
10777 => conv_std_logic_vector(1050, 16),
10778 => conv_std_logic_vector(1092, 16),
10779 => conv_std_logic_vector(1134, 16),
10780 => conv_std_logic_vector(1176, 16),
10781 => conv_std_logic_vector(1218, 16),
10782 => conv_std_logic_vector(1260, 16),
10783 => conv_std_logic_vector(1302, 16),
10784 => conv_std_logic_vector(1344, 16),
10785 => conv_std_logic_vector(1386, 16),
10786 => conv_std_logic_vector(1428, 16),
10787 => conv_std_logic_vector(1470, 16),
10788 => conv_std_logic_vector(1512, 16),
10789 => conv_std_logic_vector(1554, 16),
10790 => conv_std_logic_vector(1596, 16),
10791 => conv_std_logic_vector(1638, 16),
10792 => conv_std_logic_vector(1680, 16),
10793 => conv_std_logic_vector(1722, 16),
10794 => conv_std_logic_vector(1764, 16),
10795 => conv_std_logic_vector(1806, 16),
10796 => conv_std_logic_vector(1848, 16),
10797 => conv_std_logic_vector(1890, 16),
10798 => conv_std_logic_vector(1932, 16),
10799 => conv_std_logic_vector(1974, 16),
10800 => conv_std_logic_vector(2016, 16),
10801 => conv_std_logic_vector(2058, 16),
10802 => conv_std_logic_vector(2100, 16),
10803 => conv_std_logic_vector(2142, 16),
10804 => conv_std_logic_vector(2184, 16),
10805 => conv_std_logic_vector(2226, 16),
10806 => conv_std_logic_vector(2268, 16),
10807 => conv_std_logic_vector(2310, 16),
10808 => conv_std_logic_vector(2352, 16),
10809 => conv_std_logic_vector(2394, 16),
10810 => conv_std_logic_vector(2436, 16),
10811 => conv_std_logic_vector(2478, 16),
10812 => conv_std_logic_vector(2520, 16),
10813 => conv_std_logic_vector(2562, 16),
10814 => conv_std_logic_vector(2604, 16),
10815 => conv_std_logic_vector(2646, 16),
10816 => conv_std_logic_vector(2688, 16),
10817 => conv_std_logic_vector(2730, 16),
10818 => conv_std_logic_vector(2772, 16),
10819 => conv_std_logic_vector(2814, 16),
10820 => conv_std_logic_vector(2856, 16),
10821 => conv_std_logic_vector(2898, 16),
10822 => conv_std_logic_vector(2940, 16),
10823 => conv_std_logic_vector(2982, 16),
10824 => conv_std_logic_vector(3024, 16),
10825 => conv_std_logic_vector(3066, 16),
10826 => conv_std_logic_vector(3108, 16),
10827 => conv_std_logic_vector(3150, 16),
10828 => conv_std_logic_vector(3192, 16),
10829 => conv_std_logic_vector(3234, 16),
10830 => conv_std_logic_vector(3276, 16),
10831 => conv_std_logic_vector(3318, 16),
10832 => conv_std_logic_vector(3360, 16),
10833 => conv_std_logic_vector(3402, 16),
10834 => conv_std_logic_vector(3444, 16),
10835 => conv_std_logic_vector(3486, 16),
10836 => conv_std_logic_vector(3528, 16),
10837 => conv_std_logic_vector(3570, 16),
10838 => conv_std_logic_vector(3612, 16),
10839 => conv_std_logic_vector(3654, 16),
10840 => conv_std_logic_vector(3696, 16),
10841 => conv_std_logic_vector(3738, 16),
10842 => conv_std_logic_vector(3780, 16),
10843 => conv_std_logic_vector(3822, 16),
10844 => conv_std_logic_vector(3864, 16),
10845 => conv_std_logic_vector(3906, 16),
10846 => conv_std_logic_vector(3948, 16),
10847 => conv_std_logic_vector(3990, 16),
10848 => conv_std_logic_vector(4032, 16),
10849 => conv_std_logic_vector(4074, 16),
10850 => conv_std_logic_vector(4116, 16),
10851 => conv_std_logic_vector(4158, 16),
10852 => conv_std_logic_vector(4200, 16),
10853 => conv_std_logic_vector(4242, 16),
10854 => conv_std_logic_vector(4284, 16),
10855 => conv_std_logic_vector(4326, 16),
10856 => conv_std_logic_vector(4368, 16),
10857 => conv_std_logic_vector(4410, 16),
10858 => conv_std_logic_vector(4452, 16),
10859 => conv_std_logic_vector(4494, 16),
10860 => conv_std_logic_vector(4536, 16),
10861 => conv_std_logic_vector(4578, 16),
10862 => conv_std_logic_vector(4620, 16),
10863 => conv_std_logic_vector(4662, 16),
10864 => conv_std_logic_vector(4704, 16),
10865 => conv_std_logic_vector(4746, 16),
10866 => conv_std_logic_vector(4788, 16),
10867 => conv_std_logic_vector(4830, 16),
10868 => conv_std_logic_vector(4872, 16),
10869 => conv_std_logic_vector(4914, 16),
10870 => conv_std_logic_vector(4956, 16),
10871 => conv_std_logic_vector(4998, 16),
10872 => conv_std_logic_vector(5040, 16),
10873 => conv_std_logic_vector(5082, 16),
10874 => conv_std_logic_vector(5124, 16),
10875 => conv_std_logic_vector(5166, 16),
10876 => conv_std_logic_vector(5208, 16),
10877 => conv_std_logic_vector(5250, 16),
10878 => conv_std_logic_vector(5292, 16),
10879 => conv_std_logic_vector(5334, 16),
10880 => conv_std_logic_vector(5376, 16),
10881 => conv_std_logic_vector(5418, 16),
10882 => conv_std_logic_vector(5460, 16),
10883 => conv_std_logic_vector(5502, 16),
10884 => conv_std_logic_vector(5544, 16),
10885 => conv_std_logic_vector(5586, 16),
10886 => conv_std_logic_vector(5628, 16),
10887 => conv_std_logic_vector(5670, 16),
10888 => conv_std_logic_vector(5712, 16),
10889 => conv_std_logic_vector(5754, 16),
10890 => conv_std_logic_vector(5796, 16),
10891 => conv_std_logic_vector(5838, 16),
10892 => conv_std_logic_vector(5880, 16),
10893 => conv_std_logic_vector(5922, 16),
10894 => conv_std_logic_vector(5964, 16),
10895 => conv_std_logic_vector(6006, 16),
10896 => conv_std_logic_vector(6048, 16),
10897 => conv_std_logic_vector(6090, 16),
10898 => conv_std_logic_vector(6132, 16),
10899 => conv_std_logic_vector(6174, 16),
10900 => conv_std_logic_vector(6216, 16),
10901 => conv_std_logic_vector(6258, 16),
10902 => conv_std_logic_vector(6300, 16),
10903 => conv_std_logic_vector(6342, 16),
10904 => conv_std_logic_vector(6384, 16),
10905 => conv_std_logic_vector(6426, 16),
10906 => conv_std_logic_vector(6468, 16),
10907 => conv_std_logic_vector(6510, 16),
10908 => conv_std_logic_vector(6552, 16),
10909 => conv_std_logic_vector(6594, 16),
10910 => conv_std_logic_vector(6636, 16),
10911 => conv_std_logic_vector(6678, 16),
10912 => conv_std_logic_vector(6720, 16),
10913 => conv_std_logic_vector(6762, 16),
10914 => conv_std_logic_vector(6804, 16),
10915 => conv_std_logic_vector(6846, 16),
10916 => conv_std_logic_vector(6888, 16),
10917 => conv_std_logic_vector(6930, 16),
10918 => conv_std_logic_vector(6972, 16),
10919 => conv_std_logic_vector(7014, 16),
10920 => conv_std_logic_vector(7056, 16),
10921 => conv_std_logic_vector(7098, 16),
10922 => conv_std_logic_vector(7140, 16),
10923 => conv_std_logic_vector(7182, 16),
10924 => conv_std_logic_vector(7224, 16),
10925 => conv_std_logic_vector(7266, 16),
10926 => conv_std_logic_vector(7308, 16),
10927 => conv_std_logic_vector(7350, 16),
10928 => conv_std_logic_vector(7392, 16),
10929 => conv_std_logic_vector(7434, 16),
10930 => conv_std_logic_vector(7476, 16),
10931 => conv_std_logic_vector(7518, 16),
10932 => conv_std_logic_vector(7560, 16),
10933 => conv_std_logic_vector(7602, 16),
10934 => conv_std_logic_vector(7644, 16),
10935 => conv_std_logic_vector(7686, 16),
10936 => conv_std_logic_vector(7728, 16),
10937 => conv_std_logic_vector(7770, 16),
10938 => conv_std_logic_vector(7812, 16),
10939 => conv_std_logic_vector(7854, 16),
10940 => conv_std_logic_vector(7896, 16),
10941 => conv_std_logic_vector(7938, 16),
10942 => conv_std_logic_vector(7980, 16),
10943 => conv_std_logic_vector(8022, 16),
10944 => conv_std_logic_vector(8064, 16),
10945 => conv_std_logic_vector(8106, 16),
10946 => conv_std_logic_vector(8148, 16),
10947 => conv_std_logic_vector(8190, 16),
10948 => conv_std_logic_vector(8232, 16),
10949 => conv_std_logic_vector(8274, 16),
10950 => conv_std_logic_vector(8316, 16),
10951 => conv_std_logic_vector(8358, 16),
10952 => conv_std_logic_vector(8400, 16),
10953 => conv_std_logic_vector(8442, 16),
10954 => conv_std_logic_vector(8484, 16),
10955 => conv_std_logic_vector(8526, 16),
10956 => conv_std_logic_vector(8568, 16),
10957 => conv_std_logic_vector(8610, 16),
10958 => conv_std_logic_vector(8652, 16),
10959 => conv_std_logic_vector(8694, 16),
10960 => conv_std_logic_vector(8736, 16),
10961 => conv_std_logic_vector(8778, 16),
10962 => conv_std_logic_vector(8820, 16),
10963 => conv_std_logic_vector(8862, 16),
10964 => conv_std_logic_vector(8904, 16),
10965 => conv_std_logic_vector(8946, 16),
10966 => conv_std_logic_vector(8988, 16),
10967 => conv_std_logic_vector(9030, 16),
10968 => conv_std_logic_vector(9072, 16),
10969 => conv_std_logic_vector(9114, 16),
10970 => conv_std_logic_vector(9156, 16),
10971 => conv_std_logic_vector(9198, 16),
10972 => conv_std_logic_vector(9240, 16),
10973 => conv_std_logic_vector(9282, 16),
10974 => conv_std_logic_vector(9324, 16),
10975 => conv_std_logic_vector(9366, 16),
10976 => conv_std_logic_vector(9408, 16),
10977 => conv_std_logic_vector(9450, 16),
10978 => conv_std_logic_vector(9492, 16),
10979 => conv_std_logic_vector(9534, 16),
10980 => conv_std_logic_vector(9576, 16),
10981 => conv_std_logic_vector(9618, 16),
10982 => conv_std_logic_vector(9660, 16),
10983 => conv_std_logic_vector(9702, 16),
10984 => conv_std_logic_vector(9744, 16),
10985 => conv_std_logic_vector(9786, 16),
10986 => conv_std_logic_vector(9828, 16),
10987 => conv_std_logic_vector(9870, 16),
10988 => conv_std_logic_vector(9912, 16),
10989 => conv_std_logic_vector(9954, 16),
10990 => conv_std_logic_vector(9996, 16),
10991 => conv_std_logic_vector(10038, 16),
10992 => conv_std_logic_vector(10080, 16),
10993 => conv_std_logic_vector(10122, 16),
10994 => conv_std_logic_vector(10164, 16),
10995 => conv_std_logic_vector(10206, 16),
10996 => conv_std_logic_vector(10248, 16),
10997 => conv_std_logic_vector(10290, 16),
10998 => conv_std_logic_vector(10332, 16),
10999 => conv_std_logic_vector(10374, 16),
11000 => conv_std_logic_vector(10416, 16),
11001 => conv_std_logic_vector(10458, 16),
11002 => conv_std_logic_vector(10500, 16),
11003 => conv_std_logic_vector(10542, 16),
11004 => conv_std_logic_vector(10584, 16),
11005 => conv_std_logic_vector(10626, 16),
11006 => conv_std_logic_vector(10668, 16),
11007 => conv_std_logic_vector(10710, 16),
11008 => conv_std_logic_vector(0, 16),
11009 => conv_std_logic_vector(43, 16),
11010 => conv_std_logic_vector(86, 16),
11011 => conv_std_logic_vector(129, 16),
11012 => conv_std_logic_vector(172, 16),
11013 => conv_std_logic_vector(215, 16),
11014 => conv_std_logic_vector(258, 16),
11015 => conv_std_logic_vector(301, 16),
11016 => conv_std_logic_vector(344, 16),
11017 => conv_std_logic_vector(387, 16),
11018 => conv_std_logic_vector(430, 16),
11019 => conv_std_logic_vector(473, 16),
11020 => conv_std_logic_vector(516, 16),
11021 => conv_std_logic_vector(559, 16),
11022 => conv_std_logic_vector(602, 16),
11023 => conv_std_logic_vector(645, 16),
11024 => conv_std_logic_vector(688, 16),
11025 => conv_std_logic_vector(731, 16),
11026 => conv_std_logic_vector(774, 16),
11027 => conv_std_logic_vector(817, 16),
11028 => conv_std_logic_vector(860, 16),
11029 => conv_std_logic_vector(903, 16),
11030 => conv_std_logic_vector(946, 16),
11031 => conv_std_logic_vector(989, 16),
11032 => conv_std_logic_vector(1032, 16),
11033 => conv_std_logic_vector(1075, 16),
11034 => conv_std_logic_vector(1118, 16),
11035 => conv_std_logic_vector(1161, 16),
11036 => conv_std_logic_vector(1204, 16),
11037 => conv_std_logic_vector(1247, 16),
11038 => conv_std_logic_vector(1290, 16),
11039 => conv_std_logic_vector(1333, 16),
11040 => conv_std_logic_vector(1376, 16),
11041 => conv_std_logic_vector(1419, 16),
11042 => conv_std_logic_vector(1462, 16),
11043 => conv_std_logic_vector(1505, 16),
11044 => conv_std_logic_vector(1548, 16),
11045 => conv_std_logic_vector(1591, 16),
11046 => conv_std_logic_vector(1634, 16),
11047 => conv_std_logic_vector(1677, 16),
11048 => conv_std_logic_vector(1720, 16),
11049 => conv_std_logic_vector(1763, 16),
11050 => conv_std_logic_vector(1806, 16),
11051 => conv_std_logic_vector(1849, 16),
11052 => conv_std_logic_vector(1892, 16),
11053 => conv_std_logic_vector(1935, 16),
11054 => conv_std_logic_vector(1978, 16),
11055 => conv_std_logic_vector(2021, 16),
11056 => conv_std_logic_vector(2064, 16),
11057 => conv_std_logic_vector(2107, 16),
11058 => conv_std_logic_vector(2150, 16),
11059 => conv_std_logic_vector(2193, 16),
11060 => conv_std_logic_vector(2236, 16),
11061 => conv_std_logic_vector(2279, 16),
11062 => conv_std_logic_vector(2322, 16),
11063 => conv_std_logic_vector(2365, 16),
11064 => conv_std_logic_vector(2408, 16),
11065 => conv_std_logic_vector(2451, 16),
11066 => conv_std_logic_vector(2494, 16),
11067 => conv_std_logic_vector(2537, 16),
11068 => conv_std_logic_vector(2580, 16),
11069 => conv_std_logic_vector(2623, 16),
11070 => conv_std_logic_vector(2666, 16),
11071 => conv_std_logic_vector(2709, 16),
11072 => conv_std_logic_vector(2752, 16),
11073 => conv_std_logic_vector(2795, 16),
11074 => conv_std_logic_vector(2838, 16),
11075 => conv_std_logic_vector(2881, 16),
11076 => conv_std_logic_vector(2924, 16),
11077 => conv_std_logic_vector(2967, 16),
11078 => conv_std_logic_vector(3010, 16),
11079 => conv_std_logic_vector(3053, 16),
11080 => conv_std_logic_vector(3096, 16),
11081 => conv_std_logic_vector(3139, 16),
11082 => conv_std_logic_vector(3182, 16),
11083 => conv_std_logic_vector(3225, 16),
11084 => conv_std_logic_vector(3268, 16),
11085 => conv_std_logic_vector(3311, 16),
11086 => conv_std_logic_vector(3354, 16),
11087 => conv_std_logic_vector(3397, 16),
11088 => conv_std_logic_vector(3440, 16),
11089 => conv_std_logic_vector(3483, 16),
11090 => conv_std_logic_vector(3526, 16),
11091 => conv_std_logic_vector(3569, 16),
11092 => conv_std_logic_vector(3612, 16),
11093 => conv_std_logic_vector(3655, 16),
11094 => conv_std_logic_vector(3698, 16),
11095 => conv_std_logic_vector(3741, 16),
11096 => conv_std_logic_vector(3784, 16),
11097 => conv_std_logic_vector(3827, 16),
11098 => conv_std_logic_vector(3870, 16),
11099 => conv_std_logic_vector(3913, 16),
11100 => conv_std_logic_vector(3956, 16),
11101 => conv_std_logic_vector(3999, 16),
11102 => conv_std_logic_vector(4042, 16),
11103 => conv_std_logic_vector(4085, 16),
11104 => conv_std_logic_vector(4128, 16),
11105 => conv_std_logic_vector(4171, 16),
11106 => conv_std_logic_vector(4214, 16),
11107 => conv_std_logic_vector(4257, 16),
11108 => conv_std_logic_vector(4300, 16),
11109 => conv_std_logic_vector(4343, 16),
11110 => conv_std_logic_vector(4386, 16),
11111 => conv_std_logic_vector(4429, 16),
11112 => conv_std_logic_vector(4472, 16),
11113 => conv_std_logic_vector(4515, 16),
11114 => conv_std_logic_vector(4558, 16),
11115 => conv_std_logic_vector(4601, 16),
11116 => conv_std_logic_vector(4644, 16),
11117 => conv_std_logic_vector(4687, 16),
11118 => conv_std_logic_vector(4730, 16),
11119 => conv_std_logic_vector(4773, 16),
11120 => conv_std_logic_vector(4816, 16),
11121 => conv_std_logic_vector(4859, 16),
11122 => conv_std_logic_vector(4902, 16),
11123 => conv_std_logic_vector(4945, 16),
11124 => conv_std_logic_vector(4988, 16),
11125 => conv_std_logic_vector(5031, 16),
11126 => conv_std_logic_vector(5074, 16),
11127 => conv_std_logic_vector(5117, 16),
11128 => conv_std_logic_vector(5160, 16),
11129 => conv_std_logic_vector(5203, 16),
11130 => conv_std_logic_vector(5246, 16),
11131 => conv_std_logic_vector(5289, 16),
11132 => conv_std_logic_vector(5332, 16),
11133 => conv_std_logic_vector(5375, 16),
11134 => conv_std_logic_vector(5418, 16),
11135 => conv_std_logic_vector(5461, 16),
11136 => conv_std_logic_vector(5504, 16),
11137 => conv_std_logic_vector(5547, 16),
11138 => conv_std_logic_vector(5590, 16),
11139 => conv_std_logic_vector(5633, 16),
11140 => conv_std_logic_vector(5676, 16),
11141 => conv_std_logic_vector(5719, 16),
11142 => conv_std_logic_vector(5762, 16),
11143 => conv_std_logic_vector(5805, 16),
11144 => conv_std_logic_vector(5848, 16),
11145 => conv_std_logic_vector(5891, 16),
11146 => conv_std_logic_vector(5934, 16),
11147 => conv_std_logic_vector(5977, 16),
11148 => conv_std_logic_vector(6020, 16),
11149 => conv_std_logic_vector(6063, 16),
11150 => conv_std_logic_vector(6106, 16),
11151 => conv_std_logic_vector(6149, 16),
11152 => conv_std_logic_vector(6192, 16),
11153 => conv_std_logic_vector(6235, 16),
11154 => conv_std_logic_vector(6278, 16),
11155 => conv_std_logic_vector(6321, 16),
11156 => conv_std_logic_vector(6364, 16),
11157 => conv_std_logic_vector(6407, 16),
11158 => conv_std_logic_vector(6450, 16),
11159 => conv_std_logic_vector(6493, 16),
11160 => conv_std_logic_vector(6536, 16),
11161 => conv_std_logic_vector(6579, 16),
11162 => conv_std_logic_vector(6622, 16),
11163 => conv_std_logic_vector(6665, 16),
11164 => conv_std_logic_vector(6708, 16),
11165 => conv_std_logic_vector(6751, 16),
11166 => conv_std_logic_vector(6794, 16),
11167 => conv_std_logic_vector(6837, 16),
11168 => conv_std_logic_vector(6880, 16),
11169 => conv_std_logic_vector(6923, 16),
11170 => conv_std_logic_vector(6966, 16),
11171 => conv_std_logic_vector(7009, 16),
11172 => conv_std_logic_vector(7052, 16),
11173 => conv_std_logic_vector(7095, 16),
11174 => conv_std_logic_vector(7138, 16),
11175 => conv_std_logic_vector(7181, 16),
11176 => conv_std_logic_vector(7224, 16),
11177 => conv_std_logic_vector(7267, 16),
11178 => conv_std_logic_vector(7310, 16),
11179 => conv_std_logic_vector(7353, 16),
11180 => conv_std_logic_vector(7396, 16),
11181 => conv_std_logic_vector(7439, 16),
11182 => conv_std_logic_vector(7482, 16),
11183 => conv_std_logic_vector(7525, 16),
11184 => conv_std_logic_vector(7568, 16),
11185 => conv_std_logic_vector(7611, 16),
11186 => conv_std_logic_vector(7654, 16),
11187 => conv_std_logic_vector(7697, 16),
11188 => conv_std_logic_vector(7740, 16),
11189 => conv_std_logic_vector(7783, 16),
11190 => conv_std_logic_vector(7826, 16),
11191 => conv_std_logic_vector(7869, 16),
11192 => conv_std_logic_vector(7912, 16),
11193 => conv_std_logic_vector(7955, 16),
11194 => conv_std_logic_vector(7998, 16),
11195 => conv_std_logic_vector(8041, 16),
11196 => conv_std_logic_vector(8084, 16),
11197 => conv_std_logic_vector(8127, 16),
11198 => conv_std_logic_vector(8170, 16),
11199 => conv_std_logic_vector(8213, 16),
11200 => conv_std_logic_vector(8256, 16),
11201 => conv_std_logic_vector(8299, 16),
11202 => conv_std_logic_vector(8342, 16),
11203 => conv_std_logic_vector(8385, 16),
11204 => conv_std_logic_vector(8428, 16),
11205 => conv_std_logic_vector(8471, 16),
11206 => conv_std_logic_vector(8514, 16),
11207 => conv_std_logic_vector(8557, 16),
11208 => conv_std_logic_vector(8600, 16),
11209 => conv_std_logic_vector(8643, 16),
11210 => conv_std_logic_vector(8686, 16),
11211 => conv_std_logic_vector(8729, 16),
11212 => conv_std_logic_vector(8772, 16),
11213 => conv_std_logic_vector(8815, 16),
11214 => conv_std_logic_vector(8858, 16),
11215 => conv_std_logic_vector(8901, 16),
11216 => conv_std_logic_vector(8944, 16),
11217 => conv_std_logic_vector(8987, 16),
11218 => conv_std_logic_vector(9030, 16),
11219 => conv_std_logic_vector(9073, 16),
11220 => conv_std_logic_vector(9116, 16),
11221 => conv_std_logic_vector(9159, 16),
11222 => conv_std_logic_vector(9202, 16),
11223 => conv_std_logic_vector(9245, 16),
11224 => conv_std_logic_vector(9288, 16),
11225 => conv_std_logic_vector(9331, 16),
11226 => conv_std_logic_vector(9374, 16),
11227 => conv_std_logic_vector(9417, 16),
11228 => conv_std_logic_vector(9460, 16),
11229 => conv_std_logic_vector(9503, 16),
11230 => conv_std_logic_vector(9546, 16),
11231 => conv_std_logic_vector(9589, 16),
11232 => conv_std_logic_vector(9632, 16),
11233 => conv_std_logic_vector(9675, 16),
11234 => conv_std_logic_vector(9718, 16),
11235 => conv_std_logic_vector(9761, 16),
11236 => conv_std_logic_vector(9804, 16),
11237 => conv_std_logic_vector(9847, 16),
11238 => conv_std_logic_vector(9890, 16),
11239 => conv_std_logic_vector(9933, 16),
11240 => conv_std_logic_vector(9976, 16),
11241 => conv_std_logic_vector(10019, 16),
11242 => conv_std_logic_vector(10062, 16),
11243 => conv_std_logic_vector(10105, 16),
11244 => conv_std_logic_vector(10148, 16),
11245 => conv_std_logic_vector(10191, 16),
11246 => conv_std_logic_vector(10234, 16),
11247 => conv_std_logic_vector(10277, 16),
11248 => conv_std_logic_vector(10320, 16),
11249 => conv_std_logic_vector(10363, 16),
11250 => conv_std_logic_vector(10406, 16),
11251 => conv_std_logic_vector(10449, 16),
11252 => conv_std_logic_vector(10492, 16),
11253 => conv_std_logic_vector(10535, 16),
11254 => conv_std_logic_vector(10578, 16),
11255 => conv_std_logic_vector(10621, 16),
11256 => conv_std_logic_vector(10664, 16),
11257 => conv_std_logic_vector(10707, 16),
11258 => conv_std_logic_vector(10750, 16),
11259 => conv_std_logic_vector(10793, 16),
11260 => conv_std_logic_vector(10836, 16),
11261 => conv_std_logic_vector(10879, 16),
11262 => conv_std_logic_vector(10922, 16),
11263 => conv_std_logic_vector(10965, 16),
11264 => conv_std_logic_vector(0, 16),
11265 => conv_std_logic_vector(44, 16),
11266 => conv_std_logic_vector(88, 16),
11267 => conv_std_logic_vector(132, 16),
11268 => conv_std_logic_vector(176, 16),
11269 => conv_std_logic_vector(220, 16),
11270 => conv_std_logic_vector(264, 16),
11271 => conv_std_logic_vector(308, 16),
11272 => conv_std_logic_vector(352, 16),
11273 => conv_std_logic_vector(396, 16),
11274 => conv_std_logic_vector(440, 16),
11275 => conv_std_logic_vector(484, 16),
11276 => conv_std_logic_vector(528, 16),
11277 => conv_std_logic_vector(572, 16),
11278 => conv_std_logic_vector(616, 16),
11279 => conv_std_logic_vector(660, 16),
11280 => conv_std_logic_vector(704, 16),
11281 => conv_std_logic_vector(748, 16),
11282 => conv_std_logic_vector(792, 16),
11283 => conv_std_logic_vector(836, 16),
11284 => conv_std_logic_vector(880, 16),
11285 => conv_std_logic_vector(924, 16),
11286 => conv_std_logic_vector(968, 16),
11287 => conv_std_logic_vector(1012, 16),
11288 => conv_std_logic_vector(1056, 16),
11289 => conv_std_logic_vector(1100, 16),
11290 => conv_std_logic_vector(1144, 16),
11291 => conv_std_logic_vector(1188, 16),
11292 => conv_std_logic_vector(1232, 16),
11293 => conv_std_logic_vector(1276, 16),
11294 => conv_std_logic_vector(1320, 16),
11295 => conv_std_logic_vector(1364, 16),
11296 => conv_std_logic_vector(1408, 16),
11297 => conv_std_logic_vector(1452, 16),
11298 => conv_std_logic_vector(1496, 16),
11299 => conv_std_logic_vector(1540, 16),
11300 => conv_std_logic_vector(1584, 16),
11301 => conv_std_logic_vector(1628, 16),
11302 => conv_std_logic_vector(1672, 16),
11303 => conv_std_logic_vector(1716, 16),
11304 => conv_std_logic_vector(1760, 16),
11305 => conv_std_logic_vector(1804, 16),
11306 => conv_std_logic_vector(1848, 16),
11307 => conv_std_logic_vector(1892, 16),
11308 => conv_std_logic_vector(1936, 16),
11309 => conv_std_logic_vector(1980, 16),
11310 => conv_std_logic_vector(2024, 16),
11311 => conv_std_logic_vector(2068, 16),
11312 => conv_std_logic_vector(2112, 16),
11313 => conv_std_logic_vector(2156, 16),
11314 => conv_std_logic_vector(2200, 16),
11315 => conv_std_logic_vector(2244, 16),
11316 => conv_std_logic_vector(2288, 16),
11317 => conv_std_logic_vector(2332, 16),
11318 => conv_std_logic_vector(2376, 16),
11319 => conv_std_logic_vector(2420, 16),
11320 => conv_std_logic_vector(2464, 16),
11321 => conv_std_logic_vector(2508, 16),
11322 => conv_std_logic_vector(2552, 16),
11323 => conv_std_logic_vector(2596, 16),
11324 => conv_std_logic_vector(2640, 16),
11325 => conv_std_logic_vector(2684, 16),
11326 => conv_std_logic_vector(2728, 16),
11327 => conv_std_logic_vector(2772, 16),
11328 => conv_std_logic_vector(2816, 16),
11329 => conv_std_logic_vector(2860, 16),
11330 => conv_std_logic_vector(2904, 16),
11331 => conv_std_logic_vector(2948, 16),
11332 => conv_std_logic_vector(2992, 16),
11333 => conv_std_logic_vector(3036, 16),
11334 => conv_std_logic_vector(3080, 16),
11335 => conv_std_logic_vector(3124, 16),
11336 => conv_std_logic_vector(3168, 16),
11337 => conv_std_logic_vector(3212, 16),
11338 => conv_std_logic_vector(3256, 16),
11339 => conv_std_logic_vector(3300, 16),
11340 => conv_std_logic_vector(3344, 16),
11341 => conv_std_logic_vector(3388, 16),
11342 => conv_std_logic_vector(3432, 16),
11343 => conv_std_logic_vector(3476, 16),
11344 => conv_std_logic_vector(3520, 16),
11345 => conv_std_logic_vector(3564, 16),
11346 => conv_std_logic_vector(3608, 16),
11347 => conv_std_logic_vector(3652, 16),
11348 => conv_std_logic_vector(3696, 16),
11349 => conv_std_logic_vector(3740, 16),
11350 => conv_std_logic_vector(3784, 16),
11351 => conv_std_logic_vector(3828, 16),
11352 => conv_std_logic_vector(3872, 16),
11353 => conv_std_logic_vector(3916, 16),
11354 => conv_std_logic_vector(3960, 16),
11355 => conv_std_logic_vector(4004, 16),
11356 => conv_std_logic_vector(4048, 16),
11357 => conv_std_logic_vector(4092, 16),
11358 => conv_std_logic_vector(4136, 16),
11359 => conv_std_logic_vector(4180, 16),
11360 => conv_std_logic_vector(4224, 16),
11361 => conv_std_logic_vector(4268, 16),
11362 => conv_std_logic_vector(4312, 16),
11363 => conv_std_logic_vector(4356, 16),
11364 => conv_std_logic_vector(4400, 16),
11365 => conv_std_logic_vector(4444, 16),
11366 => conv_std_logic_vector(4488, 16),
11367 => conv_std_logic_vector(4532, 16),
11368 => conv_std_logic_vector(4576, 16),
11369 => conv_std_logic_vector(4620, 16),
11370 => conv_std_logic_vector(4664, 16),
11371 => conv_std_logic_vector(4708, 16),
11372 => conv_std_logic_vector(4752, 16),
11373 => conv_std_logic_vector(4796, 16),
11374 => conv_std_logic_vector(4840, 16),
11375 => conv_std_logic_vector(4884, 16),
11376 => conv_std_logic_vector(4928, 16),
11377 => conv_std_logic_vector(4972, 16),
11378 => conv_std_logic_vector(5016, 16),
11379 => conv_std_logic_vector(5060, 16),
11380 => conv_std_logic_vector(5104, 16),
11381 => conv_std_logic_vector(5148, 16),
11382 => conv_std_logic_vector(5192, 16),
11383 => conv_std_logic_vector(5236, 16),
11384 => conv_std_logic_vector(5280, 16),
11385 => conv_std_logic_vector(5324, 16),
11386 => conv_std_logic_vector(5368, 16),
11387 => conv_std_logic_vector(5412, 16),
11388 => conv_std_logic_vector(5456, 16),
11389 => conv_std_logic_vector(5500, 16),
11390 => conv_std_logic_vector(5544, 16),
11391 => conv_std_logic_vector(5588, 16),
11392 => conv_std_logic_vector(5632, 16),
11393 => conv_std_logic_vector(5676, 16),
11394 => conv_std_logic_vector(5720, 16),
11395 => conv_std_logic_vector(5764, 16),
11396 => conv_std_logic_vector(5808, 16),
11397 => conv_std_logic_vector(5852, 16),
11398 => conv_std_logic_vector(5896, 16),
11399 => conv_std_logic_vector(5940, 16),
11400 => conv_std_logic_vector(5984, 16),
11401 => conv_std_logic_vector(6028, 16),
11402 => conv_std_logic_vector(6072, 16),
11403 => conv_std_logic_vector(6116, 16),
11404 => conv_std_logic_vector(6160, 16),
11405 => conv_std_logic_vector(6204, 16),
11406 => conv_std_logic_vector(6248, 16),
11407 => conv_std_logic_vector(6292, 16),
11408 => conv_std_logic_vector(6336, 16),
11409 => conv_std_logic_vector(6380, 16),
11410 => conv_std_logic_vector(6424, 16),
11411 => conv_std_logic_vector(6468, 16),
11412 => conv_std_logic_vector(6512, 16),
11413 => conv_std_logic_vector(6556, 16),
11414 => conv_std_logic_vector(6600, 16),
11415 => conv_std_logic_vector(6644, 16),
11416 => conv_std_logic_vector(6688, 16),
11417 => conv_std_logic_vector(6732, 16),
11418 => conv_std_logic_vector(6776, 16),
11419 => conv_std_logic_vector(6820, 16),
11420 => conv_std_logic_vector(6864, 16),
11421 => conv_std_logic_vector(6908, 16),
11422 => conv_std_logic_vector(6952, 16),
11423 => conv_std_logic_vector(6996, 16),
11424 => conv_std_logic_vector(7040, 16),
11425 => conv_std_logic_vector(7084, 16),
11426 => conv_std_logic_vector(7128, 16),
11427 => conv_std_logic_vector(7172, 16),
11428 => conv_std_logic_vector(7216, 16),
11429 => conv_std_logic_vector(7260, 16),
11430 => conv_std_logic_vector(7304, 16),
11431 => conv_std_logic_vector(7348, 16),
11432 => conv_std_logic_vector(7392, 16),
11433 => conv_std_logic_vector(7436, 16),
11434 => conv_std_logic_vector(7480, 16),
11435 => conv_std_logic_vector(7524, 16),
11436 => conv_std_logic_vector(7568, 16),
11437 => conv_std_logic_vector(7612, 16),
11438 => conv_std_logic_vector(7656, 16),
11439 => conv_std_logic_vector(7700, 16),
11440 => conv_std_logic_vector(7744, 16),
11441 => conv_std_logic_vector(7788, 16),
11442 => conv_std_logic_vector(7832, 16),
11443 => conv_std_logic_vector(7876, 16),
11444 => conv_std_logic_vector(7920, 16),
11445 => conv_std_logic_vector(7964, 16),
11446 => conv_std_logic_vector(8008, 16),
11447 => conv_std_logic_vector(8052, 16),
11448 => conv_std_logic_vector(8096, 16),
11449 => conv_std_logic_vector(8140, 16),
11450 => conv_std_logic_vector(8184, 16),
11451 => conv_std_logic_vector(8228, 16),
11452 => conv_std_logic_vector(8272, 16),
11453 => conv_std_logic_vector(8316, 16),
11454 => conv_std_logic_vector(8360, 16),
11455 => conv_std_logic_vector(8404, 16),
11456 => conv_std_logic_vector(8448, 16),
11457 => conv_std_logic_vector(8492, 16),
11458 => conv_std_logic_vector(8536, 16),
11459 => conv_std_logic_vector(8580, 16),
11460 => conv_std_logic_vector(8624, 16),
11461 => conv_std_logic_vector(8668, 16),
11462 => conv_std_logic_vector(8712, 16),
11463 => conv_std_logic_vector(8756, 16),
11464 => conv_std_logic_vector(8800, 16),
11465 => conv_std_logic_vector(8844, 16),
11466 => conv_std_logic_vector(8888, 16),
11467 => conv_std_logic_vector(8932, 16),
11468 => conv_std_logic_vector(8976, 16),
11469 => conv_std_logic_vector(9020, 16),
11470 => conv_std_logic_vector(9064, 16),
11471 => conv_std_logic_vector(9108, 16),
11472 => conv_std_logic_vector(9152, 16),
11473 => conv_std_logic_vector(9196, 16),
11474 => conv_std_logic_vector(9240, 16),
11475 => conv_std_logic_vector(9284, 16),
11476 => conv_std_logic_vector(9328, 16),
11477 => conv_std_logic_vector(9372, 16),
11478 => conv_std_logic_vector(9416, 16),
11479 => conv_std_logic_vector(9460, 16),
11480 => conv_std_logic_vector(9504, 16),
11481 => conv_std_logic_vector(9548, 16),
11482 => conv_std_logic_vector(9592, 16),
11483 => conv_std_logic_vector(9636, 16),
11484 => conv_std_logic_vector(9680, 16),
11485 => conv_std_logic_vector(9724, 16),
11486 => conv_std_logic_vector(9768, 16),
11487 => conv_std_logic_vector(9812, 16),
11488 => conv_std_logic_vector(9856, 16),
11489 => conv_std_logic_vector(9900, 16),
11490 => conv_std_logic_vector(9944, 16),
11491 => conv_std_logic_vector(9988, 16),
11492 => conv_std_logic_vector(10032, 16),
11493 => conv_std_logic_vector(10076, 16),
11494 => conv_std_logic_vector(10120, 16),
11495 => conv_std_logic_vector(10164, 16),
11496 => conv_std_logic_vector(10208, 16),
11497 => conv_std_logic_vector(10252, 16),
11498 => conv_std_logic_vector(10296, 16),
11499 => conv_std_logic_vector(10340, 16),
11500 => conv_std_logic_vector(10384, 16),
11501 => conv_std_logic_vector(10428, 16),
11502 => conv_std_logic_vector(10472, 16),
11503 => conv_std_logic_vector(10516, 16),
11504 => conv_std_logic_vector(10560, 16),
11505 => conv_std_logic_vector(10604, 16),
11506 => conv_std_logic_vector(10648, 16),
11507 => conv_std_logic_vector(10692, 16),
11508 => conv_std_logic_vector(10736, 16),
11509 => conv_std_logic_vector(10780, 16),
11510 => conv_std_logic_vector(10824, 16),
11511 => conv_std_logic_vector(10868, 16),
11512 => conv_std_logic_vector(10912, 16),
11513 => conv_std_logic_vector(10956, 16),
11514 => conv_std_logic_vector(11000, 16),
11515 => conv_std_logic_vector(11044, 16),
11516 => conv_std_logic_vector(11088, 16),
11517 => conv_std_logic_vector(11132, 16),
11518 => conv_std_logic_vector(11176, 16),
11519 => conv_std_logic_vector(11220, 16),
11520 => conv_std_logic_vector(0, 16),
11521 => conv_std_logic_vector(45, 16),
11522 => conv_std_logic_vector(90, 16),
11523 => conv_std_logic_vector(135, 16),
11524 => conv_std_logic_vector(180, 16),
11525 => conv_std_logic_vector(225, 16),
11526 => conv_std_logic_vector(270, 16),
11527 => conv_std_logic_vector(315, 16),
11528 => conv_std_logic_vector(360, 16),
11529 => conv_std_logic_vector(405, 16),
11530 => conv_std_logic_vector(450, 16),
11531 => conv_std_logic_vector(495, 16),
11532 => conv_std_logic_vector(540, 16),
11533 => conv_std_logic_vector(585, 16),
11534 => conv_std_logic_vector(630, 16),
11535 => conv_std_logic_vector(675, 16),
11536 => conv_std_logic_vector(720, 16),
11537 => conv_std_logic_vector(765, 16),
11538 => conv_std_logic_vector(810, 16),
11539 => conv_std_logic_vector(855, 16),
11540 => conv_std_logic_vector(900, 16),
11541 => conv_std_logic_vector(945, 16),
11542 => conv_std_logic_vector(990, 16),
11543 => conv_std_logic_vector(1035, 16),
11544 => conv_std_logic_vector(1080, 16),
11545 => conv_std_logic_vector(1125, 16),
11546 => conv_std_logic_vector(1170, 16),
11547 => conv_std_logic_vector(1215, 16),
11548 => conv_std_logic_vector(1260, 16),
11549 => conv_std_logic_vector(1305, 16),
11550 => conv_std_logic_vector(1350, 16),
11551 => conv_std_logic_vector(1395, 16),
11552 => conv_std_logic_vector(1440, 16),
11553 => conv_std_logic_vector(1485, 16),
11554 => conv_std_logic_vector(1530, 16),
11555 => conv_std_logic_vector(1575, 16),
11556 => conv_std_logic_vector(1620, 16),
11557 => conv_std_logic_vector(1665, 16),
11558 => conv_std_logic_vector(1710, 16),
11559 => conv_std_logic_vector(1755, 16),
11560 => conv_std_logic_vector(1800, 16),
11561 => conv_std_logic_vector(1845, 16),
11562 => conv_std_logic_vector(1890, 16),
11563 => conv_std_logic_vector(1935, 16),
11564 => conv_std_logic_vector(1980, 16),
11565 => conv_std_logic_vector(2025, 16),
11566 => conv_std_logic_vector(2070, 16),
11567 => conv_std_logic_vector(2115, 16),
11568 => conv_std_logic_vector(2160, 16),
11569 => conv_std_logic_vector(2205, 16),
11570 => conv_std_logic_vector(2250, 16),
11571 => conv_std_logic_vector(2295, 16),
11572 => conv_std_logic_vector(2340, 16),
11573 => conv_std_logic_vector(2385, 16),
11574 => conv_std_logic_vector(2430, 16),
11575 => conv_std_logic_vector(2475, 16),
11576 => conv_std_logic_vector(2520, 16),
11577 => conv_std_logic_vector(2565, 16),
11578 => conv_std_logic_vector(2610, 16),
11579 => conv_std_logic_vector(2655, 16),
11580 => conv_std_logic_vector(2700, 16),
11581 => conv_std_logic_vector(2745, 16),
11582 => conv_std_logic_vector(2790, 16),
11583 => conv_std_logic_vector(2835, 16),
11584 => conv_std_logic_vector(2880, 16),
11585 => conv_std_logic_vector(2925, 16),
11586 => conv_std_logic_vector(2970, 16),
11587 => conv_std_logic_vector(3015, 16),
11588 => conv_std_logic_vector(3060, 16),
11589 => conv_std_logic_vector(3105, 16),
11590 => conv_std_logic_vector(3150, 16),
11591 => conv_std_logic_vector(3195, 16),
11592 => conv_std_logic_vector(3240, 16),
11593 => conv_std_logic_vector(3285, 16),
11594 => conv_std_logic_vector(3330, 16),
11595 => conv_std_logic_vector(3375, 16),
11596 => conv_std_logic_vector(3420, 16),
11597 => conv_std_logic_vector(3465, 16),
11598 => conv_std_logic_vector(3510, 16),
11599 => conv_std_logic_vector(3555, 16),
11600 => conv_std_logic_vector(3600, 16),
11601 => conv_std_logic_vector(3645, 16),
11602 => conv_std_logic_vector(3690, 16),
11603 => conv_std_logic_vector(3735, 16),
11604 => conv_std_logic_vector(3780, 16),
11605 => conv_std_logic_vector(3825, 16),
11606 => conv_std_logic_vector(3870, 16),
11607 => conv_std_logic_vector(3915, 16),
11608 => conv_std_logic_vector(3960, 16),
11609 => conv_std_logic_vector(4005, 16),
11610 => conv_std_logic_vector(4050, 16),
11611 => conv_std_logic_vector(4095, 16),
11612 => conv_std_logic_vector(4140, 16),
11613 => conv_std_logic_vector(4185, 16),
11614 => conv_std_logic_vector(4230, 16),
11615 => conv_std_logic_vector(4275, 16),
11616 => conv_std_logic_vector(4320, 16),
11617 => conv_std_logic_vector(4365, 16),
11618 => conv_std_logic_vector(4410, 16),
11619 => conv_std_logic_vector(4455, 16),
11620 => conv_std_logic_vector(4500, 16),
11621 => conv_std_logic_vector(4545, 16),
11622 => conv_std_logic_vector(4590, 16),
11623 => conv_std_logic_vector(4635, 16),
11624 => conv_std_logic_vector(4680, 16),
11625 => conv_std_logic_vector(4725, 16),
11626 => conv_std_logic_vector(4770, 16),
11627 => conv_std_logic_vector(4815, 16),
11628 => conv_std_logic_vector(4860, 16),
11629 => conv_std_logic_vector(4905, 16),
11630 => conv_std_logic_vector(4950, 16),
11631 => conv_std_logic_vector(4995, 16),
11632 => conv_std_logic_vector(5040, 16),
11633 => conv_std_logic_vector(5085, 16),
11634 => conv_std_logic_vector(5130, 16),
11635 => conv_std_logic_vector(5175, 16),
11636 => conv_std_logic_vector(5220, 16),
11637 => conv_std_logic_vector(5265, 16),
11638 => conv_std_logic_vector(5310, 16),
11639 => conv_std_logic_vector(5355, 16),
11640 => conv_std_logic_vector(5400, 16),
11641 => conv_std_logic_vector(5445, 16),
11642 => conv_std_logic_vector(5490, 16),
11643 => conv_std_logic_vector(5535, 16),
11644 => conv_std_logic_vector(5580, 16),
11645 => conv_std_logic_vector(5625, 16),
11646 => conv_std_logic_vector(5670, 16),
11647 => conv_std_logic_vector(5715, 16),
11648 => conv_std_logic_vector(5760, 16),
11649 => conv_std_logic_vector(5805, 16),
11650 => conv_std_logic_vector(5850, 16),
11651 => conv_std_logic_vector(5895, 16),
11652 => conv_std_logic_vector(5940, 16),
11653 => conv_std_logic_vector(5985, 16),
11654 => conv_std_logic_vector(6030, 16),
11655 => conv_std_logic_vector(6075, 16),
11656 => conv_std_logic_vector(6120, 16),
11657 => conv_std_logic_vector(6165, 16),
11658 => conv_std_logic_vector(6210, 16),
11659 => conv_std_logic_vector(6255, 16),
11660 => conv_std_logic_vector(6300, 16),
11661 => conv_std_logic_vector(6345, 16),
11662 => conv_std_logic_vector(6390, 16),
11663 => conv_std_logic_vector(6435, 16),
11664 => conv_std_logic_vector(6480, 16),
11665 => conv_std_logic_vector(6525, 16),
11666 => conv_std_logic_vector(6570, 16),
11667 => conv_std_logic_vector(6615, 16),
11668 => conv_std_logic_vector(6660, 16),
11669 => conv_std_logic_vector(6705, 16),
11670 => conv_std_logic_vector(6750, 16),
11671 => conv_std_logic_vector(6795, 16),
11672 => conv_std_logic_vector(6840, 16),
11673 => conv_std_logic_vector(6885, 16),
11674 => conv_std_logic_vector(6930, 16),
11675 => conv_std_logic_vector(6975, 16),
11676 => conv_std_logic_vector(7020, 16),
11677 => conv_std_logic_vector(7065, 16),
11678 => conv_std_logic_vector(7110, 16),
11679 => conv_std_logic_vector(7155, 16),
11680 => conv_std_logic_vector(7200, 16),
11681 => conv_std_logic_vector(7245, 16),
11682 => conv_std_logic_vector(7290, 16),
11683 => conv_std_logic_vector(7335, 16),
11684 => conv_std_logic_vector(7380, 16),
11685 => conv_std_logic_vector(7425, 16),
11686 => conv_std_logic_vector(7470, 16),
11687 => conv_std_logic_vector(7515, 16),
11688 => conv_std_logic_vector(7560, 16),
11689 => conv_std_logic_vector(7605, 16),
11690 => conv_std_logic_vector(7650, 16),
11691 => conv_std_logic_vector(7695, 16),
11692 => conv_std_logic_vector(7740, 16),
11693 => conv_std_logic_vector(7785, 16),
11694 => conv_std_logic_vector(7830, 16),
11695 => conv_std_logic_vector(7875, 16),
11696 => conv_std_logic_vector(7920, 16),
11697 => conv_std_logic_vector(7965, 16),
11698 => conv_std_logic_vector(8010, 16),
11699 => conv_std_logic_vector(8055, 16),
11700 => conv_std_logic_vector(8100, 16),
11701 => conv_std_logic_vector(8145, 16),
11702 => conv_std_logic_vector(8190, 16),
11703 => conv_std_logic_vector(8235, 16),
11704 => conv_std_logic_vector(8280, 16),
11705 => conv_std_logic_vector(8325, 16),
11706 => conv_std_logic_vector(8370, 16),
11707 => conv_std_logic_vector(8415, 16),
11708 => conv_std_logic_vector(8460, 16),
11709 => conv_std_logic_vector(8505, 16),
11710 => conv_std_logic_vector(8550, 16),
11711 => conv_std_logic_vector(8595, 16),
11712 => conv_std_logic_vector(8640, 16),
11713 => conv_std_logic_vector(8685, 16),
11714 => conv_std_logic_vector(8730, 16),
11715 => conv_std_logic_vector(8775, 16),
11716 => conv_std_logic_vector(8820, 16),
11717 => conv_std_logic_vector(8865, 16),
11718 => conv_std_logic_vector(8910, 16),
11719 => conv_std_logic_vector(8955, 16),
11720 => conv_std_logic_vector(9000, 16),
11721 => conv_std_logic_vector(9045, 16),
11722 => conv_std_logic_vector(9090, 16),
11723 => conv_std_logic_vector(9135, 16),
11724 => conv_std_logic_vector(9180, 16),
11725 => conv_std_logic_vector(9225, 16),
11726 => conv_std_logic_vector(9270, 16),
11727 => conv_std_logic_vector(9315, 16),
11728 => conv_std_logic_vector(9360, 16),
11729 => conv_std_logic_vector(9405, 16),
11730 => conv_std_logic_vector(9450, 16),
11731 => conv_std_logic_vector(9495, 16),
11732 => conv_std_logic_vector(9540, 16),
11733 => conv_std_logic_vector(9585, 16),
11734 => conv_std_logic_vector(9630, 16),
11735 => conv_std_logic_vector(9675, 16),
11736 => conv_std_logic_vector(9720, 16),
11737 => conv_std_logic_vector(9765, 16),
11738 => conv_std_logic_vector(9810, 16),
11739 => conv_std_logic_vector(9855, 16),
11740 => conv_std_logic_vector(9900, 16),
11741 => conv_std_logic_vector(9945, 16),
11742 => conv_std_logic_vector(9990, 16),
11743 => conv_std_logic_vector(10035, 16),
11744 => conv_std_logic_vector(10080, 16),
11745 => conv_std_logic_vector(10125, 16),
11746 => conv_std_logic_vector(10170, 16),
11747 => conv_std_logic_vector(10215, 16),
11748 => conv_std_logic_vector(10260, 16),
11749 => conv_std_logic_vector(10305, 16),
11750 => conv_std_logic_vector(10350, 16),
11751 => conv_std_logic_vector(10395, 16),
11752 => conv_std_logic_vector(10440, 16),
11753 => conv_std_logic_vector(10485, 16),
11754 => conv_std_logic_vector(10530, 16),
11755 => conv_std_logic_vector(10575, 16),
11756 => conv_std_logic_vector(10620, 16),
11757 => conv_std_logic_vector(10665, 16),
11758 => conv_std_logic_vector(10710, 16),
11759 => conv_std_logic_vector(10755, 16),
11760 => conv_std_logic_vector(10800, 16),
11761 => conv_std_logic_vector(10845, 16),
11762 => conv_std_logic_vector(10890, 16),
11763 => conv_std_logic_vector(10935, 16),
11764 => conv_std_logic_vector(10980, 16),
11765 => conv_std_logic_vector(11025, 16),
11766 => conv_std_logic_vector(11070, 16),
11767 => conv_std_logic_vector(11115, 16),
11768 => conv_std_logic_vector(11160, 16),
11769 => conv_std_logic_vector(11205, 16),
11770 => conv_std_logic_vector(11250, 16),
11771 => conv_std_logic_vector(11295, 16),
11772 => conv_std_logic_vector(11340, 16),
11773 => conv_std_logic_vector(11385, 16),
11774 => conv_std_logic_vector(11430, 16),
11775 => conv_std_logic_vector(11475, 16),
11776 => conv_std_logic_vector(0, 16),
11777 => conv_std_logic_vector(46, 16),
11778 => conv_std_logic_vector(92, 16),
11779 => conv_std_logic_vector(138, 16),
11780 => conv_std_logic_vector(184, 16),
11781 => conv_std_logic_vector(230, 16),
11782 => conv_std_logic_vector(276, 16),
11783 => conv_std_logic_vector(322, 16),
11784 => conv_std_logic_vector(368, 16),
11785 => conv_std_logic_vector(414, 16),
11786 => conv_std_logic_vector(460, 16),
11787 => conv_std_logic_vector(506, 16),
11788 => conv_std_logic_vector(552, 16),
11789 => conv_std_logic_vector(598, 16),
11790 => conv_std_logic_vector(644, 16),
11791 => conv_std_logic_vector(690, 16),
11792 => conv_std_logic_vector(736, 16),
11793 => conv_std_logic_vector(782, 16),
11794 => conv_std_logic_vector(828, 16),
11795 => conv_std_logic_vector(874, 16),
11796 => conv_std_logic_vector(920, 16),
11797 => conv_std_logic_vector(966, 16),
11798 => conv_std_logic_vector(1012, 16),
11799 => conv_std_logic_vector(1058, 16),
11800 => conv_std_logic_vector(1104, 16),
11801 => conv_std_logic_vector(1150, 16),
11802 => conv_std_logic_vector(1196, 16),
11803 => conv_std_logic_vector(1242, 16),
11804 => conv_std_logic_vector(1288, 16),
11805 => conv_std_logic_vector(1334, 16),
11806 => conv_std_logic_vector(1380, 16),
11807 => conv_std_logic_vector(1426, 16),
11808 => conv_std_logic_vector(1472, 16),
11809 => conv_std_logic_vector(1518, 16),
11810 => conv_std_logic_vector(1564, 16),
11811 => conv_std_logic_vector(1610, 16),
11812 => conv_std_logic_vector(1656, 16),
11813 => conv_std_logic_vector(1702, 16),
11814 => conv_std_logic_vector(1748, 16),
11815 => conv_std_logic_vector(1794, 16),
11816 => conv_std_logic_vector(1840, 16),
11817 => conv_std_logic_vector(1886, 16),
11818 => conv_std_logic_vector(1932, 16),
11819 => conv_std_logic_vector(1978, 16),
11820 => conv_std_logic_vector(2024, 16),
11821 => conv_std_logic_vector(2070, 16),
11822 => conv_std_logic_vector(2116, 16),
11823 => conv_std_logic_vector(2162, 16),
11824 => conv_std_logic_vector(2208, 16),
11825 => conv_std_logic_vector(2254, 16),
11826 => conv_std_logic_vector(2300, 16),
11827 => conv_std_logic_vector(2346, 16),
11828 => conv_std_logic_vector(2392, 16),
11829 => conv_std_logic_vector(2438, 16),
11830 => conv_std_logic_vector(2484, 16),
11831 => conv_std_logic_vector(2530, 16),
11832 => conv_std_logic_vector(2576, 16),
11833 => conv_std_logic_vector(2622, 16),
11834 => conv_std_logic_vector(2668, 16),
11835 => conv_std_logic_vector(2714, 16),
11836 => conv_std_logic_vector(2760, 16),
11837 => conv_std_logic_vector(2806, 16),
11838 => conv_std_logic_vector(2852, 16),
11839 => conv_std_logic_vector(2898, 16),
11840 => conv_std_logic_vector(2944, 16),
11841 => conv_std_logic_vector(2990, 16),
11842 => conv_std_logic_vector(3036, 16),
11843 => conv_std_logic_vector(3082, 16),
11844 => conv_std_logic_vector(3128, 16),
11845 => conv_std_logic_vector(3174, 16),
11846 => conv_std_logic_vector(3220, 16),
11847 => conv_std_logic_vector(3266, 16),
11848 => conv_std_logic_vector(3312, 16),
11849 => conv_std_logic_vector(3358, 16),
11850 => conv_std_logic_vector(3404, 16),
11851 => conv_std_logic_vector(3450, 16),
11852 => conv_std_logic_vector(3496, 16),
11853 => conv_std_logic_vector(3542, 16),
11854 => conv_std_logic_vector(3588, 16),
11855 => conv_std_logic_vector(3634, 16),
11856 => conv_std_logic_vector(3680, 16),
11857 => conv_std_logic_vector(3726, 16),
11858 => conv_std_logic_vector(3772, 16),
11859 => conv_std_logic_vector(3818, 16),
11860 => conv_std_logic_vector(3864, 16),
11861 => conv_std_logic_vector(3910, 16),
11862 => conv_std_logic_vector(3956, 16),
11863 => conv_std_logic_vector(4002, 16),
11864 => conv_std_logic_vector(4048, 16),
11865 => conv_std_logic_vector(4094, 16),
11866 => conv_std_logic_vector(4140, 16),
11867 => conv_std_logic_vector(4186, 16),
11868 => conv_std_logic_vector(4232, 16),
11869 => conv_std_logic_vector(4278, 16),
11870 => conv_std_logic_vector(4324, 16),
11871 => conv_std_logic_vector(4370, 16),
11872 => conv_std_logic_vector(4416, 16),
11873 => conv_std_logic_vector(4462, 16),
11874 => conv_std_logic_vector(4508, 16),
11875 => conv_std_logic_vector(4554, 16),
11876 => conv_std_logic_vector(4600, 16),
11877 => conv_std_logic_vector(4646, 16),
11878 => conv_std_logic_vector(4692, 16),
11879 => conv_std_logic_vector(4738, 16),
11880 => conv_std_logic_vector(4784, 16),
11881 => conv_std_logic_vector(4830, 16),
11882 => conv_std_logic_vector(4876, 16),
11883 => conv_std_logic_vector(4922, 16),
11884 => conv_std_logic_vector(4968, 16),
11885 => conv_std_logic_vector(5014, 16),
11886 => conv_std_logic_vector(5060, 16),
11887 => conv_std_logic_vector(5106, 16),
11888 => conv_std_logic_vector(5152, 16),
11889 => conv_std_logic_vector(5198, 16),
11890 => conv_std_logic_vector(5244, 16),
11891 => conv_std_logic_vector(5290, 16),
11892 => conv_std_logic_vector(5336, 16),
11893 => conv_std_logic_vector(5382, 16),
11894 => conv_std_logic_vector(5428, 16),
11895 => conv_std_logic_vector(5474, 16),
11896 => conv_std_logic_vector(5520, 16),
11897 => conv_std_logic_vector(5566, 16),
11898 => conv_std_logic_vector(5612, 16),
11899 => conv_std_logic_vector(5658, 16),
11900 => conv_std_logic_vector(5704, 16),
11901 => conv_std_logic_vector(5750, 16),
11902 => conv_std_logic_vector(5796, 16),
11903 => conv_std_logic_vector(5842, 16),
11904 => conv_std_logic_vector(5888, 16),
11905 => conv_std_logic_vector(5934, 16),
11906 => conv_std_logic_vector(5980, 16),
11907 => conv_std_logic_vector(6026, 16),
11908 => conv_std_logic_vector(6072, 16),
11909 => conv_std_logic_vector(6118, 16),
11910 => conv_std_logic_vector(6164, 16),
11911 => conv_std_logic_vector(6210, 16),
11912 => conv_std_logic_vector(6256, 16),
11913 => conv_std_logic_vector(6302, 16),
11914 => conv_std_logic_vector(6348, 16),
11915 => conv_std_logic_vector(6394, 16),
11916 => conv_std_logic_vector(6440, 16),
11917 => conv_std_logic_vector(6486, 16),
11918 => conv_std_logic_vector(6532, 16),
11919 => conv_std_logic_vector(6578, 16),
11920 => conv_std_logic_vector(6624, 16),
11921 => conv_std_logic_vector(6670, 16),
11922 => conv_std_logic_vector(6716, 16),
11923 => conv_std_logic_vector(6762, 16),
11924 => conv_std_logic_vector(6808, 16),
11925 => conv_std_logic_vector(6854, 16),
11926 => conv_std_logic_vector(6900, 16),
11927 => conv_std_logic_vector(6946, 16),
11928 => conv_std_logic_vector(6992, 16),
11929 => conv_std_logic_vector(7038, 16),
11930 => conv_std_logic_vector(7084, 16),
11931 => conv_std_logic_vector(7130, 16),
11932 => conv_std_logic_vector(7176, 16),
11933 => conv_std_logic_vector(7222, 16),
11934 => conv_std_logic_vector(7268, 16),
11935 => conv_std_logic_vector(7314, 16),
11936 => conv_std_logic_vector(7360, 16),
11937 => conv_std_logic_vector(7406, 16),
11938 => conv_std_logic_vector(7452, 16),
11939 => conv_std_logic_vector(7498, 16),
11940 => conv_std_logic_vector(7544, 16),
11941 => conv_std_logic_vector(7590, 16),
11942 => conv_std_logic_vector(7636, 16),
11943 => conv_std_logic_vector(7682, 16),
11944 => conv_std_logic_vector(7728, 16),
11945 => conv_std_logic_vector(7774, 16),
11946 => conv_std_logic_vector(7820, 16),
11947 => conv_std_logic_vector(7866, 16),
11948 => conv_std_logic_vector(7912, 16),
11949 => conv_std_logic_vector(7958, 16),
11950 => conv_std_logic_vector(8004, 16),
11951 => conv_std_logic_vector(8050, 16),
11952 => conv_std_logic_vector(8096, 16),
11953 => conv_std_logic_vector(8142, 16),
11954 => conv_std_logic_vector(8188, 16),
11955 => conv_std_logic_vector(8234, 16),
11956 => conv_std_logic_vector(8280, 16),
11957 => conv_std_logic_vector(8326, 16),
11958 => conv_std_logic_vector(8372, 16),
11959 => conv_std_logic_vector(8418, 16),
11960 => conv_std_logic_vector(8464, 16),
11961 => conv_std_logic_vector(8510, 16),
11962 => conv_std_logic_vector(8556, 16),
11963 => conv_std_logic_vector(8602, 16),
11964 => conv_std_logic_vector(8648, 16),
11965 => conv_std_logic_vector(8694, 16),
11966 => conv_std_logic_vector(8740, 16),
11967 => conv_std_logic_vector(8786, 16),
11968 => conv_std_logic_vector(8832, 16),
11969 => conv_std_logic_vector(8878, 16),
11970 => conv_std_logic_vector(8924, 16),
11971 => conv_std_logic_vector(8970, 16),
11972 => conv_std_logic_vector(9016, 16),
11973 => conv_std_logic_vector(9062, 16),
11974 => conv_std_logic_vector(9108, 16),
11975 => conv_std_logic_vector(9154, 16),
11976 => conv_std_logic_vector(9200, 16),
11977 => conv_std_logic_vector(9246, 16),
11978 => conv_std_logic_vector(9292, 16),
11979 => conv_std_logic_vector(9338, 16),
11980 => conv_std_logic_vector(9384, 16),
11981 => conv_std_logic_vector(9430, 16),
11982 => conv_std_logic_vector(9476, 16),
11983 => conv_std_logic_vector(9522, 16),
11984 => conv_std_logic_vector(9568, 16),
11985 => conv_std_logic_vector(9614, 16),
11986 => conv_std_logic_vector(9660, 16),
11987 => conv_std_logic_vector(9706, 16),
11988 => conv_std_logic_vector(9752, 16),
11989 => conv_std_logic_vector(9798, 16),
11990 => conv_std_logic_vector(9844, 16),
11991 => conv_std_logic_vector(9890, 16),
11992 => conv_std_logic_vector(9936, 16),
11993 => conv_std_logic_vector(9982, 16),
11994 => conv_std_logic_vector(10028, 16),
11995 => conv_std_logic_vector(10074, 16),
11996 => conv_std_logic_vector(10120, 16),
11997 => conv_std_logic_vector(10166, 16),
11998 => conv_std_logic_vector(10212, 16),
11999 => conv_std_logic_vector(10258, 16),
12000 => conv_std_logic_vector(10304, 16),
12001 => conv_std_logic_vector(10350, 16),
12002 => conv_std_logic_vector(10396, 16),
12003 => conv_std_logic_vector(10442, 16),
12004 => conv_std_logic_vector(10488, 16),
12005 => conv_std_logic_vector(10534, 16),
12006 => conv_std_logic_vector(10580, 16),
12007 => conv_std_logic_vector(10626, 16),
12008 => conv_std_logic_vector(10672, 16),
12009 => conv_std_logic_vector(10718, 16),
12010 => conv_std_logic_vector(10764, 16),
12011 => conv_std_logic_vector(10810, 16),
12012 => conv_std_logic_vector(10856, 16),
12013 => conv_std_logic_vector(10902, 16),
12014 => conv_std_logic_vector(10948, 16),
12015 => conv_std_logic_vector(10994, 16),
12016 => conv_std_logic_vector(11040, 16),
12017 => conv_std_logic_vector(11086, 16),
12018 => conv_std_logic_vector(11132, 16),
12019 => conv_std_logic_vector(11178, 16),
12020 => conv_std_logic_vector(11224, 16),
12021 => conv_std_logic_vector(11270, 16),
12022 => conv_std_logic_vector(11316, 16),
12023 => conv_std_logic_vector(11362, 16),
12024 => conv_std_logic_vector(11408, 16),
12025 => conv_std_logic_vector(11454, 16),
12026 => conv_std_logic_vector(11500, 16),
12027 => conv_std_logic_vector(11546, 16),
12028 => conv_std_logic_vector(11592, 16),
12029 => conv_std_logic_vector(11638, 16),
12030 => conv_std_logic_vector(11684, 16),
12031 => conv_std_logic_vector(11730, 16),
12032 => conv_std_logic_vector(0, 16),
12033 => conv_std_logic_vector(47, 16),
12034 => conv_std_logic_vector(94, 16),
12035 => conv_std_logic_vector(141, 16),
12036 => conv_std_logic_vector(188, 16),
12037 => conv_std_logic_vector(235, 16),
12038 => conv_std_logic_vector(282, 16),
12039 => conv_std_logic_vector(329, 16),
12040 => conv_std_logic_vector(376, 16),
12041 => conv_std_logic_vector(423, 16),
12042 => conv_std_logic_vector(470, 16),
12043 => conv_std_logic_vector(517, 16),
12044 => conv_std_logic_vector(564, 16),
12045 => conv_std_logic_vector(611, 16),
12046 => conv_std_logic_vector(658, 16),
12047 => conv_std_logic_vector(705, 16),
12048 => conv_std_logic_vector(752, 16),
12049 => conv_std_logic_vector(799, 16),
12050 => conv_std_logic_vector(846, 16),
12051 => conv_std_logic_vector(893, 16),
12052 => conv_std_logic_vector(940, 16),
12053 => conv_std_logic_vector(987, 16),
12054 => conv_std_logic_vector(1034, 16),
12055 => conv_std_logic_vector(1081, 16),
12056 => conv_std_logic_vector(1128, 16),
12057 => conv_std_logic_vector(1175, 16),
12058 => conv_std_logic_vector(1222, 16),
12059 => conv_std_logic_vector(1269, 16),
12060 => conv_std_logic_vector(1316, 16),
12061 => conv_std_logic_vector(1363, 16),
12062 => conv_std_logic_vector(1410, 16),
12063 => conv_std_logic_vector(1457, 16),
12064 => conv_std_logic_vector(1504, 16),
12065 => conv_std_logic_vector(1551, 16),
12066 => conv_std_logic_vector(1598, 16),
12067 => conv_std_logic_vector(1645, 16),
12068 => conv_std_logic_vector(1692, 16),
12069 => conv_std_logic_vector(1739, 16),
12070 => conv_std_logic_vector(1786, 16),
12071 => conv_std_logic_vector(1833, 16),
12072 => conv_std_logic_vector(1880, 16),
12073 => conv_std_logic_vector(1927, 16),
12074 => conv_std_logic_vector(1974, 16),
12075 => conv_std_logic_vector(2021, 16),
12076 => conv_std_logic_vector(2068, 16),
12077 => conv_std_logic_vector(2115, 16),
12078 => conv_std_logic_vector(2162, 16),
12079 => conv_std_logic_vector(2209, 16),
12080 => conv_std_logic_vector(2256, 16),
12081 => conv_std_logic_vector(2303, 16),
12082 => conv_std_logic_vector(2350, 16),
12083 => conv_std_logic_vector(2397, 16),
12084 => conv_std_logic_vector(2444, 16),
12085 => conv_std_logic_vector(2491, 16),
12086 => conv_std_logic_vector(2538, 16),
12087 => conv_std_logic_vector(2585, 16),
12088 => conv_std_logic_vector(2632, 16),
12089 => conv_std_logic_vector(2679, 16),
12090 => conv_std_logic_vector(2726, 16),
12091 => conv_std_logic_vector(2773, 16),
12092 => conv_std_logic_vector(2820, 16),
12093 => conv_std_logic_vector(2867, 16),
12094 => conv_std_logic_vector(2914, 16),
12095 => conv_std_logic_vector(2961, 16),
12096 => conv_std_logic_vector(3008, 16),
12097 => conv_std_logic_vector(3055, 16),
12098 => conv_std_logic_vector(3102, 16),
12099 => conv_std_logic_vector(3149, 16),
12100 => conv_std_logic_vector(3196, 16),
12101 => conv_std_logic_vector(3243, 16),
12102 => conv_std_logic_vector(3290, 16),
12103 => conv_std_logic_vector(3337, 16),
12104 => conv_std_logic_vector(3384, 16),
12105 => conv_std_logic_vector(3431, 16),
12106 => conv_std_logic_vector(3478, 16),
12107 => conv_std_logic_vector(3525, 16),
12108 => conv_std_logic_vector(3572, 16),
12109 => conv_std_logic_vector(3619, 16),
12110 => conv_std_logic_vector(3666, 16),
12111 => conv_std_logic_vector(3713, 16),
12112 => conv_std_logic_vector(3760, 16),
12113 => conv_std_logic_vector(3807, 16),
12114 => conv_std_logic_vector(3854, 16),
12115 => conv_std_logic_vector(3901, 16),
12116 => conv_std_logic_vector(3948, 16),
12117 => conv_std_logic_vector(3995, 16),
12118 => conv_std_logic_vector(4042, 16),
12119 => conv_std_logic_vector(4089, 16),
12120 => conv_std_logic_vector(4136, 16),
12121 => conv_std_logic_vector(4183, 16),
12122 => conv_std_logic_vector(4230, 16),
12123 => conv_std_logic_vector(4277, 16),
12124 => conv_std_logic_vector(4324, 16),
12125 => conv_std_logic_vector(4371, 16),
12126 => conv_std_logic_vector(4418, 16),
12127 => conv_std_logic_vector(4465, 16),
12128 => conv_std_logic_vector(4512, 16),
12129 => conv_std_logic_vector(4559, 16),
12130 => conv_std_logic_vector(4606, 16),
12131 => conv_std_logic_vector(4653, 16),
12132 => conv_std_logic_vector(4700, 16),
12133 => conv_std_logic_vector(4747, 16),
12134 => conv_std_logic_vector(4794, 16),
12135 => conv_std_logic_vector(4841, 16),
12136 => conv_std_logic_vector(4888, 16),
12137 => conv_std_logic_vector(4935, 16),
12138 => conv_std_logic_vector(4982, 16),
12139 => conv_std_logic_vector(5029, 16),
12140 => conv_std_logic_vector(5076, 16),
12141 => conv_std_logic_vector(5123, 16),
12142 => conv_std_logic_vector(5170, 16),
12143 => conv_std_logic_vector(5217, 16),
12144 => conv_std_logic_vector(5264, 16),
12145 => conv_std_logic_vector(5311, 16),
12146 => conv_std_logic_vector(5358, 16),
12147 => conv_std_logic_vector(5405, 16),
12148 => conv_std_logic_vector(5452, 16),
12149 => conv_std_logic_vector(5499, 16),
12150 => conv_std_logic_vector(5546, 16),
12151 => conv_std_logic_vector(5593, 16),
12152 => conv_std_logic_vector(5640, 16),
12153 => conv_std_logic_vector(5687, 16),
12154 => conv_std_logic_vector(5734, 16),
12155 => conv_std_logic_vector(5781, 16),
12156 => conv_std_logic_vector(5828, 16),
12157 => conv_std_logic_vector(5875, 16),
12158 => conv_std_logic_vector(5922, 16),
12159 => conv_std_logic_vector(5969, 16),
12160 => conv_std_logic_vector(6016, 16),
12161 => conv_std_logic_vector(6063, 16),
12162 => conv_std_logic_vector(6110, 16),
12163 => conv_std_logic_vector(6157, 16),
12164 => conv_std_logic_vector(6204, 16),
12165 => conv_std_logic_vector(6251, 16),
12166 => conv_std_logic_vector(6298, 16),
12167 => conv_std_logic_vector(6345, 16),
12168 => conv_std_logic_vector(6392, 16),
12169 => conv_std_logic_vector(6439, 16),
12170 => conv_std_logic_vector(6486, 16),
12171 => conv_std_logic_vector(6533, 16),
12172 => conv_std_logic_vector(6580, 16),
12173 => conv_std_logic_vector(6627, 16),
12174 => conv_std_logic_vector(6674, 16),
12175 => conv_std_logic_vector(6721, 16),
12176 => conv_std_logic_vector(6768, 16),
12177 => conv_std_logic_vector(6815, 16),
12178 => conv_std_logic_vector(6862, 16),
12179 => conv_std_logic_vector(6909, 16),
12180 => conv_std_logic_vector(6956, 16),
12181 => conv_std_logic_vector(7003, 16),
12182 => conv_std_logic_vector(7050, 16),
12183 => conv_std_logic_vector(7097, 16),
12184 => conv_std_logic_vector(7144, 16),
12185 => conv_std_logic_vector(7191, 16),
12186 => conv_std_logic_vector(7238, 16),
12187 => conv_std_logic_vector(7285, 16),
12188 => conv_std_logic_vector(7332, 16),
12189 => conv_std_logic_vector(7379, 16),
12190 => conv_std_logic_vector(7426, 16),
12191 => conv_std_logic_vector(7473, 16),
12192 => conv_std_logic_vector(7520, 16),
12193 => conv_std_logic_vector(7567, 16),
12194 => conv_std_logic_vector(7614, 16),
12195 => conv_std_logic_vector(7661, 16),
12196 => conv_std_logic_vector(7708, 16),
12197 => conv_std_logic_vector(7755, 16),
12198 => conv_std_logic_vector(7802, 16),
12199 => conv_std_logic_vector(7849, 16),
12200 => conv_std_logic_vector(7896, 16),
12201 => conv_std_logic_vector(7943, 16),
12202 => conv_std_logic_vector(7990, 16),
12203 => conv_std_logic_vector(8037, 16),
12204 => conv_std_logic_vector(8084, 16),
12205 => conv_std_logic_vector(8131, 16),
12206 => conv_std_logic_vector(8178, 16),
12207 => conv_std_logic_vector(8225, 16),
12208 => conv_std_logic_vector(8272, 16),
12209 => conv_std_logic_vector(8319, 16),
12210 => conv_std_logic_vector(8366, 16),
12211 => conv_std_logic_vector(8413, 16),
12212 => conv_std_logic_vector(8460, 16),
12213 => conv_std_logic_vector(8507, 16),
12214 => conv_std_logic_vector(8554, 16),
12215 => conv_std_logic_vector(8601, 16),
12216 => conv_std_logic_vector(8648, 16),
12217 => conv_std_logic_vector(8695, 16),
12218 => conv_std_logic_vector(8742, 16),
12219 => conv_std_logic_vector(8789, 16),
12220 => conv_std_logic_vector(8836, 16),
12221 => conv_std_logic_vector(8883, 16),
12222 => conv_std_logic_vector(8930, 16),
12223 => conv_std_logic_vector(8977, 16),
12224 => conv_std_logic_vector(9024, 16),
12225 => conv_std_logic_vector(9071, 16),
12226 => conv_std_logic_vector(9118, 16),
12227 => conv_std_logic_vector(9165, 16),
12228 => conv_std_logic_vector(9212, 16),
12229 => conv_std_logic_vector(9259, 16),
12230 => conv_std_logic_vector(9306, 16),
12231 => conv_std_logic_vector(9353, 16),
12232 => conv_std_logic_vector(9400, 16),
12233 => conv_std_logic_vector(9447, 16),
12234 => conv_std_logic_vector(9494, 16),
12235 => conv_std_logic_vector(9541, 16),
12236 => conv_std_logic_vector(9588, 16),
12237 => conv_std_logic_vector(9635, 16),
12238 => conv_std_logic_vector(9682, 16),
12239 => conv_std_logic_vector(9729, 16),
12240 => conv_std_logic_vector(9776, 16),
12241 => conv_std_logic_vector(9823, 16),
12242 => conv_std_logic_vector(9870, 16),
12243 => conv_std_logic_vector(9917, 16),
12244 => conv_std_logic_vector(9964, 16),
12245 => conv_std_logic_vector(10011, 16),
12246 => conv_std_logic_vector(10058, 16),
12247 => conv_std_logic_vector(10105, 16),
12248 => conv_std_logic_vector(10152, 16),
12249 => conv_std_logic_vector(10199, 16),
12250 => conv_std_logic_vector(10246, 16),
12251 => conv_std_logic_vector(10293, 16),
12252 => conv_std_logic_vector(10340, 16),
12253 => conv_std_logic_vector(10387, 16),
12254 => conv_std_logic_vector(10434, 16),
12255 => conv_std_logic_vector(10481, 16),
12256 => conv_std_logic_vector(10528, 16),
12257 => conv_std_logic_vector(10575, 16),
12258 => conv_std_logic_vector(10622, 16),
12259 => conv_std_logic_vector(10669, 16),
12260 => conv_std_logic_vector(10716, 16),
12261 => conv_std_logic_vector(10763, 16),
12262 => conv_std_logic_vector(10810, 16),
12263 => conv_std_logic_vector(10857, 16),
12264 => conv_std_logic_vector(10904, 16),
12265 => conv_std_logic_vector(10951, 16),
12266 => conv_std_logic_vector(10998, 16),
12267 => conv_std_logic_vector(11045, 16),
12268 => conv_std_logic_vector(11092, 16),
12269 => conv_std_logic_vector(11139, 16),
12270 => conv_std_logic_vector(11186, 16),
12271 => conv_std_logic_vector(11233, 16),
12272 => conv_std_logic_vector(11280, 16),
12273 => conv_std_logic_vector(11327, 16),
12274 => conv_std_logic_vector(11374, 16),
12275 => conv_std_logic_vector(11421, 16),
12276 => conv_std_logic_vector(11468, 16),
12277 => conv_std_logic_vector(11515, 16),
12278 => conv_std_logic_vector(11562, 16),
12279 => conv_std_logic_vector(11609, 16),
12280 => conv_std_logic_vector(11656, 16),
12281 => conv_std_logic_vector(11703, 16),
12282 => conv_std_logic_vector(11750, 16),
12283 => conv_std_logic_vector(11797, 16),
12284 => conv_std_logic_vector(11844, 16),
12285 => conv_std_logic_vector(11891, 16),
12286 => conv_std_logic_vector(11938, 16),
12287 => conv_std_logic_vector(11985, 16),
12288 => conv_std_logic_vector(0, 16),
12289 => conv_std_logic_vector(48, 16),
12290 => conv_std_logic_vector(96, 16),
12291 => conv_std_logic_vector(144, 16),
12292 => conv_std_logic_vector(192, 16),
12293 => conv_std_logic_vector(240, 16),
12294 => conv_std_logic_vector(288, 16),
12295 => conv_std_logic_vector(336, 16),
12296 => conv_std_logic_vector(384, 16),
12297 => conv_std_logic_vector(432, 16),
12298 => conv_std_logic_vector(480, 16),
12299 => conv_std_logic_vector(528, 16),
12300 => conv_std_logic_vector(576, 16),
12301 => conv_std_logic_vector(624, 16),
12302 => conv_std_logic_vector(672, 16),
12303 => conv_std_logic_vector(720, 16),
12304 => conv_std_logic_vector(768, 16),
12305 => conv_std_logic_vector(816, 16),
12306 => conv_std_logic_vector(864, 16),
12307 => conv_std_logic_vector(912, 16),
12308 => conv_std_logic_vector(960, 16),
12309 => conv_std_logic_vector(1008, 16),
12310 => conv_std_logic_vector(1056, 16),
12311 => conv_std_logic_vector(1104, 16),
12312 => conv_std_logic_vector(1152, 16),
12313 => conv_std_logic_vector(1200, 16),
12314 => conv_std_logic_vector(1248, 16),
12315 => conv_std_logic_vector(1296, 16),
12316 => conv_std_logic_vector(1344, 16),
12317 => conv_std_logic_vector(1392, 16),
12318 => conv_std_logic_vector(1440, 16),
12319 => conv_std_logic_vector(1488, 16),
12320 => conv_std_logic_vector(1536, 16),
12321 => conv_std_logic_vector(1584, 16),
12322 => conv_std_logic_vector(1632, 16),
12323 => conv_std_logic_vector(1680, 16),
12324 => conv_std_logic_vector(1728, 16),
12325 => conv_std_logic_vector(1776, 16),
12326 => conv_std_logic_vector(1824, 16),
12327 => conv_std_logic_vector(1872, 16),
12328 => conv_std_logic_vector(1920, 16),
12329 => conv_std_logic_vector(1968, 16),
12330 => conv_std_logic_vector(2016, 16),
12331 => conv_std_logic_vector(2064, 16),
12332 => conv_std_logic_vector(2112, 16),
12333 => conv_std_logic_vector(2160, 16),
12334 => conv_std_logic_vector(2208, 16),
12335 => conv_std_logic_vector(2256, 16),
12336 => conv_std_logic_vector(2304, 16),
12337 => conv_std_logic_vector(2352, 16),
12338 => conv_std_logic_vector(2400, 16),
12339 => conv_std_logic_vector(2448, 16),
12340 => conv_std_logic_vector(2496, 16),
12341 => conv_std_logic_vector(2544, 16),
12342 => conv_std_logic_vector(2592, 16),
12343 => conv_std_logic_vector(2640, 16),
12344 => conv_std_logic_vector(2688, 16),
12345 => conv_std_logic_vector(2736, 16),
12346 => conv_std_logic_vector(2784, 16),
12347 => conv_std_logic_vector(2832, 16),
12348 => conv_std_logic_vector(2880, 16),
12349 => conv_std_logic_vector(2928, 16),
12350 => conv_std_logic_vector(2976, 16),
12351 => conv_std_logic_vector(3024, 16),
12352 => conv_std_logic_vector(3072, 16),
12353 => conv_std_logic_vector(3120, 16),
12354 => conv_std_logic_vector(3168, 16),
12355 => conv_std_logic_vector(3216, 16),
12356 => conv_std_logic_vector(3264, 16),
12357 => conv_std_logic_vector(3312, 16),
12358 => conv_std_logic_vector(3360, 16),
12359 => conv_std_logic_vector(3408, 16),
12360 => conv_std_logic_vector(3456, 16),
12361 => conv_std_logic_vector(3504, 16),
12362 => conv_std_logic_vector(3552, 16),
12363 => conv_std_logic_vector(3600, 16),
12364 => conv_std_logic_vector(3648, 16),
12365 => conv_std_logic_vector(3696, 16),
12366 => conv_std_logic_vector(3744, 16),
12367 => conv_std_logic_vector(3792, 16),
12368 => conv_std_logic_vector(3840, 16),
12369 => conv_std_logic_vector(3888, 16),
12370 => conv_std_logic_vector(3936, 16),
12371 => conv_std_logic_vector(3984, 16),
12372 => conv_std_logic_vector(4032, 16),
12373 => conv_std_logic_vector(4080, 16),
12374 => conv_std_logic_vector(4128, 16),
12375 => conv_std_logic_vector(4176, 16),
12376 => conv_std_logic_vector(4224, 16),
12377 => conv_std_logic_vector(4272, 16),
12378 => conv_std_logic_vector(4320, 16),
12379 => conv_std_logic_vector(4368, 16),
12380 => conv_std_logic_vector(4416, 16),
12381 => conv_std_logic_vector(4464, 16),
12382 => conv_std_logic_vector(4512, 16),
12383 => conv_std_logic_vector(4560, 16),
12384 => conv_std_logic_vector(4608, 16),
12385 => conv_std_logic_vector(4656, 16),
12386 => conv_std_logic_vector(4704, 16),
12387 => conv_std_logic_vector(4752, 16),
12388 => conv_std_logic_vector(4800, 16),
12389 => conv_std_logic_vector(4848, 16),
12390 => conv_std_logic_vector(4896, 16),
12391 => conv_std_logic_vector(4944, 16),
12392 => conv_std_logic_vector(4992, 16),
12393 => conv_std_logic_vector(5040, 16),
12394 => conv_std_logic_vector(5088, 16),
12395 => conv_std_logic_vector(5136, 16),
12396 => conv_std_logic_vector(5184, 16),
12397 => conv_std_logic_vector(5232, 16),
12398 => conv_std_logic_vector(5280, 16),
12399 => conv_std_logic_vector(5328, 16),
12400 => conv_std_logic_vector(5376, 16),
12401 => conv_std_logic_vector(5424, 16),
12402 => conv_std_logic_vector(5472, 16),
12403 => conv_std_logic_vector(5520, 16),
12404 => conv_std_logic_vector(5568, 16),
12405 => conv_std_logic_vector(5616, 16),
12406 => conv_std_logic_vector(5664, 16),
12407 => conv_std_logic_vector(5712, 16),
12408 => conv_std_logic_vector(5760, 16),
12409 => conv_std_logic_vector(5808, 16),
12410 => conv_std_logic_vector(5856, 16),
12411 => conv_std_logic_vector(5904, 16),
12412 => conv_std_logic_vector(5952, 16),
12413 => conv_std_logic_vector(6000, 16),
12414 => conv_std_logic_vector(6048, 16),
12415 => conv_std_logic_vector(6096, 16),
12416 => conv_std_logic_vector(6144, 16),
12417 => conv_std_logic_vector(6192, 16),
12418 => conv_std_logic_vector(6240, 16),
12419 => conv_std_logic_vector(6288, 16),
12420 => conv_std_logic_vector(6336, 16),
12421 => conv_std_logic_vector(6384, 16),
12422 => conv_std_logic_vector(6432, 16),
12423 => conv_std_logic_vector(6480, 16),
12424 => conv_std_logic_vector(6528, 16),
12425 => conv_std_logic_vector(6576, 16),
12426 => conv_std_logic_vector(6624, 16),
12427 => conv_std_logic_vector(6672, 16),
12428 => conv_std_logic_vector(6720, 16),
12429 => conv_std_logic_vector(6768, 16),
12430 => conv_std_logic_vector(6816, 16),
12431 => conv_std_logic_vector(6864, 16),
12432 => conv_std_logic_vector(6912, 16),
12433 => conv_std_logic_vector(6960, 16),
12434 => conv_std_logic_vector(7008, 16),
12435 => conv_std_logic_vector(7056, 16),
12436 => conv_std_logic_vector(7104, 16),
12437 => conv_std_logic_vector(7152, 16),
12438 => conv_std_logic_vector(7200, 16),
12439 => conv_std_logic_vector(7248, 16),
12440 => conv_std_logic_vector(7296, 16),
12441 => conv_std_logic_vector(7344, 16),
12442 => conv_std_logic_vector(7392, 16),
12443 => conv_std_logic_vector(7440, 16),
12444 => conv_std_logic_vector(7488, 16),
12445 => conv_std_logic_vector(7536, 16),
12446 => conv_std_logic_vector(7584, 16),
12447 => conv_std_logic_vector(7632, 16),
12448 => conv_std_logic_vector(7680, 16),
12449 => conv_std_logic_vector(7728, 16),
12450 => conv_std_logic_vector(7776, 16),
12451 => conv_std_logic_vector(7824, 16),
12452 => conv_std_logic_vector(7872, 16),
12453 => conv_std_logic_vector(7920, 16),
12454 => conv_std_logic_vector(7968, 16),
12455 => conv_std_logic_vector(8016, 16),
12456 => conv_std_logic_vector(8064, 16),
12457 => conv_std_logic_vector(8112, 16),
12458 => conv_std_logic_vector(8160, 16),
12459 => conv_std_logic_vector(8208, 16),
12460 => conv_std_logic_vector(8256, 16),
12461 => conv_std_logic_vector(8304, 16),
12462 => conv_std_logic_vector(8352, 16),
12463 => conv_std_logic_vector(8400, 16),
12464 => conv_std_logic_vector(8448, 16),
12465 => conv_std_logic_vector(8496, 16),
12466 => conv_std_logic_vector(8544, 16),
12467 => conv_std_logic_vector(8592, 16),
12468 => conv_std_logic_vector(8640, 16),
12469 => conv_std_logic_vector(8688, 16),
12470 => conv_std_logic_vector(8736, 16),
12471 => conv_std_logic_vector(8784, 16),
12472 => conv_std_logic_vector(8832, 16),
12473 => conv_std_logic_vector(8880, 16),
12474 => conv_std_logic_vector(8928, 16),
12475 => conv_std_logic_vector(8976, 16),
12476 => conv_std_logic_vector(9024, 16),
12477 => conv_std_logic_vector(9072, 16),
12478 => conv_std_logic_vector(9120, 16),
12479 => conv_std_logic_vector(9168, 16),
12480 => conv_std_logic_vector(9216, 16),
12481 => conv_std_logic_vector(9264, 16),
12482 => conv_std_logic_vector(9312, 16),
12483 => conv_std_logic_vector(9360, 16),
12484 => conv_std_logic_vector(9408, 16),
12485 => conv_std_logic_vector(9456, 16),
12486 => conv_std_logic_vector(9504, 16),
12487 => conv_std_logic_vector(9552, 16),
12488 => conv_std_logic_vector(9600, 16),
12489 => conv_std_logic_vector(9648, 16),
12490 => conv_std_logic_vector(9696, 16),
12491 => conv_std_logic_vector(9744, 16),
12492 => conv_std_logic_vector(9792, 16),
12493 => conv_std_logic_vector(9840, 16),
12494 => conv_std_logic_vector(9888, 16),
12495 => conv_std_logic_vector(9936, 16),
12496 => conv_std_logic_vector(9984, 16),
12497 => conv_std_logic_vector(10032, 16),
12498 => conv_std_logic_vector(10080, 16),
12499 => conv_std_logic_vector(10128, 16),
12500 => conv_std_logic_vector(10176, 16),
12501 => conv_std_logic_vector(10224, 16),
12502 => conv_std_logic_vector(10272, 16),
12503 => conv_std_logic_vector(10320, 16),
12504 => conv_std_logic_vector(10368, 16),
12505 => conv_std_logic_vector(10416, 16),
12506 => conv_std_logic_vector(10464, 16),
12507 => conv_std_logic_vector(10512, 16),
12508 => conv_std_logic_vector(10560, 16),
12509 => conv_std_logic_vector(10608, 16),
12510 => conv_std_logic_vector(10656, 16),
12511 => conv_std_logic_vector(10704, 16),
12512 => conv_std_logic_vector(10752, 16),
12513 => conv_std_logic_vector(10800, 16),
12514 => conv_std_logic_vector(10848, 16),
12515 => conv_std_logic_vector(10896, 16),
12516 => conv_std_logic_vector(10944, 16),
12517 => conv_std_logic_vector(10992, 16),
12518 => conv_std_logic_vector(11040, 16),
12519 => conv_std_logic_vector(11088, 16),
12520 => conv_std_logic_vector(11136, 16),
12521 => conv_std_logic_vector(11184, 16),
12522 => conv_std_logic_vector(11232, 16),
12523 => conv_std_logic_vector(11280, 16),
12524 => conv_std_logic_vector(11328, 16),
12525 => conv_std_logic_vector(11376, 16),
12526 => conv_std_logic_vector(11424, 16),
12527 => conv_std_logic_vector(11472, 16),
12528 => conv_std_logic_vector(11520, 16),
12529 => conv_std_logic_vector(11568, 16),
12530 => conv_std_logic_vector(11616, 16),
12531 => conv_std_logic_vector(11664, 16),
12532 => conv_std_logic_vector(11712, 16),
12533 => conv_std_logic_vector(11760, 16),
12534 => conv_std_logic_vector(11808, 16),
12535 => conv_std_logic_vector(11856, 16),
12536 => conv_std_logic_vector(11904, 16),
12537 => conv_std_logic_vector(11952, 16),
12538 => conv_std_logic_vector(12000, 16),
12539 => conv_std_logic_vector(12048, 16),
12540 => conv_std_logic_vector(12096, 16),
12541 => conv_std_logic_vector(12144, 16),
12542 => conv_std_logic_vector(12192, 16),
12543 => conv_std_logic_vector(12240, 16),
12544 => conv_std_logic_vector(0, 16),
12545 => conv_std_logic_vector(49, 16),
12546 => conv_std_logic_vector(98, 16),
12547 => conv_std_logic_vector(147, 16),
12548 => conv_std_logic_vector(196, 16),
12549 => conv_std_logic_vector(245, 16),
12550 => conv_std_logic_vector(294, 16),
12551 => conv_std_logic_vector(343, 16),
12552 => conv_std_logic_vector(392, 16),
12553 => conv_std_logic_vector(441, 16),
12554 => conv_std_logic_vector(490, 16),
12555 => conv_std_logic_vector(539, 16),
12556 => conv_std_logic_vector(588, 16),
12557 => conv_std_logic_vector(637, 16),
12558 => conv_std_logic_vector(686, 16),
12559 => conv_std_logic_vector(735, 16),
12560 => conv_std_logic_vector(784, 16),
12561 => conv_std_logic_vector(833, 16),
12562 => conv_std_logic_vector(882, 16),
12563 => conv_std_logic_vector(931, 16),
12564 => conv_std_logic_vector(980, 16),
12565 => conv_std_logic_vector(1029, 16),
12566 => conv_std_logic_vector(1078, 16),
12567 => conv_std_logic_vector(1127, 16),
12568 => conv_std_logic_vector(1176, 16),
12569 => conv_std_logic_vector(1225, 16),
12570 => conv_std_logic_vector(1274, 16),
12571 => conv_std_logic_vector(1323, 16),
12572 => conv_std_logic_vector(1372, 16),
12573 => conv_std_logic_vector(1421, 16),
12574 => conv_std_logic_vector(1470, 16),
12575 => conv_std_logic_vector(1519, 16),
12576 => conv_std_logic_vector(1568, 16),
12577 => conv_std_logic_vector(1617, 16),
12578 => conv_std_logic_vector(1666, 16),
12579 => conv_std_logic_vector(1715, 16),
12580 => conv_std_logic_vector(1764, 16),
12581 => conv_std_logic_vector(1813, 16),
12582 => conv_std_logic_vector(1862, 16),
12583 => conv_std_logic_vector(1911, 16),
12584 => conv_std_logic_vector(1960, 16),
12585 => conv_std_logic_vector(2009, 16),
12586 => conv_std_logic_vector(2058, 16),
12587 => conv_std_logic_vector(2107, 16),
12588 => conv_std_logic_vector(2156, 16),
12589 => conv_std_logic_vector(2205, 16),
12590 => conv_std_logic_vector(2254, 16),
12591 => conv_std_logic_vector(2303, 16),
12592 => conv_std_logic_vector(2352, 16),
12593 => conv_std_logic_vector(2401, 16),
12594 => conv_std_logic_vector(2450, 16),
12595 => conv_std_logic_vector(2499, 16),
12596 => conv_std_logic_vector(2548, 16),
12597 => conv_std_logic_vector(2597, 16),
12598 => conv_std_logic_vector(2646, 16),
12599 => conv_std_logic_vector(2695, 16),
12600 => conv_std_logic_vector(2744, 16),
12601 => conv_std_logic_vector(2793, 16),
12602 => conv_std_logic_vector(2842, 16),
12603 => conv_std_logic_vector(2891, 16),
12604 => conv_std_logic_vector(2940, 16),
12605 => conv_std_logic_vector(2989, 16),
12606 => conv_std_logic_vector(3038, 16),
12607 => conv_std_logic_vector(3087, 16),
12608 => conv_std_logic_vector(3136, 16),
12609 => conv_std_logic_vector(3185, 16),
12610 => conv_std_logic_vector(3234, 16),
12611 => conv_std_logic_vector(3283, 16),
12612 => conv_std_logic_vector(3332, 16),
12613 => conv_std_logic_vector(3381, 16),
12614 => conv_std_logic_vector(3430, 16),
12615 => conv_std_logic_vector(3479, 16),
12616 => conv_std_logic_vector(3528, 16),
12617 => conv_std_logic_vector(3577, 16),
12618 => conv_std_logic_vector(3626, 16),
12619 => conv_std_logic_vector(3675, 16),
12620 => conv_std_logic_vector(3724, 16),
12621 => conv_std_logic_vector(3773, 16),
12622 => conv_std_logic_vector(3822, 16),
12623 => conv_std_logic_vector(3871, 16),
12624 => conv_std_logic_vector(3920, 16),
12625 => conv_std_logic_vector(3969, 16),
12626 => conv_std_logic_vector(4018, 16),
12627 => conv_std_logic_vector(4067, 16),
12628 => conv_std_logic_vector(4116, 16),
12629 => conv_std_logic_vector(4165, 16),
12630 => conv_std_logic_vector(4214, 16),
12631 => conv_std_logic_vector(4263, 16),
12632 => conv_std_logic_vector(4312, 16),
12633 => conv_std_logic_vector(4361, 16),
12634 => conv_std_logic_vector(4410, 16),
12635 => conv_std_logic_vector(4459, 16),
12636 => conv_std_logic_vector(4508, 16),
12637 => conv_std_logic_vector(4557, 16),
12638 => conv_std_logic_vector(4606, 16),
12639 => conv_std_logic_vector(4655, 16),
12640 => conv_std_logic_vector(4704, 16),
12641 => conv_std_logic_vector(4753, 16),
12642 => conv_std_logic_vector(4802, 16),
12643 => conv_std_logic_vector(4851, 16),
12644 => conv_std_logic_vector(4900, 16),
12645 => conv_std_logic_vector(4949, 16),
12646 => conv_std_logic_vector(4998, 16),
12647 => conv_std_logic_vector(5047, 16),
12648 => conv_std_logic_vector(5096, 16),
12649 => conv_std_logic_vector(5145, 16),
12650 => conv_std_logic_vector(5194, 16),
12651 => conv_std_logic_vector(5243, 16),
12652 => conv_std_logic_vector(5292, 16),
12653 => conv_std_logic_vector(5341, 16),
12654 => conv_std_logic_vector(5390, 16),
12655 => conv_std_logic_vector(5439, 16),
12656 => conv_std_logic_vector(5488, 16),
12657 => conv_std_logic_vector(5537, 16),
12658 => conv_std_logic_vector(5586, 16),
12659 => conv_std_logic_vector(5635, 16),
12660 => conv_std_logic_vector(5684, 16),
12661 => conv_std_logic_vector(5733, 16),
12662 => conv_std_logic_vector(5782, 16),
12663 => conv_std_logic_vector(5831, 16),
12664 => conv_std_logic_vector(5880, 16),
12665 => conv_std_logic_vector(5929, 16),
12666 => conv_std_logic_vector(5978, 16),
12667 => conv_std_logic_vector(6027, 16),
12668 => conv_std_logic_vector(6076, 16),
12669 => conv_std_logic_vector(6125, 16),
12670 => conv_std_logic_vector(6174, 16),
12671 => conv_std_logic_vector(6223, 16),
12672 => conv_std_logic_vector(6272, 16),
12673 => conv_std_logic_vector(6321, 16),
12674 => conv_std_logic_vector(6370, 16),
12675 => conv_std_logic_vector(6419, 16),
12676 => conv_std_logic_vector(6468, 16),
12677 => conv_std_logic_vector(6517, 16),
12678 => conv_std_logic_vector(6566, 16),
12679 => conv_std_logic_vector(6615, 16),
12680 => conv_std_logic_vector(6664, 16),
12681 => conv_std_logic_vector(6713, 16),
12682 => conv_std_logic_vector(6762, 16),
12683 => conv_std_logic_vector(6811, 16),
12684 => conv_std_logic_vector(6860, 16),
12685 => conv_std_logic_vector(6909, 16),
12686 => conv_std_logic_vector(6958, 16),
12687 => conv_std_logic_vector(7007, 16),
12688 => conv_std_logic_vector(7056, 16),
12689 => conv_std_logic_vector(7105, 16),
12690 => conv_std_logic_vector(7154, 16),
12691 => conv_std_logic_vector(7203, 16),
12692 => conv_std_logic_vector(7252, 16),
12693 => conv_std_logic_vector(7301, 16),
12694 => conv_std_logic_vector(7350, 16),
12695 => conv_std_logic_vector(7399, 16),
12696 => conv_std_logic_vector(7448, 16),
12697 => conv_std_logic_vector(7497, 16),
12698 => conv_std_logic_vector(7546, 16),
12699 => conv_std_logic_vector(7595, 16),
12700 => conv_std_logic_vector(7644, 16),
12701 => conv_std_logic_vector(7693, 16),
12702 => conv_std_logic_vector(7742, 16),
12703 => conv_std_logic_vector(7791, 16),
12704 => conv_std_logic_vector(7840, 16),
12705 => conv_std_logic_vector(7889, 16),
12706 => conv_std_logic_vector(7938, 16),
12707 => conv_std_logic_vector(7987, 16),
12708 => conv_std_logic_vector(8036, 16),
12709 => conv_std_logic_vector(8085, 16),
12710 => conv_std_logic_vector(8134, 16),
12711 => conv_std_logic_vector(8183, 16),
12712 => conv_std_logic_vector(8232, 16),
12713 => conv_std_logic_vector(8281, 16),
12714 => conv_std_logic_vector(8330, 16),
12715 => conv_std_logic_vector(8379, 16),
12716 => conv_std_logic_vector(8428, 16),
12717 => conv_std_logic_vector(8477, 16),
12718 => conv_std_logic_vector(8526, 16),
12719 => conv_std_logic_vector(8575, 16),
12720 => conv_std_logic_vector(8624, 16),
12721 => conv_std_logic_vector(8673, 16),
12722 => conv_std_logic_vector(8722, 16),
12723 => conv_std_logic_vector(8771, 16),
12724 => conv_std_logic_vector(8820, 16),
12725 => conv_std_logic_vector(8869, 16),
12726 => conv_std_logic_vector(8918, 16),
12727 => conv_std_logic_vector(8967, 16),
12728 => conv_std_logic_vector(9016, 16),
12729 => conv_std_logic_vector(9065, 16),
12730 => conv_std_logic_vector(9114, 16),
12731 => conv_std_logic_vector(9163, 16),
12732 => conv_std_logic_vector(9212, 16),
12733 => conv_std_logic_vector(9261, 16),
12734 => conv_std_logic_vector(9310, 16),
12735 => conv_std_logic_vector(9359, 16),
12736 => conv_std_logic_vector(9408, 16),
12737 => conv_std_logic_vector(9457, 16),
12738 => conv_std_logic_vector(9506, 16),
12739 => conv_std_logic_vector(9555, 16),
12740 => conv_std_logic_vector(9604, 16),
12741 => conv_std_logic_vector(9653, 16),
12742 => conv_std_logic_vector(9702, 16),
12743 => conv_std_logic_vector(9751, 16),
12744 => conv_std_logic_vector(9800, 16),
12745 => conv_std_logic_vector(9849, 16),
12746 => conv_std_logic_vector(9898, 16),
12747 => conv_std_logic_vector(9947, 16),
12748 => conv_std_logic_vector(9996, 16),
12749 => conv_std_logic_vector(10045, 16),
12750 => conv_std_logic_vector(10094, 16),
12751 => conv_std_logic_vector(10143, 16),
12752 => conv_std_logic_vector(10192, 16),
12753 => conv_std_logic_vector(10241, 16),
12754 => conv_std_logic_vector(10290, 16),
12755 => conv_std_logic_vector(10339, 16),
12756 => conv_std_logic_vector(10388, 16),
12757 => conv_std_logic_vector(10437, 16),
12758 => conv_std_logic_vector(10486, 16),
12759 => conv_std_logic_vector(10535, 16),
12760 => conv_std_logic_vector(10584, 16),
12761 => conv_std_logic_vector(10633, 16),
12762 => conv_std_logic_vector(10682, 16),
12763 => conv_std_logic_vector(10731, 16),
12764 => conv_std_logic_vector(10780, 16),
12765 => conv_std_logic_vector(10829, 16),
12766 => conv_std_logic_vector(10878, 16),
12767 => conv_std_logic_vector(10927, 16),
12768 => conv_std_logic_vector(10976, 16),
12769 => conv_std_logic_vector(11025, 16),
12770 => conv_std_logic_vector(11074, 16),
12771 => conv_std_logic_vector(11123, 16),
12772 => conv_std_logic_vector(11172, 16),
12773 => conv_std_logic_vector(11221, 16),
12774 => conv_std_logic_vector(11270, 16),
12775 => conv_std_logic_vector(11319, 16),
12776 => conv_std_logic_vector(11368, 16),
12777 => conv_std_logic_vector(11417, 16),
12778 => conv_std_logic_vector(11466, 16),
12779 => conv_std_logic_vector(11515, 16),
12780 => conv_std_logic_vector(11564, 16),
12781 => conv_std_logic_vector(11613, 16),
12782 => conv_std_logic_vector(11662, 16),
12783 => conv_std_logic_vector(11711, 16),
12784 => conv_std_logic_vector(11760, 16),
12785 => conv_std_logic_vector(11809, 16),
12786 => conv_std_logic_vector(11858, 16),
12787 => conv_std_logic_vector(11907, 16),
12788 => conv_std_logic_vector(11956, 16),
12789 => conv_std_logic_vector(12005, 16),
12790 => conv_std_logic_vector(12054, 16),
12791 => conv_std_logic_vector(12103, 16),
12792 => conv_std_logic_vector(12152, 16),
12793 => conv_std_logic_vector(12201, 16),
12794 => conv_std_logic_vector(12250, 16),
12795 => conv_std_logic_vector(12299, 16),
12796 => conv_std_logic_vector(12348, 16),
12797 => conv_std_logic_vector(12397, 16),
12798 => conv_std_logic_vector(12446, 16),
12799 => conv_std_logic_vector(12495, 16),
12800 => conv_std_logic_vector(0, 16),
12801 => conv_std_logic_vector(50, 16),
12802 => conv_std_logic_vector(100, 16),
12803 => conv_std_logic_vector(150, 16),
12804 => conv_std_logic_vector(200, 16),
12805 => conv_std_logic_vector(250, 16),
12806 => conv_std_logic_vector(300, 16),
12807 => conv_std_logic_vector(350, 16),
12808 => conv_std_logic_vector(400, 16),
12809 => conv_std_logic_vector(450, 16),
12810 => conv_std_logic_vector(500, 16),
12811 => conv_std_logic_vector(550, 16),
12812 => conv_std_logic_vector(600, 16),
12813 => conv_std_logic_vector(650, 16),
12814 => conv_std_logic_vector(700, 16),
12815 => conv_std_logic_vector(750, 16),
12816 => conv_std_logic_vector(800, 16),
12817 => conv_std_logic_vector(850, 16),
12818 => conv_std_logic_vector(900, 16),
12819 => conv_std_logic_vector(950, 16),
12820 => conv_std_logic_vector(1000, 16),
12821 => conv_std_logic_vector(1050, 16),
12822 => conv_std_logic_vector(1100, 16),
12823 => conv_std_logic_vector(1150, 16),
12824 => conv_std_logic_vector(1200, 16),
12825 => conv_std_logic_vector(1250, 16),
12826 => conv_std_logic_vector(1300, 16),
12827 => conv_std_logic_vector(1350, 16),
12828 => conv_std_logic_vector(1400, 16),
12829 => conv_std_logic_vector(1450, 16),
12830 => conv_std_logic_vector(1500, 16),
12831 => conv_std_logic_vector(1550, 16),
12832 => conv_std_logic_vector(1600, 16),
12833 => conv_std_logic_vector(1650, 16),
12834 => conv_std_logic_vector(1700, 16),
12835 => conv_std_logic_vector(1750, 16),
12836 => conv_std_logic_vector(1800, 16),
12837 => conv_std_logic_vector(1850, 16),
12838 => conv_std_logic_vector(1900, 16),
12839 => conv_std_logic_vector(1950, 16),
12840 => conv_std_logic_vector(2000, 16),
12841 => conv_std_logic_vector(2050, 16),
12842 => conv_std_logic_vector(2100, 16),
12843 => conv_std_logic_vector(2150, 16),
12844 => conv_std_logic_vector(2200, 16),
12845 => conv_std_logic_vector(2250, 16),
12846 => conv_std_logic_vector(2300, 16),
12847 => conv_std_logic_vector(2350, 16),
12848 => conv_std_logic_vector(2400, 16),
12849 => conv_std_logic_vector(2450, 16),
12850 => conv_std_logic_vector(2500, 16),
12851 => conv_std_logic_vector(2550, 16),
12852 => conv_std_logic_vector(2600, 16),
12853 => conv_std_logic_vector(2650, 16),
12854 => conv_std_logic_vector(2700, 16),
12855 => conv_std_logic_vector(2750, 16),
12856 => conv_std_logic_vector(2800, 16),
12857 => conv_std_logic_vector(2850, 16),
12858 => conv_std_logic_vector(2900, 16),
12859 => conv_std_logic_vector(2950, 16),
12860 => conv_std_logic_vector(3000, 16),
12861 => conv_std_logic_vector(3050, 16),
12862 => conv_std_logic_vector(3100, 16),
12863 => conv_std_logic_vector(3150, 16),
12864 => conv_std_logic_vector(3200, 16),
12865 => conv_std_logic_vector(3250, 16),
12866 => conv_std_logic_vector(3300, 16),
12867 => conv_std_logic_vector(3350, 16),
12868 => conv_std_logic_vector(3400, 16),
12869 => conv_std_logic_vector(3450, 16),
12870 => conv_std_logic_vector(3500, 16),
12871 => conv_std_logic_vector(3550, 16),
12872 => conv_std_logic_vector(3600, 16),
12873 => conv_std_logic_vector(3650, 16),
12874 => conv_std_logic_vector(3700, 16),
12875 => conv_std_logic_vector(3750, 16),
12876 => conv_std_logic_vector(3800, 16),
12877 => conv_std_logic_vector(3850, 16),
12878 => conv_std_logic_vector(3900, 16),
12879 => conv_std_logic_vector(3950, 16),
12880 => conv_std_logic_vector(4000, 16),
12881 => conv_std_logic_vector(4050, 16),
12882 => conv_std_logic_vector(4100, 16),
12883 => conv_std_logic_vector(4150, 16),
12884 => conv_std_logic_vector(4200, 16),
12885 => conv_std_logic_vector(4250, 16),
12886 => conv_std_logic_vector(4300, 16),
12887 => conv_std_logic_vector(4350, 16),
12888 => conv_std_logic_vector(4400, 16),
12889 => conv_std_logic_vector(4450, 16),
12890 => conv_std_logic_vector(4500, 16),
12891 => conv_std_logic_vector(4550, 16),
12892 => conv_std_logic_vector(4600, 16),
12893 => conv_std_logic_vector(4650, 16),
12894 => conv_std_logic_vector(4700, 16),
12895 => conv_std_logic_vector(4750, 16),
12896 => conv_std_logic_vector(4800, 16),
12897 => conv_std_logic_vector(4850, 16),
12898 => conv_std_logic_vector(4900, 16),
12899 => conv_std_logic_vector(4950, 16),
12900 => conv_std_logic_vector(5000, 16),
12901 => conv_std_logic_vector(5050, 16),
12902 => conv_std_logic_vector(5100, 16),
12903 => conv_std_logic_vector(5150, 16),
12904 => conv_std_logic_vector(5200, 16),
12905 => conv_std_logic_vector(5250, 16),
12906 => conv_std_logic_vector(5300, 16),
12907 => conv_std_logic_vector(5350, 16),
12908 => conv_std_logic_vector(5400, 16),
12909 => conv_std_logic_vector(5450, 16),
12910 => conv_std_logic_vector(5500, 16),
12911 => conv_std_logic_vector(5550, 16),
12912 => conv_std_logic_vector(5600, 16),
12913 => conv_std_logic_vector(5650, 16),
12914 => conv_std_logic_vector(5700, 16),
12915 => conv_std_logic_vector(5750, 16),
12916 => conv_std_logic_vector(5800, 16),
12917 => conv_std_logic_vector(5850, 16),
12918 => conv_std_logic_vector(5900, 16),
12919 => conv_std_logic_vector(5950, 16),
12920 => conv_std_logic_vector(6000, 16),
12921 => conv_std_logic_vector(6050, 16),
12922 => conv_std_logic_vector(6100, 16),
12923 => conv_std_logic_vector(6150, 16),
12924 => conv_std_logic_vector(6200, 16),
12925 => conv_std_logic_vector(6250, 16),
12926 => conv_std_logic_vector(6300, 16),
12927 => conv_std_logic_vector(6350, 16),
12928 => conv_std_logic_vector(6400, 16),
12929 => conv_std_logic_vector(6450, 16),
12930 => conv_std_logic_vector(6500, 16),
12931 => conv_std_logic_vector(6550, 16),
12932 => conv_std_logic_vector(6600, 16),
12933 => conv_std_logic_vector(6650, 16),
12934 => conv_std_logic_vector(6700, 16),
12935 => conv_std_logic_vector(6750, 16),
12936 => conv_std_logic_vector(6800, 16),
12937 => conv_std_logic_vector(6850, 16),
12938 => conv_std_logic_vector(6900, 16),
12939 => conv_std_logic_vector(6950, 16),
12940 => conv_std_logic_vector(7000, 16),
12941 => conv_std_logic_vector(7050, 16),
12942 => conv_std_logic_vector(7100, 16),
12943 => conv_std_logic_vector(7150, 16),
12944 => conv_std_logic_vector(7200, 16),
12945 => conv_std_logic_vector(7250, 16),
12946 => conv_std_logic_vector(7300, 16),
12947 => conv_std_logic_vector(7350, 16),
12948 => conv_std_logic_vector(7400, 16),
12949 => conv_std_logic_vector(7450, 16),
12950 => conv_std_logic_vector(7500, 16),
12951 => conv_std_logic_vector(7550, 16),
12952 => conv_std_logic_vector(7600, 16),
12953 => conv_std_logic_vector(7650, 16),
12954 => conv_std_logic_vector(7700, 16),
12955 => conv_std_logic_vector(7750, 16),
12956 => conv_std_logic_vector(7800, 16),
12957 => conv_std_logic_vector(7850, 16),
12958 => conv_std_logic_vector(7900, 16),
12959 => conv_std_logic_vector(7950, 16),
12960 => conv_std_logic_vector(8000, 16),
12961 => conv_std_logic_vector(8050, 16),
12962 => conv_std_logic_vector(8100, 16),
12963 => conv_std_logic_vector(8150, 16),
12964 => conv_std_logic_vector(8200, 16),
12965 => conv_std_logic_vector(8250, 16),
12966 => conv_std_logic_vector(8300, 16),
12967 => conv_std_logic_vector(8350, 16),
12968 => conv_std_logic_vector(8400, 16),
12969 => conv_std_logic_vector(8450, 16),
12970 => conv_std_logic_vector(8500, 16),
12971 => conv_std_logic_vector(8550, 16),
12972 => conv_std_logic_vector(8600, 16),
12973 => conv_std_logic_vector(8650, 16),
12974 => conv_std_logic_vector(8700, 16),
12975 => conv_std_logic_vector(8750, 16),
12976 => conv_std_logic_vector(8800, 16),
12977 => conv_std_logic_vector(8850, 16),
12978 => conv_std_logic_vector(8900, 16),
12979 => conv_std_logic_vector(8950, 16),
12980 => conv_std_logic_vector(9000, 16),
12981 => conv_std_logic_vector(9050, 16),
12982 => conv_std_logic_vector(9100, 16),
12983 => conv_std_logic_vector(9150, 16),
12984 => conv_std_logic_vector(9200, 16),
12985 => conv_std_logic_vector(9250, 16),
12986 => conv_std_logic_vector(9300, 16),
12987 => conv_std_logic_vector(9350, 16),
12988 => conv_std_logic_vector(9400, 16),
12989 => conv_std_logic_vector(9450, 16),
12990 => conv_std_logic_vector(9500, 16),
12991 => conv_std_logic_vector(9550, 16),
12992 => conv_std_logic_vector(9600, 16),
12993 => conv_std_logic_vector(9650, 16),
12994 => conv_std_logic_vector(9700, 16),
12995 => conv_std_logic_vector(9750, 16),
12996 => conv_std_logic_vector(9800, 16),
12997 => conv_std_logic_vector(9850, 16),
12998 => conv_std_logic_vector(9900, 16),
12999 => conv_std_logic_vector(9950, 16),
13000 => conv_std_logic_vector(10000, 16),
13001 => conv_std_logic_vector(10050, 16),
13002 => conv_std_logic_vector(10100, 16),
13003 => conv_std_logic_vector(10150, 16),
13004 => conv_std_logic_vector(10200, 16),
13005 => conv_std_logic_vector(10250, 16),
13006 => conv_std_logic_vector(10300, 16),
13007 => conv_std_logic_vector(10350, 16),
13008 => conv_std_logic_vector(10400, 16),
13009 => conv_std_logic_vector(10450, 16),
13010 => conv_std_logic_vector(10500, 16),
13011 => conv_std_logic_vector(10550, 16),
13012 => conv_std_logic_vector(10600, 16),
13013 => conv_std_logic_vector(10650, 16),
13014 => conv_std_logic_vector(10700, 16),
13015 => conv_std_logic_vector(10750, 16),
13016 => conv_std_logic_vector(10800, 16),
13017 => conv_std_logic_vector(10850, 16),
13018 => conv_std_logic_vector(10900, 16),
13019 => conv_std_logic_vector(10950, 16),
13020 => conv_std_logic_vector(11000, 16),
13021 => conv_std_logic_vector(11050, 16),
13022 => conv_std_logic_vector(11100, 16),
13023 => conv_std_logic_vector(11150, 16),
13024 => conv_std_logic_vector(11200, 16),
13025 => conv_std_logic_vector(11250, 16),
13026 => conv_std_logic_vector(11300, 16),
13027 => conv_std_logic_vector(11350, 16),
13028 => conv_std_logic_vector(11400, 16),
13029 => conv_std_logic_vector(11450, 16),
13030 => conv_std_logic_vector(11500, 16),
13031 => conv_std_logic_vector(11550, 16),
13032 => conv_std_logic_vector(11600, 16),
13033 => conv_std_logic_vector(11650, 16),
13034 => conv_std_logic_vector(11700, 16),
13035 => conv_std_logic_vector(11750, 16),
13036 => conv_std_logic_vector(11800, 16),
13037 => conv_std_logic_vector(11850, 16),
13038 => conv_std_logic_vector(11900, 16),
13039 => conv_std_logic_vector(11950, 16),
13040 => conv_std_logic_vector(12000, 16),
13041 => conv_std_logic_vector(12050, 16),
13042 => conv_std_logic_vector(12100, 16),
13043 => conv_std_logic_vector(12150, 16),
13044 => conv_std_logic_vector(12200, 16),
13045 => conv_std_logic_vector(12250, 16),
13046 => conv_std_logic_vector(12300, 16),
13047 => conv_std_logic_vector(12350, 16),
13048 => conv_std_logic_vector(12400, 16),
13049 => conv_std_logic_vector(12450, 16),
13050 => conv_std_logic_vector(12500, 16),
13051 => conv_std_logic_vector(12550, 16),
13052 => conv_std_logic_vector(12600, 16),
13053 => conv_std_logic_vector(12650, 16),
13054 => conv_std_logic_vector(12700, 16),
13055 => conv_std_logic_vector(12750, 16),
13056 => conv_std_logic_vector(0, 16),
13057 => conv_std_logic_vector(51, 16),
13058 => conv_std_logic_vector(102, 16),
13059 => conv_std_logic_vector(153, 16),
13060 => conv_std_logic_vector(204, 16),
13061 => conv_std_logic_vector(255, 16),
13062 => conv_std_logic_vector(306, 16),
13063 => conv_std_logic_vector(357, 16),
13064 => conv_std_logic_vector(408, 16),
13065 => conv_std_logic_vector(459, 16),
13066 => conv_std_logic_vector(510, 16),
13067 => conv_std_logic_vector(561, 16),
13068 => conv_std_logic_vector(612, 16),
13069 => conv_std_logic_vector(663, 16),
13070 => conv_std_logic_vector(714, 16),
13071 => conv_std_logic_vector(765, 16),
13072 => conv_std_logic_vector(816, 16),
13073 => conv_std_logic_vector(867, 16),
13074 => conv_std_logic_vector(918, 16),
13075 => conv_std_logic_vector(969, 16),
13076 => conv_std_logic_vector(1020, 16),
13077 => conv_std_logic_vector(1071, 16),
13078 => conv_std_logic_vector(1122, 16),
13079 => conv_std_logic_vector(1173, 16),
13080 => conv_std_logic_vector(1224, 16),
13081 => conv_std_logic_vector(1275, 16),
13082 => conv_std_logic_vector(1326, 16),
13083 => conv_std_logic_vector(1377, 16),
13084 => conv_std_logic_vector(1428, 16),
13085 => conv_std_logic_vector(1479, 16),
13086 => conv_std_logic_vector(1530, 16),
13087 => conv_std_logic_vector(1581, 16),
13088 => conv_std_logic_vector(1632, 16),
13089 => conv_std_logic_vector(1683, 16),
13090 => conv_std_logic_vector(1734, 16),
13091 => conv_std_logic_vector(1785, 16),
13092 => conv_std_logic_vector(1836, 16),
13093 => conv_std_logic_vector(1887, 16),
13094 => conv_std_logic_vector(1938, 16),
13095 => conv_std_logic_vector(1989, 16),
13096 => conv_std_logic_vector(2040, 16),
13097 => conv_std_logic_vector(2091, 16),
13098 => conv_std_logic_vector(2142, 16),
13099 => conv_std_logic_vector(2193, 16),
13100 => conv_std_logic_vector(2244, 16),
13101 => conv_std_logic_vector(2295, 16),
13102 => conv_std_logic_vector(2346, 16),
13103 => conv_std_logic_vector(2397, 16),
13104 => conv_std_logic_vector(2448, 16),
13105 => conv_std_logic_vector(2499, 16),
13106 => conv_std_logic_vector(2550, 16),
13107 => conv_std_logic_vector(2601, 16),
13108 => conv_std_logic_vector(2652, 16),
13109 => conv_std_logic_vector(2703, 16),
13110 => conv_std_logic_vector(2754, 16),
13111 => conv_std_logic_vector(2805, 16),
13112 => conv_std_logic_vector(2856, 16),
13113 => conv_std_logic_vector(2907, 16),
13114 => conv_std_logic_vector(2958, 16),
13115 => conv_std_logic_vector(3009, 16),
13116 => conv_std_logic_vector(3060, 16),
13117 => conv_std_logic_vector(3111, 16),
13118 => conv_std_logic_vector(3162, 16),
13119 => conv_std_logic_vector(3213, 16),
13120 => conv_std_logic_vector(3264, 16),
13121 => conv_std_logic_vector(3315, 16),
13122 => conv_std_logic_vector(3366, 16),
13123 => conv_std_logic_vector(3417, 16),
13124 => conv_std_logic_vector(3468, 16),
13125 => conv_std_logic_vector(3519, 16),
13126 => conv_std_logic_vector(3570, 16),
13127 => conv_std_logic_vector(3621, 16),
13128 => conv_std_logic_vector(3672, 16),
13129 => conv_std_logic_vector(3723, 16),
13130 => conv_std_logic_vector(3774, 16),
13131 => conv_std_logic_vector(3825, 16),
13132 => conv_std_logic_vector(3876, 16),
13133 => conv_std_logic_vector(3927, 16),
13134 => conv_std_logic_vector(3978, 16),
13135 => conv_std_logic_vector(4029, 16),
13136 => conv_std_logic_vector(4080, 16),
13137 => conv_std_logic_vector(4131, 16),
13138 => conv_std_logic_vector(4182, 16),
13139 => conv_std_logic_vector(4233, 16),
13140 => conv_std_logic_vector(4284, 16),
13141 => conv_std_logic_vector(4335, 16),
13142 => conv_std_logic_vector(4386, 16),
13143 => conv_std_logic_vector(4437, 16),
13144 => conv_std_logic_vector(4488, 16),
13145 => conv_std_logic_vector(4539, 16),
13146 => conv_std_logic_vector(4590, 16),
13147 => conv_std_logic_vector(4641, 16),
13148 => conv_std_logic_vector(4692, 16),
13149 => conv_std_logic_vector(4743, 16),
13150 => conv_std_logic_vector(4794, 16),
13151 => conv_std_logic_vector(4845, 16),
13152 => conv_std_logic_vector(4896, 16),
13153 => conv_std_logic_vector(4947, 16),
13154 => conv_std_logic_vector(4998, 16),
13155 => conv_std_logic_vector(5049, 16),
13156 => conv_std_logic_vector(5100, 16),
13157 => conv_std_logic_vector(5151, 16),
13158 => conv_std_logic_vector(5202, 16),
13159 => conv_std_logic_vector(5253, 16),
13160 => conv_std_logic_vector(5304, 16),
13161 => conv_std_logic_vector(5355, 16),
13162 => conv_std_logic_vector(5406, 16),
13163 => conv_std_logic_vector(5457, 16),
13164 => conv_std_logic_vector(5508, 16),
13165 => conv_std_logic_vector(5559, 16),
13166 => conv_std_logic_vector(5610, 16),
13167 => conv_std_logic_vector(5661, 16),
13168 => conv_std_logic_vector(5712, 16),
13169 => conv_std_logic_vector(5763, 16),
13170 => conv_std_logic_vector(5814, 16),
13171 => conv_std_logic_vector(5865, 16),
13172 => conv_std_logic_vector(5916, 16),
13173 => conv_std_logic_vector(5967, 16),
13174 => conv_std_logic_vector(6018, 16),
13175 => conv_std_logic_vector(6069, 16),
13176 => conv_std_logic_vector(6120, 16),
13177 => conv_std_logic_vector(6171, 16),
13178 => conv_std_logic_vector(6222, 16),
13179 => conv_std_logic_vector(6273, 16),
13180 => conv_std_logic_vector(6324, 16),
13181 => conv_std_logic_vector(6375, 16),
13182 => conv_std_logic_vector(6426, 16),
13183 => conv_std_logic_vector(6477, 16),
13184 => conv_std_logic_vector(6528, 16),
13185 => conv_std_logic_vector(6579, 16),
13186 => conv_std_logic_vector(6630, 16),
13187 => conv_std_logic_vector(6681, 16),
13188 => conv_std_logic_vector(6732, 16),
13189 => conv_std_logic_vector(6783, 16),
13190 => conv_std_logic_vector(6834, 16),
13191 => conv_std_logic_vector(6885, 16),
13192 => conv_std_logic_vector(6936, 16),
13193 => conv_std_logic_vector(6987, 16),
13194 => conv_std_logic_vector(7038, 16),
13195 => conv_std_logic_vector(7089, 16),
13196 => conv_std_logic_vector(7140, 16),
13197 => conv_std_logic_vector(7191, 16),
13198 => conv_std_logic_vector(7242, 16),
13199 => conv_std_logic_vector(7293, 16),
13200 => conv_std_logic_vector(7344, 16),
13201 => conv_std_logic_vector(7395, 16),
13202 => conv_std_logic_vector(7446, 16),
13203 => conv_std_logic_vector(7497, 16),
13204 => conv_std_logic_vector(7548, 16),
13205 => conv_std_logic_vector(7599, 16),
13206 => conv_std_logic_vector(7650, 16),
13207 => conv_std_logic_vector(7701, 16),
13208 => conv_std_logic_vector(7752, 16),
13209 => conv_std_logic_vector(7803, 16),
13210 => conv_std_logic_vector(7854, 16),
13211 => conv_std_logic_vector(7905, 16),
13212 => conv_std_logic_vector(7956, 16),
13213 => conv_std_logic_vector(8007, 16),
13214 => conv_std_logic_vector(8058, 16),
13215 => conv_std_logic_vector(8109, 16),
13216 => conv_std_logic_vector(8160, 16),
13217 => conv_std_logic_vector(8211, 16),
13218 => conv_std_logic_vector(8262, 16),
13219 => conv_std_logic_vector(8313, 16),
13220 => conv_std_logic_vector(8364, 16),
13221 => conv_std_logic_vector(8415, 16),
13222 => conv_std_logic_vector(8466, 16),
13223 => conv_std_logic_vector(8517, 16),
13224 => conv_std_logic_vector(8568, 16),
13225 => conv_std_logic_vector(8619, 16),
13226 => conv_std_logic_vector(8670, 16),
13227 => conv_std_logic_vector(8721, 16),
13228 => conv_std_logic_vector(8772, 16),
13229 => conv_std_logic_vector(8823, 16),
13230 => conv_std_logic_vector(8874, 16),
13231 => conv_std_logic_vector(8925, 16),
13232 => conv_std_logic_vector(8976, 16),
13233 => conv_std_logic_vector(9027, 16),
13234 => conv_std_logic_vector(9078, 16),
13235 => conv_std_logic_vector(9129, 16),
13236 => conv_std_logic_vector(9180, 16),
13237 => conv_std_logic_vector(9231, 16),
13238 => conv_std_logic_vector(9282, 16),
13239 => conv_std_logic_vector(9333, 16),
13240 => conv_std_logic_vector(9384, 16),
13241 => conv_std_logic_vector(9435, 16),
13242 => conv_std_logic_vector(9486, 16),
13243 => conv_std_logic_vector(9537, 16),
13244 => conv_std_logic_vector(9588, 16),
13245 => conv_std_logic_vector(9639, 16),
13246 => conv_std_logic_vector(9690, 16),
13247 => conv_std_logic_vector(9741, 16),
13248 => conv_std_logic_vector(9792, 16),
13249 => conv_std_logic_vector(9843, 16),
13250 => conv_std_logic_vector(9894, 16),
13251 => conv_std_logic_vector(9945, 16),
13252 => conv_std_logic_vector(9996, 16),
13253 => conv_std_logic_vector(10047, 16),
13254 => conv_std_logic_vector(10098, 16),
13255 => conv_std_logic_vector(10149, 16),
13256 => conv_std_logic_vector(10200, 16),
13257 => conv_std_logic_vector(10251, 16),
13258 => conv_std_logic_vector(10302, 16),
13259 => conv_std_logic_vector(10353, 16),
13260 => conv_std_logic_vector(10404, 16),
13261 => conv_std_logic_vector(10455, 16),
13262 => conv_std_logic_vector(10506, 16),
13263 => conv_std_logic_vector(10557, 16),
13264 => conv_std_logic_vector(10608, 16),
13265 => conv_std_logic_vector(10659, 16),
13266 => conv_std_logic_vector(10710, 16),
13267 => conv_std_logic_vector(10761, 16),
13268 => conv_std_logic_vector(10812, 16),
13269 => conv_std_logic_vector(10863, 16),
13270 => conv_std_logic_vector(10914, 16),
13271 => conv_std_logic_vector(10965, 16),
13272 => conv_std_logic_vector(11016, 16),
13273 => conv_std_logic_vector(11067, 16),
13274 => conv_std_logic_vector(11118, 16),
13275 => conv_std_logic_vector(11169, 16),
13276 => conv_std_logic_vector(11220, 16),
13277 => conv_std_logic_vector(11271, 16),
13278 => conv_std_logic_vector(11322, 16),
13279 => conv_std_logic_vector(11373, 16),
13280 => conv_std_logic_vector(11424, 16),
13281 => conv_std_logic_vector(11475, 16),
13282 => conv_std_logic_vector(11526, 16),
13283 => conv_std_logic_vector(11577, 16),
13284 => conv_std_logic_vector(11628, 16),
13285 => conv_std_logic_vector(11679, 16),
13286 => conv_std_logic_vector(11730, 16),
13287 => conv_std_logic_vector(11781, 16),
13288 => conv_std_logic_vector(11832, 16),
13289 => conv_std_logic_vector(11883, 16),
13290 => conv_std_logic_vector(11934, 16),
13291 => conv_std_logic_vector(11985, 16),
13292 => conv_std_logic_vector(12036, 16),
13293 => conv_std_logic_vector(12087, 16),
13294 => conv_std_logic_vector(12138, 16),
13295 => conv_std_logic_vector(12189, 16),
13296 => conv_std_logic_vector(12240, 16),
13297 => conv_std_logic_vector(12291, 16),
13298 => conv_std_logic_vector(12342, 16),
13299 => conv_std_logic_vector(12393, 16),
13300 => conv_std_logic_vector(12444, 16),
13301 => conv_std_logic_vector(12495, 16),
13302 => conv_std_logic_vector(12546, 16),
13303 => conv_std_logic_vector(12597, 16),
13304 => conv_std_logic_vector(12648, 16),
13305 => conv_std_logic_vector(12699, 16),
13306 => conv_std_logic_vector(12750, 16),
13307 => conv_std_logic_vector(12801, 16),
13308 => conv_std_logic_vector(12852, 16),
13309 => conv_std_logic_vector(12903, 16),
13310 => conv_std_logic_vector(12954, 16),
13311 => conv_std_logic_vector(13005, 16),
13312 => conv_std_logic_vector(0, 16),
13313 => conv_std_logic_vector(52, 16),
13314 => conv_std_logic_vector(104, 16),
13315 => conv_std_logic_vector(156, 16),
13316 => conv_std_logic_vector(208, 16),
13317 => conv_std_logic_vector(260, 16),
13318 => conv_std_logic_vector(312, 16),
13319 => conv_std_logic_vector(364, 16),
13320 => conv_std_logic_vector(416, 16),
13321 => conv_std_logic_vector(468, 16),
13322 => conv_std_logic_vector(520, 16),
13323 => conv_std_logic_vector(572, 16),
13324 => conv_std_logic_vector(624, 16),
13325 => conv_std_logic_vector(676, 16),
13326 => conv_std_logic_vector(728, 16),
13327 => conv_std_logic_vector(780, 16),
13328 => conv_std_logic_vector(832, 16),
13329 => conv_std_logic_vector(884, 16),
13330 => conv_std_logic_vector(936, 16),
13331 => conv_std_logic_vector(988, 16),
13332 => conv_std_logic_vector(1040, 16),
13333 => conv_std_logic_vector(1092, 16),
13334 => conv_std_logic_vector(1144, 16),
13335 => conv_std_logic_vector(1196, 16),
13336 => conv_std_logic_vector(1248, 16),
13337 => conv_std_logic_vector(1300, 16),
13338 => conv_std_logic_vector(1352, 16),
13339 => conv_std_logic_vector(1404, 16),
13340 => conv_std_logic_vector(1456, 16),
13341 => conv_std_logic_vector(1508, 16),
13342 => conv_std_logic_vector(1560, 16),
13343 => conv_std_logic_vector(1612, 16),
13344 => conv_std_logic_vector(1664, 16),
13345 => conv_std_logic_vector(1716, 16),
13346 => conv_std_logic_vector(1768, 16),
13347 => conv_std_logic_vector(1820, 16),
13348 => conv_std_logic_vector(1872, 16),
13349 => conv_std_logic_vector(1924, 16),
13350 => conv_std_logic_vector(1976, 16),
13351 => conv_std_logic_vector(2028, 16),
13352 => conv_std_logic_vector(2080, 16),
13353 => conv_std_logic_vector(2132, 16),
13354 => conv_std_logic_vector(2184, 16),
13355 => conv_std_logic_vector(2236, 16),
13356 => conv_std_logic_vector(2288, 16),
13357 => conv_std_logic_vector(2340, 16),
13358 => conv_std_logic_vector(2392, 16),
13359 => conv_std_logic_vector(2444, 16),
13360 => conv_std_logic_vector(2496, 16),
13361 => conv_std_logic_vector(2548, 16),
13362 => conv_std_logic_vector(2600, 16),
13363 => conv_std_logic_vector(2652, 16),
13364 => conv_std_logic_vector(2704, 16),
13365 => conv_std_logic_vector(2756, 16),
13366 => conv_std_logic_vector(2808, 16),
13367 => conv_std_logic_vector(2860, 16),
13368 => conv_std_logic_vector(2912, 16),
13369 => conv_std_logic_vector(2964, 16),
13370 => conv_std_logic_vector(3016, 16),
13371 => conv_std_logic_vector(3068, 16),
13372 => conv_std_logic_vector(3120, 16),
13373 => conv_std_logic_vector(3172, 16),
13374 => conv_std_logic_vector(3224, 16),
13375 => conv_std_logic_vector(3276, 16),
13376 => conv_std_logic_vector(3328, 16),
13377 => conv_std_logic_vector(3380, 16),
13378 => conv_std_logic_vector(3432, 16),
13379 => conv_std_logic_vector(3484, 16),
13380 => conv_std_logic_vector(3536, 16),
13381 => conv_std_logic_vector(3588, 16),
13382 => conv_std_logic_vector(3640, 16),
13383 => conv_std_logic_vector(3692, 16),
13384 => conv_std_logic_vector(3744, 16),
13385 => conv_std_logic_vector(3796, 16),
13386 => conv_std_logic_vector(3848, 16),
13387 => conv_std_logic_vector(3900, 16),
13388 => conv_std_logic_vector(3952, 16),
13389 => conv_std_logic_vector(4004, 16),
13390 => conv_std_logic_vector(4056, 16),
13391 => conv_std_logic_vector(4108, 16),
13392 => conv_std_logic_vector(4160, 16),
13393 => conv_std_logic_vector(4212, 16),
13394 => conv_std_logic_vector(4264, 16),
13395 => conv_std_logic_vector(4316, 16),
13396 => conv_std_logic_vector(4368, 16),
13397 => conv_std_logic_vector(4420, 16),
13398 => conv_std_logic_vector(4472, 16),
13399 => conv_std_logic_vector(4524, 16),
13400 => conv_std_logic_vector(4576, 16),
13401 => conv_std_logic_vector(4628, 16),
13402 => conv_std_logic_vector(4680, 16),
13403 => conv_std_logic_vector(4732, 16),
13404 => conv_std_logic_vector(4784, 16),
13405 => conv_std_logic_vector(4836, 16),
13406 => conv_std_logic_vector(4888, 16),
13407 => conv_std_logic_vector(4940, 16),
13408 => conv_std_logic_vector(4992, 16),
13409 => conv_std_logic_vector(5044, 16),
13410 => conv_std_logic_vector(5096, 16),
13411 => conv_std_logic_vector(5148, 16),
13412 => conv_std_logic_vector(5200, 16),
13413 => conv_std_logic_vector(5252, 16),
13414 => conv_std_logic_vector(5304, 16),
13415 => conv_std_logic_vector(5356, 16),
13416 => conv_std_logic_vector(5408, 16),
13417 => conv_std_logic_vector(5460, 16),
13418 => conv_std_logic_vector(5512, 16),
13419 => conv_std_logic_vector(5564, 16),
13420 => conv_std_logic_vector(5616, 16),
13421 => conv_std_logic_vector(5668, 16),
13422 => conv_std_logic_vector(5720, 16),
13423 => conv_std_logic_vector(5772, 16),
13424 => conv_std_logic_vector(5824, 16),
13425 => conv_std_logic_vector(5876, 16),
13426 => conv_std_logic_vector(5928, 16),
13427 => conv_std_logic_vector(5980, 16),
13428 => conv_std_logic_vector(6032, 16),
13429 => conv_std_logic_vector(6084, 16),
13430 => conv_std_logic_vector(6136, 16),
13431 => conv_std_logic_vector(6188, 16),
13432 => conv_std_logic_vector(6240, 16),
13433 => conv_std_logic_vector(6292, 16),
13434 => conv_std_logic_vector(6344, 16),
13435 => conv_std_logic_vector(6396, 16),
13436 => conv_std_logic_vector(6448, 16),
13437 => conv_std_logic_vector(6500, 16),
13438 => conv_std_logic_vector(6552, 16),
13439 => conv_std_logic_vector(6604, 16),
13440 => conv_std_logic_vector(6656, 16),
13441 => conv_std_logic_vector(6708, 16),
13442 => conv_std_logic_vector(6760, 16),
13443 => conv_std_logic_vector(6812, 16),
13444 => conv_std_logic_vector(6864, 16),
13445 => conv_std_logic_vector(6916, 16),
13446 => conv_std_logic_vector(6968, 16),
13447 => conv_std_logic_vector(7020, 16),
13448 => conv_std_logic_vector(7072, 16),
13449 => conv_std_logic_vector(7124, 16),
13450 => conv_std_logic_vector(7176, 16),
13451 => conv_std_logic_vector(7228, 16),
13452 => conv_std_logic_vector(7280, 16),
13453 => conv_std_logic_vector(7332, 16),
13454 => conv_std_logic_vector(7384, 16),
13455 => conv_std_logic_vector(7436, 16),
13456 => conv_std_logic_vector(7488, 16),
13457 => conv_std_logic_vector(7540, 16),
13458 => conv_std_logic_vector(7592, 16),
13459 => conv_std_logic_vector(7644, 16),
13460 => conv_std_logic_vector(7696, 16),
13461 => conv_std_logic_vector(7748, 16),
13462 => conv_std_logic_vector(7800, 16),
13463 => conv_std_logic_vector(7852, 16),
13464 => conv_std_logic_vector(7904, 16),
13465 => conv_std_logic_vector(7956, 16),
13466 => conv_std_logic_vector(8008, 16),
13467 => conv_std_logic_vector(8060, 16),
13468 => conv_std_logic_vector(8112, 16),
13469 => conv_std_logic_vector(8164, 16),
13470 => conv_std_logic_vector(8216, 16),
13471 => conv_std_logic_vector(8268, 16),
13472 => conv_std_logic_vector(8320, 16),
13473 => conv_std_logic_vector(8372, 16),
13474 => conv_std_logic_vector(8424, 16),
13475 => conv_std_logic_vector(8476, 16),
13476 => conv_std_logic_vector(8528, 16),
13477 => conv_std_logic_vector(8580, 16),
13478 => conv_std_logic_vector(8632, 16),
13479 => conv_std_logic_vector(8684, 16),
13480 => conv_std_logic_vector(8736, 16),
13481 => conv_std_logic_vector(8788, 16),
13482 => conv_std_logic_vector(8840, 16),
13483 => conv_std_logic_vector(8892, 16),
13484 => conv_std_logic_vector(8944, 16),
13485 => conv_std_logic_vector(8996, 16),
13486 => conv_std_logic_vector(9048, 16),
13487 => conv_std_logic_vector(9100, 16),
13488 => conv_std_logic_vector(9152, 16),
13489 => conv_std_logic_vector(9204, 16),
13490 => conv_std_logic_vector(9256, 16),
13491 => conv_std_logic_vector(9308, 16),
13492 => conv_std_logic_vector(9360, 16),
13493 => conv_std_logic_vector(9412, 16),
13494 => conv_std_logic_vector(9464, 16),
13495 => conv_std_logic_vector(9516, 16),
13496 => conv_std_logic_vector(9568, 16),
13497 => conv_std_logic_vector(9620, 16),
13498 => conv_std_logic_vector(9672, 16),
13499 => conv_std_logic_vector(9724, 16),
13500 => conv_std_logic_vector(9776, 16),
13501 => conv_std_logic_vector(9828, 16),
13502 => conv_std_logic_vector(9880, 16),
13503 => conv_std_logic_vector(9932, 16),
13504 => conv_std_logic_vector(9984, 16),
13505 => conv_std_logic_vector(10036, 16),
13506 => conv_std_logic_vector(10088, 16),
13507 => conv_std_logic_vector(10140, 16),
13508 => conv_std_logic_vector(10192, 16),
13509 => conv_std_logic_vector(10244, 16),
13510 => conv_std_logic_vector(10296, 16),
13511 => conv_std_logic_vector(10348, 16),
13512 => conv_std_logic_vector(10400, 16),
13513 => conv_std_logic_vector(10452, 16),
13514 => conv_std_logic_vector(10504, 16),
13515 => conv_std_logic_vector(10556, 16),
13516 => conv_std_logic_vector(10608, 16),
13517 => conv_std_logic_vector(10660, 16),
13518 => conv_std_logic_vector(10712, 16),
13519 => conv_std_logic_vector(10764, 16),
13520 => conv_std_logic_vector(10816, 16),
13521 => conv_std_logic_vector(10868, 16),
13522 => conv_std_logic_vector(10920, 16),
13523 => conv_std_logic_vector(10972, 16),
13524 => conv_std_logic_vector(11024, 16),
13525 => conv_std_logic_vector(11076, 16),
13526 => conv_std_logic_vector(11128, 16),
13527 => conv_std_logic_vector(11180, 16),
13528 => conv_std_logic_vector(11232, 16),
13529 => conv_std_logic_vector(11284, 16),
13530 => conv_std_logic_vector(11336, 16),
13531 => conv_std_logic_vector(11388, 16),
13532 => conv_std_logic_vector(11440, 16),
13533 => conv_std_logic_vector(11492, 16),
13534 => conv_std_logic_vector(11544, 16),
13535 => conv_std_logic_vector(11596, 16),
13536 => conv_std_logic_vector(11648, 16),
13537 => conv_std_logic_vector(11700, 16),
13538 => conv_std_logic_vector(11752, 16),
13539 => conv_std_logic_vector(11804, 16),
13540 => conv_std_logic_vector(11856, 16),
13541 => conv_std_logic_vector(11908, 16),
13542 => conv_std_logic_vector(11960, 16),
13543 => conv_std_logic_vector(12012, 16),
13544 => conv_std_logic_vector(12064, 16),
13545 => conv_std_logic_vector(12116, 16),
13546 => conv_std_logic_vector(12168, 16),
13547 => conv_std_logic_vector(12220, 16),
13548 => conv_std_logic_vector(12272, 16),
13549 => conv_std_logic_vector(12324, 16),
13550 => conv_std_logic_vector(12376, 16),
13551 => conv_std_logic_vector(12428, 16),
13552 => conv_std_logic_vector(12480, 16),
13553 => conv_std_logic_vector(12532, 16),
13554 => conv_std_logic_vector(12584, 16),
13555 => conv_std_logic_vector(12636, 16),
13556 => conv_std_logic_vector(12688, 16),
13557 => conv_std_logic_vector(12740, 16),
13558 => conv_std_logic_vector(12792, 16),
13559 => conv_std_logic_vector(12844, 16),
13560 => conv_std_logic_vector(12896, 16),
13561 => conv_std_logic_vector(12948, 16),
13562 => conv_std_logic_vector(13000, 16),
13563 => conv_std_logic_vector(13052, 16),
13564 => conv_std_logic_vector(13104, 16),
13565 => conv_std_logic_vector(13156, 16),
13566 => conv_std_logic_vector(13208, 16),
13567 => conv_std_logic_vector(13260, 16),
13568 => conv_std_logic_vector(0, 16),
13569 => conv_std_logic_vector(53, 16),
13570 => conv_std_logic_vector(106, 16),
13571 => conv_std_logic_vector(159, 16),
13572 => conv_std_logic_vector(212, 16),
13573 => conv_std_logic_vector(265, 16),
13574 => conv_std_logic_vector(318, 16),
13575 => conv_std_logic_vector(371, 16),
13576 => conv_std_logic_vector(424, 16),
13577 => conv_std_logic_vector(477, 16),
13578 => conv_std_logic_vector(530, 16),
13579 => conv_std_logic_vector(583, 16),
13580 => conv_std_logic_vector(636, 16),
13581 => conv_std_logic_vector(689, 16),
13582 => conv_std_logic_vector(742, 16),
13583 => conv_std_logic_vector(795, 16),
13584 => conv_std_logic_vector(848, 16),
13585 => conv_std_logic_vector(901, 16),
13586 => conv_std_logic_vector(954, 16),
13587 => conv_std_logic_vector(1007, 16),
13588 => conv_std_logic_vector(1060, 16),
13589 => conv_std_logic_vector(1113, 16),
13590 => conv_std_logic_vector(1166, 16),
13591 => conv_std_logic_vector(1219, 16),
13592 => conv_std_logic_vector(1272, 16),
13593 => conv_std_logic_vector(1325, 16),
13594 => conv_std_logic_vector(1378, 16),
13595 => conv_std_logic_vector(1431, 16),
13596 => conv_std_logic_vector(1484, 16),
13597 => conv_std_logic_vector(1537, 16),
13598 => conv_std_logic_vector(1590, 16),
13599 => conv_std_logic_vector(1643, 16),
13600 => conv_std_logic_vector(1696, 16),
13601 => conv_std_logic_vector(1749, 16),
13602 => conv_std_logic_vector(1802, 16),
13603 => conv_std_logic_vector(1855, 16),
13604 => conv_std_logic_vector(1908, 16),
13605 => conv_std_logic_vector(1961, 16),
13606 => conv_std_logic_vector(2014, 16),
13607 => conv_std_logic_vector(2067, 16),
13608 => conv_std_logic_vector(2120, 16),
13609 => conv_std_logic_vector(2173, 16),
13610 => conv_std_logic_vector(2226, 16),
13611 => conv_std_logic_vector(2279, 16),
13612 => conv_std_logic_vector(2332, 16),
13613 => conv_std_logic_vector(2385, 16),
13614 => conv_std_logic_vector(2438, 16),
13615 => conv_std_logic_vector(2491, 16),
13616 => conv_std_logic_vector(2544, 16),
13617 => conv_std_logic_vector(2597, 16),
13618 => conv_std_logic_vector(2650, 16),
13619 => conv_std_logic_vector(2703, 16),
13620 => conv_std_logic_vector(2756, 16),
13621 => conv_std_logic_vector(2809, 16),
13622 => conv_std_logic_vector(2862, 16),
13623 => conv_std_logic_vector(2915, 16),
13624 => conv_std_logic_vector(2968, 16),
13625 => conv_std_logic_vector(3021, 16),
13626 => conv_std_logic_vector(3074, 16),
13627 => conv_std_logic_vector(3127, 16),
13628 => conv_std_logic_vector(3180, 16),
13629 => conv_std_logic_vector(3233, 16),
13630 => conv_std_logic_vector(3286, 16),
13631 => conv_std_logic_vector(3339, 16),
13632 => conv_std_logic_vector(3392, 16),
13633 => conv_std_logic_vector(3445, 16),
13634 => conv_std_logic_vector(3498, 16),
13635 => conv_std_logic_vector(3551, 16),
13636 => conv_std_logic_vector(3604, 16),
13637 => conv_std_logic_vector(3657, 16),
13638 => conv_std_logic_vector(3710, 16),
13639 => conv_std_logic_vector(3763, 16),
13640 => conv_std_logic_vector(3816, 16),
13641 => conv_std_logic_vector(3869, 16),
13642 => conv_std_logic_vector(3922, 16),
13643 => conv_std_logic_vector(3975, 16),
13644 => conv_std_logic_vector(4028, 16),
13645 => conv_std_logic_vector(4081, 16),
13646 => conv_std_logic_vector(4134, 16),
13647 => conv_std_logic_vector(4187, 16),
13648 => conv_std_logic_vector(4240, 16),
13649 => conv_std_logic_vector(4293, 16),
13650 => conv_std_logic_vector(4346, 16),
13651 => conv_std_logic_vector(4399, 16),
13652 => conv_std_logic_vector(4452, 16),
13653 => conv_std_logic_vector(4505, 16),
13654 => conv_std_logic_vector(4558, 16),
13655 => conv_std_logic_vector(4611, 16),
13656 => conv_std_logic_vector(4664, 16),
13657 => conv_std_logic_vector(4717, 16),
13658 => conv_std_logic_vector(4770, 16),
13659 => conv_std_logic_vector(4823, 16),
13660 => conv_std_logic_vector(4876, 16),
13661 => conv_std_logic_vector(4929, 16),
13662 => conv_std_logic_vector(4982, 16),
13663 => conv_std_logic_vector(5035, 16),
13664 => conv_std_logic_vector(5088, 16),
13665 => conv_std_logic_vector(5141, 16),
13666 => conv_std_logic_vector(5194, 16),
13667 => conv_std_logic_vector(5247, 16),
13668 => conv_std_logic_vector(5300, 16),
13669 => conv_std_logic_vector(5353, 16),
13670 => conv_std_logic_vector(5406, 16),
13671 => conv_std_logic_vector(5459, 16),
13672 => conv_std_logic_vector(5512, 16),
13673 => conv_std_logic_vector(5565, 16),
13674 => conv_std_logic_vector(5618, 16),
13675 => conv_std_logic_vector(5671, 16),
13676 => conv_std_logic_vector(5724, 16),
13677 => conv_std_logic_vector(5777, 16),
13678 => conv_std_logic_vector(5830, 16),
13679 => conv_std_logic_vector(5883, 16),
13680 => conv_std_logic_vector(5936, 16),
13681 => conv_std_logic_vector(5989, 16),
13682 => conv_std_logic_vector(6042, 16),
13683 => conv_std_logic_vector(6095, 16),
13684 => conv_std_logic_vector(6148, 16),
13685 => conv_std_logic_vector(6201, 16),
13686 => conv_std_logic_vector(6254, 16),
13687 => conv_std_logic_vector(6307, 16),
13688 => conv_std_logic_vector(6360, 16),
13689 => conv_std_logic_vector(6413, 16),
13690 => conv_std_logic_vector(6466, 16),
13691 => conv_std_logic_vector(6519, 16),
13692 => conv_std_logic_vector(6572, 16),
13693 => conv_std_logic_vector(6625, 16),
13694 => conv_std_logic_vector(6678, 16),
13695 => conv_std_logic_vector(6731, 16),
13696 => conv_std_logic_vector(6784, 16),
13697 => conv_std_logic_vector(6837, 16),
13698 => conv_std_logic_vector(6890, 16),
13699 => conv_std_logic_vector(6943, 16),
13700 => conv_std_logic_vector(6996, 16),
13701 => conv_std_logic_vector(7049, 16),
13702 => conv_std_logic_vector(7102, 16),
13703 => conv_std_logic_vector(7155, 16),
13704 => conv_std_logic_vector(7208, 16),
13705 => conv_std_logic_vector(7261, 16),
13706 => conv_std_logic_vector(7314, 16),
13707 => conv_std_logic_vector(7367, 16),
13708 => conv_std_logic_vector(7420, 16),
13709 => conv_std_logic_vector(7473, 16),
13710 => conv_std_logic_vector(7526, 16),
13711 => conv_std_logic_vector(7579, 16),
13712 => conv_std_logic_vector(7632, 16),
13713 => conv_std_logic_vector(7685, 16),
13714 => conv_std_logic_vector(7738, 16),
13715 => conv_std_logic_vector(7791, 16),
13716 => conv_std_logic_vector(7844, 16),
13717 => conv_std_logic_vector(7897, 16),
13718 => conv_std_logic_vector(7950, 16),
13719 => conv_std_logic_vector(8003, 16),
13720 => conv_std_logic_vector(8056, 16),
13721 => conv_std_logic_vector(8109, 16),
13722 => conv_std_logic_vector(8162, 16),
13723 => conv_std_logic_vector(8215, 16),
13724 => conv_std_logic_vector(8268, 16),
13725 => conv_std_logic_vector(8321, 16),
13726 => conv_std_logic_vector(8374, 16),
13727 => conv_std_logic_vector(8427, 16),
13728 => conv_std_logic_vector(8480, 16),
13729 => conv_std_logic_vector(8533, 16),
13730 => conv_std_logic_vector(8586, 16),
13731 => conv_std_logic_vector(8639, 16),
13732 => conv_std_logic_vector(8692, 16),
13733 => conv_std_logic_vector(8745, 16),
13734 => conv_std_logic_vector(8798, 16),
13735 => conv_std_logic_vector(8851, 16),
13736 => conv_std_logic_vector(8904, 16),
13737 => conv_std_logic_vector(8957, 16),
13738 => conv_std_logic_vector(9010, 16),
13739 => conv_std_logic_vector(9063, 16),
13740 => conv_std_logic_vector(9116, 16),
13741 => conv_std_logic_vector(9169, 16),
13742 => conv_std_logic_vector(9222, 16),
13743 => conv_std_logic_vector(9275, 16),
13744 => conv_std_logic_vector(9328, 16),
13745 => conv_std_logic_vector(9381, 16),
13746 => conv_std_logic_vector(9434, 16),
13747 => conv_std_logic_vector(9487, 16),
13748 => conv_std_logic_vector(9540, 16),
13749 => conv_std_logic_vector(9593, 16),
13750 => conv_std_logic_vector(9646, 16),
13751 => conv_std_logic_vector(9699, 16),
13752 => conv_std_logic_vector(9752, 16),
13753 => conv_std_logic_vector(9805, 16),
13754 => conv_std_logic_vector(9858, 16),
13755 => conv_std_logic_vector(9911, 16),
13756 => conv_std_logic_vector(9964, 16),
13757 => conv_std_logic_vector(10017, 16),
13758 => conv_std_logic_vector(10070, 16),
13759 => conv_std_logic_vector(10123, 16),
13760 => conv_std_logic_vector(10176, 16),
13761 => conv_std_logic_vector(10229, 16),
13762 => conv_std_logic_vector(10282, 16),
13763 => conv_std_logic_vector(10335, 16),
13764 => conv_std_logic_vector(10388, 16),
13765 => conv_std_logic_vector(10441, 16),
13766 => conv_std_logic_vector(10494, 16),
13767 => conv_std_logic_vector(10547, 16),
13768 => conv_std_logic_vector(10600, 16),
13769 => conv_std_logic_vector(10653, 16),
13770 => conv_std_logic_vector(10706, 16),
13771 => conv_std_logic_vector(10759, 16),
13772 => conv_std_logic_vector(10812, 16),
13773 => conv_std_logic_vector(10865, 16),
13774 => conv_std_logic_vector(10918, 16),
13775 => conv_std_logic_vector(10971, 16),
13776 => conv_std_logic_vector(11024, 16),
13777 => conv_std_logic_vector(11077, 16),
13778 => conv_std_logic_vector(11130, 16),
13779 => conv_std_logic_vector(11183, 16),
13780 => conv_std_logic_vector(11236, 16),
13781 => conv_std_logic_vector(11289, 16),
13782 => conv_std_logic_vector(11342, 16),
13783 => conv_std_logic_vector(11395, 16),
13784 => conv_std_logic_vector(11448, 16),
13785 => conv_std_logic_vector(11501, 16),
13786 => conv_std_logic_vector(11554, 16),
13787 => conv_std_logic_vector(11607, 16),
13788 => conv_std_logic_vector(11660, 16),
13789 => conv_std_logic_vector(11713, 16),
13790 => conv_std_logic_vector(11766, 16),
13791 => conv_std_logic_vector(11819, 16),
13792 => conv_std_logic_vector(11872, 16),
13793 => conv_std_logic_vector(11925, 16),
13794 => conv_std_logic_vector(11978, 16),
13795 => conv_std_logic_vector(12031, 16),
13796 => conv_std_logic_vector(12084, 16),
13797 => conv_std_logic_vector(12137, 16),
13798 => conv_std_logic_vector(12190, 16),
13799 => conv_std_logic_vector(12243, 16),
13800 => conv_std_logic_vector(12296, 16),
13801 => conv_std_logic_vector(12349, 16),
13802 => conv_std_logic_vector(12402, 16),
13803 => conv_std_logic_vector(12455, 16),
13804 => conv_std_logic_vector(12508, 16),
13805 => conv_std_logic_vector(12561, 16),
13806 => conv_std_logic_vector(12614, 16),
13807 => conv_std_logic_vector(12667, 16),
13808 => conv_std_logic_vector(12720, 16),
13809 => conv_std_logic_vector(12773, 16),
13810 => conv_std_logic_vector(12826, 16),
13811 => conv_std_logic_vector(12879, 16),
13812 => conv_std_logic_vector(12932, 16),
13813 => conv_std_logic_vector(12985, 16),
13814 => conv_std_logic_vector(13038, 16),
13815 => conv_std_logic_vector(13091, 16),
13816 => conv_std_logic_vector(13144, 16),
13817 => conv_std_logic_vector(13197, 16),
13818 => conv_std_logic_vector(13250, 16),
13819 => conv_std_logic_vector(13303, 16),
13820 => conv_std_logic_vector(13356, 16),
13821 => conv_std_logic_vector(13409, 16),
13822 => conv_std_logic_vector(13462, 16),
13823 => conv_std_logic_vector(13515, 16),
13824 => conv_std_logic_vector(0, 16),
13825 => conv_std_logic_vector(54, 16),
13826 => conv_std_logic_vector(108, 16),
13827 => conv_std_logic_vector(162, 16),
13828 => conv_std_logic_vector(216, 16),
13829 => conv_std_logic_vector(270, 16),
13830 => conv_std_logic_vector(324, 16),
13831 => conv_std_logic_vector(378, 16),
13832 => conv_std_logic_vector(432, 16),
13833 => conv_std_logic_vector(486, 16),
13834 => conv_std_logic_vector(540, 16),
13835 => conv_std_logic_vector(594, 16),
13836 => conv_std_logic_vector(648, 16),
13837 => conv_std_logic_vector(702, 16),
13838 => conv_std_logic_vector(756, 16),
13839 => conv_std_logic_vector(810, 16),
13840 => conv_std_logic_vector(864, 16),
13841 => conv_std_logic_vector(918, 16),
13842 => conv_std_logic_vector(972, 16),
13843 => conv_std_logic_vector(1026, 16),
13844 => conv_std_logic_vector(1080, 16),
13845 => conv_std_logic_vector(1134, 16),
13846 => conv_std_logic_vector(1188, 16),
13847 => conv_std_logic_vector(1242, 16),
13848 => conv_std_logic_vector(1296, 16),
13849 => conv_std_logic_vector(1350, 16),
13850 => conv_std_logic_vector(1404, 16),
13851 => conv_std_logic_vector(1458, 16),
13852 => conv_std_logic_vector(1512, 16),
13853 => conv_std_logic_vector(1566, 16),
13854 => conv_std_logic_vector(1620, 16),
13855 => conv_std_logic_vector(1674, 16),
13856 => conv_std_logic_vector(1728, 16),
13857 => conv_std_logic_vector(1782, 16),
13858 => conv_std_logic_vector(1836, 16),
13859 => conv_std_logic_vector(1890, 16),
13860 => conv_std_logic_vector(1944, 16),
13861 => conv_std_logic_vector(1998, 16),
13862 => conv_std_logic_vector(2052, 16),
13863 => conv_std_logic_vector(2106, 16),
13864 => conv_std_logic_vector(2160, 16),
13865 => conv_std_logic_vector(2214, 16),
13866 => conv_std_logic_vector(2268, 16),
13867 => conv_std_logic_vector(2322, 16),
13868 => conv_std_logic_vector(2376, 16),
13869 => conv_std_logic_vector(2430, 16),
13870 => conv_std_logic_vector(2484, 16),
13871 => conv_std_logic_vector(2538, 16),
13872 => conv_std_logic_vector(2592, 16),
13873 => conv_std_logic_vector(2646, 16),
13874 => conv_std_logic_vector(2700, 16),
13875 => conv_std_logic_vector(2754, 16),
13876 => conv_std_logic_vector(2808, 16),
13877 => conv_std_logic_vector(2862, 16),
13878 => conv_std_logic_vector(2916, 16),
13879 => conv_std_logic_vector(2970, 16),
13880 => conv_std_logic_vector(3024, 16),
13881 => conv_std_logic_vector(3078, 16),
13882 => conv_std_logic_vector(3132, 16),
13883 => conv_std_logic_vector(3186, 16),
13884 => conv_std_logic_vector(3240, 16),
13885 => conv_std_logic_vector(3294, 16),
13886 => conv_std_logic_vector(3348, 16),
13887 => conv_std_logic_vector(3402, 16),
13888 => conv_std_logic_vector(3456, 16),
13889 => conv_std_logic_vector(3510, 16),
13890 => conv_std_logic_vector(3564, 16),
13891 => conv_std_logic_vector(3618, 16),
13892 => conv_std_logic_vector(3672, 16),
13893 => conv_std_logic_vector(3726, 16),
13894 => conv_std_logic_vector(3780, 16),
13895 => conv_std_logic_vector(3834, 16),
13896 => conv_std_logic_vector(3888, 16),
13897 => conv_std_logic_vector(3942, 16),
13898 => conv_std_logic_vector(3996, 16),
13899 => conv_std_logic_vector(4050, 16),
13900 => conv_std_logic_vector(4104, 16),
13901 => conv_std_logic_vector(4158, 16),
13902 => conv_std_logic_vector(4212, 16),
13903 => conv_std_logic_vector(4266, 16),
13904 => conv_std_logic_vector(4320, 16),
13905 => conv_std_logic_vector(4374, 16),
13906 => conv_std_logic_vector(4428, 16),
13907 => conv_std_logic_vector(4482, 16),
13908 => conv_std_logic_vector(4536, 16),
13909 => conv_std_logic_vector(4590, 16),
13910 => conv_std_logic_vector(4644, 16),
13911 => conv_std_logic_vector(4698, 16),
13912 => conv_std_logic_vector(4752, 16),
13913 => conv_std_logic_vector(4806, 16),
13914 => conv_std_logic_vector(4860, 16),
13915 => conv_std_logic_vector(4914, 16),
13916 => conv_std_logic_vector(4968, 16),
13917 => conv_std_logic_vector(5022, 16),
13918 => conv_std_logic_vector(5076, 16),
13919 => conv_std_logic_vector(5130, 16),
13920 => conv_std_logic_vector(5184, 16),
13921 => conv_std_logic_vector(5238, 16),
13922 => conv_std_logic_vector(5292, 16),
13923 => conv_std_logic_vector(5346, 16),
13924 => conv_std_logic_vector(5400, 16),
13925 => conv_std_logic_vector(5454, 16),
13926 => conv_std_logic_vector(5508, 16),
13927 => conv_std_logic_vector(5562, 16),
13928 => conv_std_logic_vector(5616, 16),
13929 => conv_std_logic_vector(5670, 16),
13930 => conv_std_logic_vector(5724, 16),
13931 => conv_std_logic_vector(5778, 16),
13932 => conv_std_logic_vector(5832, 16),
13933 => conv_std_logic_vector(5886, 16),
13934 => conv_std_logic_vector(5940, 16),
13935 => conv_std_logic_vector(5994, 16),
13936 => conv_std_logic_vector(6048, 16),
13937 => conv_std_logic_vector(6102, 16),
13938 => conv_std_logic_vector(6156, 16),
13939 => conv_std_logic_vector(6210, 16),
13940 => conv_std_logic_vector(6264, 16),
13941 => conv_std_logic_vector(6318, 16),
13942 => conv_std_logic_vector(6372, 16),
13943 => conv_std_logic_vector(6426, 16),
13944 => conv_std_logic_vector(6480, 16),
13945 => conv_std_logic_vector(6534, 16),
13946 => conv_std_logic_vector(6588, 16),
13947 => conv_std_logic_vector(6642, 16),
13948 => conv_std_logic_vector(6696, 16),
13949 => conv_std_logic_vector(6750, 16),
13950 => conv_std_logic_vector(6804, 16),
13951 => conv_std_logic_vector(6858, 16),
13952 => conv_std_logic_vector(6912, 16),
13953 => conv_std_logic_vector(6966, 16),
13954 => conv_std_logic_vector(7020, 16),
13955 => conv_std_logic_vector(7074, 16),
13956 => conv_std_logic_vector(7128, 16),
13957 => conv_std_logic_vector(7182, 16),
13958 => conv_std_logic_vector(7236, 16),
13959 => conv_std_logic_vector(7290, 16),
13960 => conv_std_logic_vector(7344, 16),
13961 => conv_std_logic_vector(7398, 16),
13962 => conv_std_logic_vector(7452, 16),
13963 => conv_std_logic_vector(7506, 16),
13964 => conv_std_logic_vector(7560, 16),
13965 => conv_std_logic_vector(7614, 16),
13966 => conv_std_logic_vector(7668, 16),
13967 => conv_std_logic_vector(7722, 16),
13968 => conv_std_logic_vector(7776, 16),
13969 => conv_std_logic_vector(7830, 16),
13970 => conv_std_logic_vector(7884, 16),
13971 => conv_std_logic_vector(7938, 16),
13972 => conv_std_logic_vector(7992, 16),
13973 => conv_std_logic_vector(8046, 16),
13974 => conv_std_logic_vector(8100, 16),
13975 => conv_std_logic_vector(8154, 16),
13976 => conv_std_logic_vector(8208, 16),
13977 => conv_std_logic_vector(8262, 16),
13978 => conv_std_logic_vector(8316, 16),
13979 => conv_std_logic_vector(8370, 16),
13980 => conv_std_logic_vector(8424, 16),
13981 => conv_std_logic_vector(8478, 16),
13982 => conv_std_logic_vector(8532, 16),
13983 => conv_std_logic_vector(8586, 16),
13984 => conv_std_logic_vector(8640, 16),
13985 => conv_std_logic_vector(8694, 16),
13986 => conv_std_logic_vector(8748, 16),
13987 => conv_std_logic_vector(8802, 16),
13988 => conv_std_logic_vector(8856, 16),
13989 => conv_std_logic_vector(8910, 16),
13990 => conv_std_logic_vector(8964, 16),
13991 => conv_std_logic_vector(9018, 16),
13992 => conv_std_logic_vector(9072, 16),
13993 => conv_std_logic_vector(9126, 16),
13994 => conv_std_logic_vector(9180, 16),
13995 => conv_std_logic_vector(9234, 16),
13996 => conv_std_logic_vector(9288, 16),
13997 => conv_std_logic_vector(9342, 16),
13998 => conv_std_logic_vector(9396, 16),
13999 => conv_std_logic_vector(9450, 16),
14000 => conv_std_logic_vector(9504, 16),
14001 => conv_std_logic_vector(9558, 16),
14002 => conv_std_logic_vector(9612, 16),
14003 => conv_std_logic_vector(9666, 16),
14004 => conv_std_logic_vector(9720, 16),
14005 => conv_std_logic_vector(9774, 16),
14006 => conv_std_logic_vector(9828, 16),
14007 => conv_std_logic_vector(9882, 16),
14008 => conv_std_logic_vector(9936, 16),
14009 => conv_std_logic_vector(9990, 16),
14010 => conv_std_logic_vector(10044, 16),
14011 => conv_std_logic_vector(10098, 16),
14012 => conv_std_logic_vector(10152, 16),
14013 => conv_std_logic_vector(10206, 16),
14014 => conv_std_logic_vector(10260, 16),
14015 => conv_std_logic_vector(10314, 16),
14016 => conv_std_logic_vector(10368, 16),
14017 => conv_std_logic_vector(10422, 16),
14018 => conv_std_logic_vector(10476, 16),
14019 => conv_std_logic_vector(10530, 16),
14020 => conv_std_logic_vector(10584, 16),
14021 => conv_std_logic_vector(10638, 16),
14022 => conv_std_logic_vector(10692, 16),
14023 => conv_std_logic_vector(10746, 16),
14024 => conv_std_logic_vector(10800, 16),
14025 => conv_std_logic_vector(10854, 16),
14026 => conv_std_logic_vector(10908, 16),
14027 => conv_std_logic_vector(10962, 16),
14028 => conv_std_logic_vector(11016, 16),
14029 => conv_std_logic_vector(11070, 16),
14030 => conv_std_logic_vector(11124, 16),
14031 => conv_std_logic_vector(11178, 16),
14032 => conv_std_logic_vector(11232, 16),
14033 => conv_std_logic_vector(11286, 16),
14034 => conv_std_logic_vector(11340, 16),
14035 => conv_std_logic_vector(11394, 16),
14036 => conv_std_logic_vector(11448, 16),
14037 => conv_std_logic_vector(11502, 16),
14038 => conv_std_logic_vector(11556, 16),
14039 => conv_std_logic_vector(11610, 16),
14040 => conv_std_logic_vector(11664, 16),
14041 => conv_std_logic_vector(11718, 16),
14042 => conv_std_logic_vector(11772, 16),
14043 => conv_std_logic_vector(11826, 16),
14044 => conv_std_logic_vector(11880, 16),
14045 => conv_std_logic_vector(11934, 16),
14046 => conv_std_logic_vector(11988, 16),
14047 => conv_std_logic_vector(12042, 16),
14048 => conv_std_logic_vector(12096, 16),
14049 => conv_std_logic_vector(12150, 16),
14050 => conv_std_logic_vector(12204, 16),
14051 => conv_std_logic_vector(12258, 16),
14052 => conv_std_logic_vector(12312, 16),
14053 => conv_std_logic_vector(12366, 16),
14054 => conv_std_logic_vector(12420, 16),
14055 => conv_std_logic_vector(12474, 16),
14056 => conv_std_logic_vector(12528, 16),
14057 => conv_std_logic_vector(12582, 16),
14058 => conv_std_logic_vector(12636, 16),
14059 => conv_std_logic_vector(12690, 16),
14060 => conv_std_logic_vector(12744, 16),
14061 => conv_std_logic_vector(12798, 16),
14062 => conv_std_logic_vector(12852, 16),
14063 => conv_std_logic_vector(12906, 16),
14064 => conv_std_logic_vector(12960, 16),
14065 => conv_std_logic_vector(13014, 16),
14066 => conv_std_logic_vector(13068, 16),
14067 => conv_std_logic_vector(13122, 16),
14068 => conv_std_logic_vector(13176, 16),
14069 => conv_std_logic_vector(13230, 16),
14070 => conv_std_logic_vector(13284, 16),
14071 => conv_std_logic_vector(13338, 16),
14072 => conv_std_logic_vector(13392, 16),
14073 => conv_std_logic_vector(13446, 16),
14074 => conv_std_logic_vector(13500, 16),
14075 => conv_std_logic_vector(13554, 16),
14076 => conv_std_logic_vector(13608, 16),
14077 => conv_std_logic_vector(13662, 16),
14078 => conv_std_logic_vector(13716, 16),
14079 => conv_std_logic_vector(13770, 16),
14080 => conv_std_logic_vector(0, 16),
14081 => conv_std_logic_vector(55, 16),
14082 => conv_std_logic_vector(110, 16),
14083 => conv_std_logic_vector(165, 16),
14084 => conv_std_logic_vector(220, 16),
14085 => conv_std_logic_vector(275, 16),
14086 => conv_std_logic_vector(330, 16),
14087 => conv_std_logic_vector(385, 16),
14088 => conv_std_logic_vector(440, 16),
14089 => conv_std_logic_vector(495, 16),
14090 => conv_std_logic_vector(550, 16),
14091 => conv_std_logic_vector(605, 16),
14092 => conv_std_logic_vector(660, 16),
14093 => conv_std_logic_vector(715, 16),
14094 => conv_std_logic_vector(770, 16),
14095 => conv_std_logic_vector(825, 16),
14096 => conv_std_logic_vector(880, 16),
14097 => conv_std_logic_vector(935, 16),
14098 => conv_std_logic_vector(990, 16),
14099 => conv_std_logic_vector(1045, 16),
14100 => conv_std_logic_vector(1100, 16),
14101 => conv_std_logic_vector(1155, 16),
14102 => conv_std_logic_vector(1210, 16),
14103 => conv_std_logic_vector(1265, 16),
14104 => conv_std_logic_vector(1320, 16),
14105 => conv_std_logic_vector(1375, 16),
14106 => conv_std_logic_vector(1430, 16),
14107 => conv_std_logic_vector(1485, 16),
14108 => conv_std_logic_vector(1540, 16),
14109 => conv_std_logic_vector(1595, 16),
14110 => conv_std_logic_vector(1650, 16),
14111 => conv_std_logic_vector(1705, 16),
14112 => conv_std_logic_vector(1760, 16),
14113 => conv_std_logic_vector(1815, 16),
14114 => conv_std_logic_vector(1870, 16),
14115 => conv_std_logic_vector(1925, 16),
14116 => conv_std_logic_vector(1980, 16),
14117 => conv_std_logic_vector(2035, 16),
14118 => conv_std_logic_vector(2090, 16),
14119 => conv_std_logic_vector(2145, 16),
14120 => conv_std_logic_vector(2200, 16),
14121 => conv_std_logic_vector(2255, 16),
14122 => conv_std_logic_vector(2310, 16),
14123 => conv_std_logic_vector(2365, 16),
14124 => conv_std_logic_vector(2420, 16),
14125 => conv_std_logic_vector(2475, 16),
14126 => conv_std_logic_vector(2530, 16),
14127 => conv_std_logic_vector(2585, 16),
14128 => conv_std_logic_vector(2640, 16),
14129 => conv_std_logic_vector(2695, 16),
14130 => conv_std_logic_vector(2750, 16),
14131 => conv_std_logic_vector(2805, 16),
14132 => conv_std_logic_vector(2860, 16),
14133 => conv_std_logic_vector(2915, 16),
14134 => conv_std_logic_vector(2970, 16),
14135 => conv_std_logic_vector(3025, 16),
14136 => conv_std_logic_vector(3080, 16),
14137 => conv_std_logic_vector(3135, 16),
14138 => conv_std_logic_vector(3190, 16),
14139 => conv_std_logic_vector(3245, 16),
14140 => conv_std_logic_vector(3300, 16),
14141 => conv_std_logic_vector(3355, 16),
14142 => conv_std_logic_vector(3410, 16),
14143 => conv_std_logic_vector(3465, 16),
14144 => conv_std_logic_vector(3520, 16),
14145 => conv_std_logic_vector(3575, 16),
14146 => conv_std_logic_vector(3630, 16),
14147 => conv_std_logic_vector(3685, 16),
14148 => conv_std_logic_vector(3740, 16),
14149 => conv_std_logic_vector(3795, 16),
14150 => conv_std_logic_vector(3850, 16),
14151 => conv_std_logic_vector(3905, 16),
14152 => conv_std_logic_vector(3960, 16),
14153 => conv_std_logic_vector(4015, 16),
14154 => conv_std_logic_vector(4070, 16),
14155 => conv_std_logic_vector(4125, 16),
14156 => conv_std_logic_vector(4180, 16),
14157 => conv_std_logic_vector(4235, 16),
14158 => conv_std_logic_vector(4290, 16),
14159 => conv_std_logic_vector(4345, 16),
14160 => conv_std_logic_vector(4400, 16),
14161 => conv_std_logic_vector(4455, 16),
14162 => conv_std_logic_vector(4510, 16),
14163 => conv_std_logic_vector(4565, 16),
14164 => conv_std_logic_vector(4620, 16),
14165 => conv_std_logic_vector(4675, 16),
14166 => conv_std_logic_vector(4730, 16),
14167 => conv_std_logic_vector(4785, 16),
14168 => conv_std_logic_vector(4840, 16),
14169 => conv_std_logic_vector(4895, 16),
14170 => conv_std_logic_vector(4950, 16),
14171 => conv_std_logic_vector(5005, 16),
14172 => conv_std_logic_vector(5060, 16),
14173 => conv_std_logic_vector(5115, 16),
14174 => conv_std_logic_vector(5170, 16),
14175 => conv_std_logic_vector(5225, 16),
14176 => conv_std_logic_vector(5280, 16),
14177 => conv_std_logic_vector(5335, 16),
14178 => conv_std_logic_vector(5390, 16),
14179 => conv_std_logic_vector(5445, 16),
14180 => conv_std_logic_vector(5500, 16),
14181 => conv_std_logic_vector(5555, 16),
14182 => conv_std_logic_vector(5610, 16),
14183 => conv_std_logic_vector(5665, 16),
14184 => conv_std_logic_vector(5720, 16),
14185 => conv_std_logic_vector(5775, 16),
14186 => conv_std_logic_vector(5830, 16),
14187 => conv_std_logic_vector(5885, 16),
14188 => conv_std_logic_vector(5940, 16),
14189 => conv_std_logic_vector(5995, 16),
14190 => conv_std_logic_vector(6050, 16),
14191 => conv_std_logic_vector(6105, 16),
14192 => conv_std_logic_vector(6160, 16),
14193 => conv_std_logic_vector(6215, 16),
14194 => conv_std_logic_vector(6270, 16),
14195 => conv_std_logic_vector(6325, 16),
14196 => conv_std_logic_vector(6380, 16),
14197 => conv_std_logic_vector(6435, 16),
14198 => conv_std_logic_vector(6490, 16),
14199 => conv_std_logic_vector(6545, 16),
14200 => conv_std_logic_vector(6600, 16),
14201 => conv_std_logic_vector(6655, 16),
14202 => conv_std_logic_vector(6710, 16),
14203 => conv_std_logic_vector(6765, 16),
14204 => conv_std_logic_vector(6820, 16),
14205 => conv_std_logic_vector(6875, 16),
14206 => conv_std_logic_vector(6930, 16),
14207 => conv_std_logic_vector(6985, 16),
14208 => conv_std_logic_vector(7040, 16),
14209 => conv_std_logic_vector(7095, 16),
14210 => conv_std_logic_vector(7150, 16),
14211 => conv_std_logic_vector(7205, 16),
14212 => conv_std_logic_vector(7260, 16),
14213 => conv_std_logic_vector(7315, 16),
14214 => conv_std_logic_vector(7370, 16),
14215 => conv_std_logic_vector(7425, 16),
14216 => conv_std_logic_vector(7480, 16),
14217 => conv_std_logic_vector(7535, 16),
14218 => conv_std_logic_vector(7590, 16),
14219 => conv_std_logic_vector(7645, 16),
14220 => conv_std_logic_vector(7700, 16),
14221 => conv_std_logic_vector(7755, 16),
14222 => conv_std_logic_vector(7810, 16),
14223 => conv_std_logic_vector(7865, 16),
14224 => conv_std_logic_vector(7920, 16),
14225 => conv_std_logic_vector(7975, 16),
14226 => conv_std_logic_vector(8030, 16),
14227 => conv_std_logic_vector(8085, 16),
14228 => conv_std_logic_vector(8140, 16),
14229 => conv_std_logic_vector(8195, 16),
14230 => conv_std_logic_vector(8250, 16),
14231 => conv_std_logic_vector(8305, 16),
14232 => conv_std_logic_vector(8360, 16),
14233 => conv_std_logic_vector(8415, 16),
14234 => conv_std_logic_vector(8470, 16),
14235 => conv_std_logic_vector(8525, 16),
14236 => conv_std_logic_vector(8580, 16),
14237 => conv_std_logic_vector(8635, 16),
14238 => conv_std_logic_vector(8690, 16),
14239 => conv_std_logic_vector(8745, 16),
14240 => conv_std_logic_vector(8800, 16),
14241 => conv_std_logic_vector(8855, 16),
14242 => conv_std_logic_vector(8910, 16),
14243 => conv_std_logic_vector(8965, 16),
14244 => conv_std_logic_vector(9020, 16),
14245 => conv_std_logic_vector(9075, 16),
14246 => conv_std_logic_vector(9130, 16),
14247 => conv_std_logic_vector(9185, 16),
14248 => conv_std_logic_vector(9240, 16),
14249 => conv_std_logic_vector(9295, 16),
14250 => conv_std_logic_vector(9350, 16),
14251 => conv_std_logic_vector(9405, 16),
14252 => conv_std_logic_vector(9460, 16),
14253 => conv_std_logic_vector(9515, 16),
14254 => conv_std_logic_vector(9570, 16),
14255 => conv_std_logic_vector(9625, 16),
14256 => conv_std_logic_vector(9680, 16),
14257 => conv_std_logic_vector(9735, 16),
14258 => conv_std_logic_vector(9790, 16),
14259 => conv_std_logic_vector(9845, 16),
14260 => conv_std_logic_vector(9900, 16),
14261 => conv_std_logic_vector(9955, 16),
14262 => conv_std_logic_vector(10010, 16),
14263 => conv_std_logic_vector(10065, 16),
14264 => conv_std_logic_vector(10120, 16),
14265 => conv_std_logic_vector(10175, 16),
14266 => conv_std_logic_vector(10230, 16),
14267 => conv_std_logic_vector(10285, 16),
14268 => conv_std_logic_vector(10340, 16),
14269 => conv_std_logic_vector(10395, 16),
14270 => conv_std_logic_vector(10450, 16),
14271 => conv_std_logic_vector(10505, 16),
14272 => conv_std_logic_vector(10560, 16),
14273 => conv_std_logic_vector(10615, 16),
14274 => conv_std_logic_vector(10670, 16),
14275 => conv_std_logic_vector(10725, 16),
14276 => conv_std_logic_vector(10780, 16),
14277 => conv_std_logic_vector(10835, 16),
14278 => conv_std_logic_vector(10890, 16),
14279 => conv_std_logic_vector(10945, 16),
14280 => conv_std_logic_vector(11000, 16),
14281 => conv_std_logic_vector(11055, 16),
14282 => conv_std_logic_vector(11110, 16),
14283 => conv_std_logic_vector(11165, 16),
14284 => conv_std_logic_vector(11220, 16),
14285 => conv_std_logic_vector(11275, 16),
14286 => conv_std_logic_vector(11330, 16),
14287 => conv_std_logic_vector(11385, 16),
14288 => conv_std_logic_vector(11440, 16),
14289 => conv_std_logic_vector(11495, 16),
14290 => conv_std_logic_vector(11550, 16),
14291 => conv_std_logic_vector(11605, 16),
14292 => conv_std_logic_vector(11660, 16),
14293 => conv_std_logic_vector(11715, 16),
14294 => conv_std_logic_vector(11770, 16),
14295 => conv_std_logic_vector(11825, 16),
14296 => conv_std_logic_vector(11880, 16),
14297 => conv_std_logic_vector(11935, 16),
14298 => conv_std_logic_vector(11990, 16),
14299 => conv_std_logic_vector(12045, 16),
14300 => conv_std_logic_vector(12100, 16),
14301 => conv_std_logic_vector(12155, 16),
14302 => conv_std_logic_vector(12210, 16),
14303 => conv_std_logic_vector(12265, 16),
14304 => conv_std_logic_vector(12320, 16),
14305 => conv_std_logic_vector(12375, 16),
14306 => conv_std_logic_vector(12430, 16),
14307 => conv_std_logic_vector(12485, 16),
14308 => conv_std_logic_vector(12540, 16),
14309 => conv_std_logic_vector(12595, 16),
14310 => conv_std_logic_vector(12650, 16),
14311 => conv_std_logic_vector(12705, 16),
14312 => conv_std_logic_vector(12760, 16),
14313 => conv_std_logic_vector(12815, 16),
14314 => conv_std_logic_vector(12870, 16),
14315 => conv_std_logic_vector(12925, 16),
14316 => conv_std_logic_vector(12980, 16),
14317 => conv_std_logic_vector(13035, 16),
14318 => conv_std_logic_vector(13090, 16),
14319 => conv_std_logic_vector(13145, 16),
14320 => conv_std_logic_vector(13200, 16),
14321 => conv_std_logic_vector(13255, 16),
14322 => conv_std_logic_vector(13310, 16),
14323 => conv_std_logic_vector(13365, 16),
14324 => conv_std_logic_vector(13420, 16),
14325 => conv_std_logic_vector(13475, 16),
14326 => conv_std_logic_vector(13530, 16),
14327 => conv_std_logic_vector(13585, 16),
14328 => conv_std_logic_vector(13640, 16),
14329 => conv_std_logic_vector(13695, 16),
14330 => conv_std_logic_vector(13750, 16),
14331 => conv_std_logic_vector(13805, 16),
14332 => conv_std_logic_vector(13860, 16),
14333 => conv_std_logic_vector(13915, 16),
14334 => conv_std_logic_vector(13970, 16),
14335 => conv_std_logic_vector(14025, 16),
14336 => conv_std_logic_vector(0, 16),
14337 => conv_std_logic_vector(56, 16),
14338 => conv_std_logic_vector(112, 16),
14339 => conv_std_logic_vector(168, 16),
14340 => conv_std_logic_vector(224, 16),
14341 => conv_std_logic_vector(280, 16),
14342 => conv_std_logic_vector(336, 16),
14343 => conv_std_logic_vector(392, 16),
14344 => conv_std_logic_vector(448, 16),
14345 => conv_std_logic_vector(504, 16),
14346 => conv_std_logic_vector(560, 16),
14347 => conv_std_logic_vector(616, 16),
14348 => conv_std_logic_vector(672, 16),
14349 => conv_std_logic_vector(728, 16),
14350 => conv_std_logic_vector(784, 16),
14351 => conv_std_logic_vector(840, 16),
14352 => conv_std_logic_vector(896, 16),
14353 => conv_std_logic_vector(952, 16),
14354 => conv_std_logic_vector(1008, 16),
14355 => conv_std_logic_vector(1064, 16),
14356 => conv_std_logic_vector(1120, 16),
14357 => conv_std_logic_vector(1176, 16),
14358 => conv_std_logic_vector(1232, 16),
14359 => conv_std_logic_vector(1288, 16),
14360 => conv_std_logic_vector(1344, 16),
14361 => conv_std_logic_vector(1400, 16),
14362 => conv_std_logic_vector(1456, 16),
14363 => conv_std_logic_vector(1512, 16),
14364 => conv_std_logic_vector(1568, 16),
14365 => conv_std_logic_vector(1624, 16),
14366 => conv_std_logic_vector(1680, 16),
14367 => conv_std_logic_vector(1736, 16),
14368 => conv_std_logic_vector(1792, 16),
14369 => conv_std_logic_vector(1848, 16),
14370 => conv_std_logic_vector(1904, 16),
14371 => conv_std_logic_vector(1960, 16),
14372 => conv_std_logic_vector(2016, 16),
14373 => conv_std_logic_vector(2072, 16),
14374 => conv_std_logic_vector(2128, 16),
14375 => conv_std_logic_vector(2184, 16),
14376 => conv_std_logic_vector(2240, 16),
14377 => conv_std_logic_vector(2296, 16),
14378 => conv_std_logic_vector(2352, 16),
14379 => conv_std_logic_vector(2408, 16),
14380 => conv_std_logic_vector(2464, 16),
14381 => conv_std_logic_vector(2520, 16),
14382 => conv_std_logic_vector(2576, 16),
14383 => conv_std_logic_vector(2632, 16),
14384 => conv_std_logic_vector(2688, 16),
14385 => conv_std_logic_vector(2744, 16),
14386 => conv_std_logic_vector(2800, 16),
14387 => conv_std_logic_vector(2856, 16),
14388 => conv_std_logic_vector(2912, 16),
14389 => conv_std_logic_vector(2968, 16),
14390 => conv_std_logic_vector(3024, 16),
14391 => conv_std_logic_vector(3080, 16),
14392 => conv_std_logic_vector(3136, 16),
14393 => conv_std_logic_vector(3192, 16),
14394 => conv_std_logic_vector(3248, 16),
14395 => conv_std_logic_vector(3304, 16),
14396 => conv_std_logic_vector(3360, 16),
14397 => conv_std_logic_vector(3416, 16),
14398 => conv_std_logic_vector(3472, 16),
14399 => conv_std_logic_vector(3528, 16),
14400 => conv_std_logic_vector(3584, 16),
14401 => conv_std_logic_vector(3640, 16),
14402 => conv_std_logic_vector(3696, 16),
14403 => conv_std_logic_vector(3752, 16),
14404 => conv_std_logic_vector(3808, 16),
14405 => conv_std_logic_vector(3864, 16),
14406 => conv_std_logic_vector(3920, 16),
14407 => conv_std_logic_vector(3976, 16),
14408 => conv_std_logic_vector(4032, 16),
14409 => conv_std_logic_vector(4088, 16),
14410 => conv_std_logic_vector(4144, 16),
14411 => conv_std_logic_vector(4200, 16),
14412 => conv_std_logic_vector(4256, 16),
14413 => conv_std_logic_vector(4312, 16),
14414 => conv_std_logic_vector(4368, 16),
14415 => conv_std_logic_vector(4424, 16),
14416 => conv_std_logic_vector(4480, 16),
14417 => conv_std_logic_vector(4536, 16),
14418 => conv_std_logic_vector(4592, 16),
14419 => conv_std_logic_vector(4648, 16),
14420 => conv_std_logic_vector(4704, 16),
14421 => conv_std_logic_vector(4760, 16),
14422 => conv_std_logic_vector(4816, 16),
14423 => conv_std_logic_vector(4872, 16),
14424 => conv_std_logic_vector(4928, 16),
14425 => conv_std_logic_vector(4984, 16),
14426 => conv_std_logic_vector(5040, 16),
14427 => conv_std_logic_vector(5096, 16),
14428 => conv_std_logic_vector(5152, 16),
14429 => conv_std_logic_vector(5208, 16),
14430 => conv_std_logic_vector(5264, 16),
14431 => conv_std_logic_vector(5320, 16),
14432 => conv_std_logic_vector(5376, 16),
14433 => conv_std_logic_vector(5432, 16),
14434 => conv_std_logic_vector(5488, 16),
14435 => conv_std_logic_vector(5544, 16),
14436 => conv_std_logic_vector(5600, 16),
14437 => conv_std_logic_vector(5656, 16),
14438 => conv_std_logic_vector(5712, 16),
14439 => conv_std_logic_vector(5768, 16),
14440 => conv_std_logic_vector(5824, 16),
14441 => conv_std_logic_vector(5880, 16),
14442 => conv_std_logic_vector(5936, 16),
14443 => conv_std_logic_vector(5992, 16),
14444 => conv_std_logic_vector(6048, 16),
14445 => conv_std_logic_vector(6104, 16),
14446 => conv_std_logic_vector(6160, 16),
14447 => conv_std_logic_vector(6216, 16),
14448 => conv_std_logic_vector(6272, 16),
14449 => conv_std_logic_vector(6328, 16),
14450 => conv_std_logic_vector(6384, 16),
14451 => conv_std_logic_vector(6440, 16),
14452 => conv_std_logic_vector(6496, 16),
14453 => conv_std_logic_vector(6552, 16),
14454 => conv_std_logic_vector(6608, 16),
14455 => conv_std_logic_vector(6664, 16),
14456 => conv_std_logic_vector(6720, 16),
14457 => conv_std_logic_vector(6776, 16),
14458 => conv_std_logic_vector(6832, 16),
14459 => conv_std_logic_vector(6888, 16),
14460 => conv_std_logic_vector(6944, 16),
14461 => conv_std_logic_vector(7000, 16),
14462 => conv_std_logic_vector(7056, 16),
14463 => conv_std_logic_vector(7112, 16),
14464 => conv_std_logic_vector(7168, 16),
14465 => conv_std_logic_vector(7224, 16),
14466 => conv_std_logic_vector(7280, 16),
14467 => conv_std_logic_vector(7336, 16),
14468 => conv_std_logic_vector(7392, 16),
14469 => conv_std_logic_vector(7448, 16),
14470 => conv_std_logic_vector(7504, 16),
14471 => conv_std_logic_vector(7560, 16),
14472 => conv_std_logic_vector(7616, 16),
14473 => conv_std_logic_vector(7672, 16),
14474 => conv_std_logic_vector(7728, 16),
14475 => conv_std_logic_vector(7784, 16),
14476 => conv_std_logic_vector(7840, 16),
14477 => conv_std_logic_vector(7896, 16),
14478 => conv_std_logic_vector(7952, 16),
14479 => conv_std_logic_vector(8008, 16),
14480 => conv_std_logic_vector(8064, 16),
14481 => conv_std_logic_vector(8120, 16),
14482 => conv_std_logic_vector(8176, 16),
14483 => conv_std_logic_vector(8232, 16),
14484 => conv_std_logic_vector(8288, 16),
14485 => conv_std_logic_vector(8344, 16),
14486 => conv_std_logic_vector(8400, 16),
14487 => conv_std_logic_vector(8456, 16),
14488 => conv_std_logic_vector(8512, 16),
14489 => conv_std_logic_vector(8568, 16),
14490 => conv_std_logic_vector(8624, 16),
14491 => conv_std_logic_vector(8680, 16),
14492 => conv_std_logic_vector(8736, 16),
14493 => conv_std_logic_vector(8792, 16),
14494 => conv_std_logic_vector(8848, 16),
14495 => conv_std_logic_vector(8904, 16),
14496 => conv_std_logic_vector(8960, 16),
14497 => conv_std_logic_vector(9016, 16),
14498 => conv_std_logic_vector(9072, 16),
14499 => conv_std_logic_vector(9128, 16),
14500 => conv_std_logic_vector(9184, 16),
14501 => conv_std_logic_vector(9240, 16),
14502 => conv_std_logic_vector(9296, 16),
14503 => conv_std_logic_vector(9352, 16),
14504 => conv_std_logic_vector(9408, 16),
14505 => conv_std_logic_vector(9464, 16),
14506 => conv_std_logic_vector(9520, 16),
14507 => conv_std_logic_vector(9576, 16),
14508 => conv_std_logic_vector(9632, 16),
14509 => conv_std_logic_vector(9688, 16),
14510 => conv_std_logic_vector(9744, 16),
14511 => conv_std_logic_vector(9800, 16),
14512 => conv_std_logic_vector(9856, 16),
14513 => conv_std_logic_vector(9912, 16),
14514 => conv_std_logic_vector(9968, 16),
14515 => conv_std_logic_vector(10024, 16),
14516 => conv_std_logic_vector(10080, 16),
14517 => conv_std_logic_vector(10136, 16),
14518 => conv_std_logic_vector(10192, 16),
14519 => conv_std_logic_vector(10248, 16),
14520 => conv_std_logic_vector(10304, 16),
14521 => conv_std_logic_vector(10360, 16),
14522 => conv_std_logic_vector(10416, 16),
14523 => conv_std_logic_vector(10472, 16),
14524 => conv_std_logic_vector(10528, 16),
14525 => conv_std_logic_vector(10584, 16),
14526 => conv_std_logic_vector(10640, 16),
14527 => conv_std_logic_vector(10696, 16),
14528 => conv_std_logic_vector(10752, 16),
14529 => conv_std_logic_vector(10808, 16),
14530 => conv_std_logic_vector(10864, 16),
14531 => conv_std_logic_vector(10920, 16),
14532 => conv_std_logic_vector(10976, 16),
14533 => conv_std_logic_vector(11032, 16),
14534 => conv_std_logic_vector(11088, 16),
14535 => conv_std_logic_vector(11144, 16),
14536 => conv_std_logic_vector(11200, 16),
14537 => conv_std_logic_vector(11256, 16),
14538 => conv_std_logic_vector(11312, 16),
14539 => conv_std_logic_vector(11368, 16),
14540 => conv_std_logic_vector(11424, 16),
14541 => conv_std_logic_vector(11480, 16),
14542 => conv_std_logic_vector(11536, 16),
14543 => conv_std_logic_vector(11592, 16),
14544 => conv_std_logic_vector(11648, 16),
14545 => conv_std_logic_vector(11704, 16),
14546 => conv_std_logic_vector(11760, 16),
14547 => conv_std_logic_vector(11816, 16),
14548 => conv_std_logic_vector(11872, 16),
14549 => conv_std_logic_vector(11928, 16),
14550 => conv_std_logic_vector(11984, 16),
14551 => conv_std_logic_vector(12040, 16),
14552 => conv_std_logic_vector(12096, 16),
14553 => conv_std_logic_vector(12152, 16),
14554 => conv_std_logic_vector(12208, 16),
14555 => conv_std_logic_vector(12264, 16),
14556 => conv_std_logic_vector(12320, 16),
14557 => conv_std_logic_vector(12376, 16),
14558 => conv_std_logic_vector(12432, 16),
14559 => conv_std_logic_vector(12488, 16),
14560 => conv_std_logic_vector(12544, 16),
14561 => conv_std_logic_vector(12600, 16),
14562 => conv_std_logic_vector(12656, 16),
14563 => conv_std_logic_vector(12712, 16),
14564 => conv_std_logic_vector(12768, 16),
14565 => conv_std_logic_vector(12824, 16),
14566 => conv_std_logic_vector(12880, 16),
14567 => conv_std_logic_vector(12936, 16),
14568 => conv_std_logic_vector(12992, 16),
14569 => conv_std_logic_vector(13048, 16),
14570 => conv_std_logic_vector(13104, 16),
14571 => conv_std_logic_vector(13160, 16),
14572 => conv_std_logic_vector(13216, 16),
14573 => conv_std_logic_vector(13272, 16),
14574 => conv_std_logic_vector(13328, 16),
14575 => conv_std_logic_vector(13384, 16),
14576 => conv_std_logic_vector(13440, 16),
14577 => conv_std_logic_vector(13496, 16),
14578 => conv_std_logic_vector(13552, 16),
14579 => conv_std_logic_vector(13608, 16),
14580 => conv_std_logic_vector(13664, 16),
14581 => conv_std_logic_vector(13720, 16),
14582 => conv_std_logic_vector(13776, 16),
14583 => conv_std_logic_vector(13832, 16),
14584 => conv_std_logic_vector(13888, 16),
14585 => conv_std_logic_vector(13944, 16),
14586 => conv_std_logic_vector(14000, 16),
14587 => conv_std_logic_vector(14056, 16),
14588 => conv_std_logic_vector(14112, 16),
14589 => conv_std_logic_vector(14168, 16),
14590 => conv_std_logic_vector(14224, 16),
14591 => conv_std_logic_vector(14280, 16),
14592 => conv_std_logic_vector(0, 16),
14593 => conv_std_logic_vector(57, 16),
14594 => conv_std_logic_vector(114, 16),
14595 => conv_std_logic_vector(171, 16),
14596 => conv_std_logic_vector(228, 16),
14597 => conv_std_logic_vector(285, 16),
14598 => conv_std_logic_vector(342, 16),
14599 => conv_std_logic_vector(399, 16),
14600 => conv_std_logic_vector(456, 16),
14601 => conv_std_logic_vector(513, 16),
14602 => conv_std_logic_vector(570, 16),
14603 => conv_std_logic_vector(627, 16),
14604 => conv_std_logic_vector(684, 16),
14605 => conv_std_logic_vector(741, 16),
14606 => conv_std_logic_vector(798, 16),
14607 => conv_std_logic_vector(855, 16),
14608 => conv_std_logic_vector(912, 16),
14609 => conv_std_logic_vector(969, 16),
14610 => conv_std_logic_vector(1026, 16),
14611 => conv_std_logic_vector(1083, 16),
14612 => conv_std_logic_vector(1140, 16),
14613 => conv_std_logic_vector(1197, 16),
14614 => conv_std_logic_vector(1254, 16),
14615 => conv_std_logic_vector(1311, 16),
14616 => conv_std_logic_vector(1368, 16),
14617 => conv_std_logic_vector(1425, 16),
14618 => conv_std_logic_vector(1482, 16),
14619 => conv_std_logic_vector(1539, 16),
14620 => conv_std_logic_vector(1596, 16),
14621 => conv_std_logic_vector(1653, 16),
14622 => conv_std_logic_vector(1710, 16),
14623 => conv_std_logic_vector(1767, 16),
14624 => conv_std_logic_vector(1824, 16),
14625 => conv_std_logic_vector(1881, 16),
14626 => conv_std_logic_vector(1938, 16),
14627 => conv_std_logic_vector(1995, 16),
14628 => conv_std_logic_vector(2052, 16),
14629 => conv_std_logic_vector(2109, 16),
14630 => conv_std_logic_vector(2166, 16),
14631 => conv_std_logic_vector(2223, 16),
14632 => conv_std_logic_vector(2280, 16),
14633 => conv_std_logic_vector(2337, 16),
14634 => conv_std_logic_vector(2394, 16),
14635 => conv_std_logic_vector(2451, 16),
14636 => conv_std_logic_vector(2508, 16),
14637 => conv_std_logic_vector(2565, 16),
14638 => conv_std_logic_vector(2622, 16),
14639 => conv_std_logic_vector(2679, 16),
14640 => conv_std_logic_vector(2736, 16),
14641 => conv_std_logic_vector(2793, 16),
14642 => conv_std_logic_vector(2850, 16),
14643 => conv_std_logic_vector(2907, 16),
14644 => conv_std_logic_vector(2964, 16),
14645 => conv_std_logic_vector(3021, 16),
14646 => conv_std_logic_vector(3078, 16),
14647 => conv_std_logic_vector(3135, 16),
14648 => conv_std_logic_vector(3192, 16),
14649 => conv_std_logic_vector(3249, 16),
14650 => conv_std_logic_vector(3306, 16),
14651 => conv_std_logic_vector(3363, 16),
14652 => conv_std_logic_vector(3420, 16),
14653 => conv_std_logic_vector(3477, 16),
14654 => conv_std_logic_vector(3534, 16),
14655 => conv_std_logic_vector(3591, 16),
14656 => conv_std_logic_vector(3648, 16),
14657 => conv_std_logic_vector(3705, 16),
14658 => conv_std_logic_vector(3762, 16),
14659 => conv_std_logic_vector(3819, 16),
14660 => conv_std_logic_vector(3876, 16),
14661 => conv_std_logic_vector(3933, 16),
14662 => conv_std_logic_vector(3990, 16),
14663 => conv_std_logic_vector(4047, 16),
14664 => conv_std_logic_vector(4104, 16),
14665 => conv_std_logic_vector(4161, 16),
14666 => conv_std_logic_vector(4218, 16),
14667 => conv_std_logic_vector(4275, 16),
14668 => conv_std_logic_vector(4332, 16),
14669 => conv_std_logic_vector(4389, 16),
14670 => conv_std_logic_vector(4446, 16),
14671 => conv_std_logic_vector(4503, 16),
14672 => conv_std_logic_vector(4560, 16),
14673 => conv_std_logic_vector(4617, 16),
14674 => conv_std_logic_vector(4674, 16),
14675 => conv_std_logic_vector(4731, 16),
14676 => conv_std_logic_vector(4788, 16),
14677 => conv_std_logic_vector(4845, 16),
14678 => conv_std_logic_vector(4902, 16),
14679 => conv_std_logic_vector(4959, 16),
14680 => conv_std_logic_vector(5016, 16),
14681 => conv_std_logic_vector(5073, 16),
14682 => conv_std_logic_vector(5130, 16),
14683 => conv_std_logic_vector(5187, 16),
14684 => conv_std_logic_vector(5244, 16),
14685 => conv_std_logic_vector(5301, 16),
14686 => conv_std_logic_vector(5358, 16),
14687 => conv_std_logic_vector(5415, 16),
14688 => conv_std_logic_vector(5472, 16),
14689 => conv_std_logic_vector(5529, 16),
14690 => conv_std_logic_vector(5586, 16),
14691 => conv_std_logic_vector(5643, 16),
14692 => conv_std_logic_vector(5700, 16),
14693 => conv_std_logic_vector(5757, 16),
14694 => conv_std_logic_vector(5814, 16),
14695 => conv_std_logic_vector(5871, 16),
14696 => conv_std_logic_vector(5928, 16),
14697 => conv_std_logic_vector(5985, 16),
14698 => conv_std_logic_vector(6042, 16),
14699 => conv_std_logic_vector(6099, 16),
14700 => conv_std_logic_vector(6156, 16),
14701 => conv_std_logic_vector(6213, 16),
14702 => conv_std_logic_vector(6270, 16),
14703 => conv_std_logic_vector(6327, 16),
14704 => conv_std_logic_vector(6384, 16),
14705 => conv_std_logic_vector(6441, 16),
14706 => conv_std_logic_vector(6498, 16),
14707 => conv_std_logic_vector(6555, 16),
14708 => conv_std_logic_vector(6612, 16),
14709 => conv_std_logic_vector(6669, 16),
14710 => conv_std_logic_vector(6726, 16),
14711 => conv_std_logic_vector(6783, 16),
14712 => conv_std_logic_vector(6840, 16),
14713 => conv_std_logic_vector(6897, 16),
14714 => conv_std_logic_vector(6954, 16),
14715 => conv_std_logic_vector(7011, 16),
14716 => conv_std_logic_vector(7068, 16),
14717 => conv_std_logic_vector(7125, 16),
14718 => conv_std_logic_vector(7182, 16),
14719 => conv_std_logic_vector(7239, 16),
14720 => conv_std_logic_vector(7296, 16),
14721 => conv_std_logic_vector(7353, 16),
14722 => conv_std_logic_vector(7410, 16),
14723 => conv_std_logic_vector(7467, 16),
14724 => conv_std_logic_vector(7524, 16),
14725 => conv_std_logic_vector(7581, 16),
14726 => conv_std_logic_vector(7638, 16),
14727 => conv_std_logic_vector(7695, 16),
14728 => conv_std_logic_vector(7752, 16),
14729 => conv_std_logic_vector(7809, 16),
14730 => conv_std_logic_vector(7866, 16),
14731 => conv_std_logic_vector(7923, 16),
14732 => conv_std_logic_vector(7980, 16),
14733 => conv_std_logic_vector(8037, 16),
14734 => conv_std_logic_vector(8094, 16),
14735 => conv_std_logic_vector(8151, 16),
14736 => conv_std_logic_vector(8208, 16),
14737 => conv_std_logic_vector(8265, 16),
14738 => conv_std_logic_vector(8322, 16),
14739 => conv_std_logic_vector(8379, 16),
14740 => conv_std_logic_vector(8436, 16),
14741 => conv_std_logic_vector(8493, 16),
14742 => conv_std_logic_vector(8550, 16),
14743 => conv_std_logic_vector(8607, 16),
14744 => conv_std_logic_vector(8664, 16),
14745 => conv_std_logic_vector(8721, 16),
14746 => conv_std_logic_vector(8778, 16),
14747 => conv_std_logic_vector(8835, 16),
14748 => conv_std_logic_vector(8892, 16),
14749 => conv_std_logic_vector(8949, 16),
14750 => conv_std_logic_vector(9006, 16),
14751 => conv_std_logic_vector(9063, 16),
14752 => conv_std_logic_vector(9120, 16),
14753 => conv_std_logic_vector(9177, 16),
14754 => conv_std_logic_vector(9234, 16),
14755 => conv_std_logic_vector(9291, 16),
14756 => conv_std_logic_vector(9348, 16),
14757 => conv_std_logic_vector(9405, 16),
14758 => conv_std_logic_vector(9462, 16),
14759 => conv_std_logic_vector(9519, 16),
14760 => conv_std_logic_vector(9576, 16),
14761 => conv_std_logic_vector(9633, 16),
14762 => conv_std_logic_vector(9690, 16),
14763 => conv_std_logic_vector(9747, 16),
14764 => conv_std_logic_vector(9804, 16),
14765 => conv_std_logic_vector(9861, 16),
14766 => conv_std_logic_vector(9918, 16),
14767 => conv_std_logic_vector(9975, 16),
14768 => conv_std_logic_vector(10032, 16),
14769 => conv_std_logic_vector(10089, 16),
14770 => conv_std_logic_vector(10146, 16),
14771 => conv_std_logic_vector(10203, 16),
14772 => conv_std_logic_vector(10260, 16),
14773 => conv_std_logic_vector(10317, 16),
14774 => conv_std_logic_vector(10374, 16),
14775 => conv_std_logic_vector(10431, 16),
14776 => conv_std_logic_vector(10488, 16),
14777 => conv_std_logic_vector(10545, 16),
14778 => conv_std_logic_vector(10602, 16),
14779 => conv_std_logic_vector(10659, 16),
14780 => conv_std_logic_vector(10716, 16),
14781 => conv_std_logic_vector(10773, 16),
14782 => conv_std_logic_vector(10830, 16),
14783 => conv_std_logic_vector(10887, 16),
14784 => conv_std_logic_vector(10944, 16),
14785 => conv_std_logic_vector(11001, 16),
14786 => conv_std_logic_vector(11058, 16),
14787 => conv_std_logic_vector(11115, 16),
14788 => conv_std_logic_vector(11172, 16),
14789 => conv_std_logic_vector(11229, 16),
14790 => conv_std_logic_vector(11286, 16),
14791 => conv_std_logic_vector(11343, 16),
14792 => conv_std_logic_vector(11400, 16),
14793 => conv_std_logic_vector(11457, 16),
14794 => conv_std_logic_vector(11514, 16),
14795 => conv_std_logic_vector(11571, 16),
14796 => conv_std_logic_vector(11628, 16),
14797 => conv_std_logic_vector(11685, 16),
14798 => conv_std_logic_vector(11742, 16),
14799 => conv_std_logic_vector(11799, 16),
14800 => conv_std_logic_vector(11856, 16),
14801 => conv_std_logic_vector(11913, 16),
14802 => conv_std_logic_vector(11970, 16),
14803 => conv_std_logic_vector(12027, 16),
14804 => conv_std_logic_vector(12084, 16),
14805 => conv_std_logic_vector(12141, 16),
14806 => conv_std_logic_vector(12198, 16),
14807 => conv_std_logic_vector(12255, 16),
14808 => conv_std_logic_vector(12312, 16),
14809 => conv_std_logic_vector(12369, 16),
14810 => conv_std_logic_vector(12426, 16),
14811 => conv_std_logic_vector(12483, 16),
14812 => conv_std_logic_vector(12540, 16),
14813 => conv_std_logic_vector(12597, 16),
14814 => conv_std_logic_vector(12654, 16),
14815 => conv_std_logic_vector(12711, 16),
14816 => conv_std_logic_vector(12768, 16),
14817 => conv_std_logic_vector(12825, 16),
14818 => conv_std_logic_vector(12882, 16),
14819 => conv_std_logic_vector(12939, 16),
14820 => conv_std_logic_vector(12996, 16),
14821 => conv_std_logic_vector(13053, 16),
14822 => conv_std_logic_vector(13110, 16),
14823 => conv_std_logic_vector(13167, 16),
14824 => conv_std_logic_vector(13224, 16),
14825 => conv_std_logic_vector(13281, 16),
14826 => conv_std_logic_vector(13338, 16),
14827 => conv_std_logic_vector(13395, 16),
14828 => conv_std_logic_vector(13452, 16),
14829 => conv_std_logic_vector(13509, 16),
14830 => conv_std_logic_vector(13566, 16),
14831 => conv_std_logic_vector(13623, 16),
14832 => conv_std_logic_vector(13680, 16),
14833 => conv_std_logic_vector(13737, 16),
14834 => conv_std_logic_vector(13794, 16),
14835 => conv_std_logic_vector(13851, 16),
14836 => conv_std_logic_vector(13908, 16),
14837 => conv_std_logic_vector(13965, 16),
14838 => conv_std_logic_vector(14022, 16),
14839 => conv_std_logic_vector(14079, 16),
14840 => conv_std_logic_vector(14136, 16),
14841 => conv_std_logic_vector(14193, 16),
14842 => conv_std_logic_vector(14250, 16),
14843 => conv_std_logic_vector(14307, 16),
14844 => conv_std_logic_vector(14364, 16),
14845 => conv_std_logic_vector(14421, 16),
14846 => conv_std_logic_vector(14478, 16),
14847 => conv_std_logic_vector(14535, 16),
14848 => conv_std_logic_vector(0, 16),
14849 => conv_std_logic_vector(58, 16),
14850 => conv_std_logic_vector(116, 16),
14851 => conv_std_logic_vector(174, 16),
14852 => conv_std_logic_vector(232, 16),
14853 => conv_std_logic_vector(290, 16),
14854 => conv_std_logic_vector(348, 16),
14855 => conv_std_logic_vector(406, 16),
14856 => conv_std_logic_vector(464, 16),
14857 => conv_std_logic_vector(522, 16),
14858 => conv_std_logic_vector(580, 16),
14859 => conv_std_logic_vector(638, 16),
14860 => conv_std_logic_vector(696, 16),
14861 => conv_std_logic_vector(754, 16),
14862 => conv_std_logic_vector(812, 16),
14863 => conv_std_logic_vector(870, 16),
14864 => conv_std_logic_vector(928, 16),
14865 => conv_std_logic_vector(986, 16),
14866 => conv_std_logic_vector(1044, 16),
14867 => conv_std_logic_vector(1102, 16),
14868 => conv_std_logic_vector(1160, 16),
14869 => conv_std_logic_vector(1218, 16),
14870 => conv_std_logic_vector(1276, 16),
14871 => conv_std_logic_vector(1334, 16),
14872 => conv_std_logic_vector(1392, 16),
14873 => conv_std_logic_vector(1450, 16),
14874 => conv_std_logic_vector(1508, 16),
14875 => conv_std_logic_vector(1566, 16),
14876 => conv_std_logic_vector(1624, 16),
14877 => conv_std_logic_vector(1682, 16),
14878 => conv_std_logic_vector(1740, 16),
14879 => conv_std_logic_vector(1798, 16),
14880 => conv_std_logic_vector(1856, 16),
14881 => conv_std_logic_vector(1914, 16),
14882 => conv_std_logic_vector(1972, 16),
14883 => conv_std_logic_vector(2030, 16),
14884 => conv_std_logic_vector(2088, 16),
14885 => conv_std_logic_vector(2146, 16),
14886 => conv_std_logic_vector(2204, 16),
14887 => conv_std_logic_vector(2262, 16),
14888 => conv_std_logic_vector(2320, 16),
14889 => conv_std_logic_vector(2378, 16),
14890 => conv_std_logic_vector(2436, 16),
14891 => conv_std_logic_vector(2494, 16),
14892 => conv_std_logic_vector(2552, 16),
14893 => conv_std_logic_vector(2610, 16),
14894 => conv_std_logic_vector(2668, 16),
14895 => conv_std_logic_vector(2726, 16),
14896 => conv_std_logic_vector(2784, 16),
14897 => conv_std_logic_vector(2842, 16),
14898 => conv_std_logic_vector(2900, 16),
14899 => conv_std_logic_vector(2958, 16),
14900 => conv_std_logic_vector(3016, 16),
14901 => conv_std_logic_vector(3074, 16),
14902 => conv_std_logic_vector(3132, 16),
14903 => conv_std_logic_vector(3190, 16),
14904 => conv_std_logic_vector(3248, 16),
14905 => conv_std_logic_vector(3306, 16),
14906 => conv_std_logic_vector(3364, 16),
14907 => conv_std_logic_vector(3422, 16),
14908 => conv_std_logic_vector(3480, 16),
14909 => conv_std_logic_vector(3538, 16),
14910 => conv_std_logic_vector(3596, 16),
14911 => conv_std_logic_vector(3654, 16),
14912 => conv_std_logic_vector(3712, 16),
14913 => conv_std_logic_vector(3770, 16),
14914 => conv_std_logic_vector(3828, 16),
14915 => conv_std_logic_vector(3886, 16),
14916 => conv_std_logic_vector(3944, 16),
14917 => conv_std_logic_vector(4002, 16),
14918 => conv_std_logic_vector(4060, 16),
14919 => conv_std_logic_vector(4118, 16),
14920 => conv_std_logic_vector(4176, 16),
14921 => conv_std_logic_vector(4234, 16),
14922 => conv_std_logic_vector(4292, 16),
14923 => conv_std_logic_vector(4350, 16),
14924 => conv_std_logic_vector(4408, 16),
14925 => conv_std_logic_vector(4466, 16),
14926 => conv_std_logic_vector(4524, 16),
14927 => conv_std_logic_vector(4582, 16),
14928 => conv_std_logic_vector(4640, 16),
14929 => conv_std_logic_vector(4698, 16),
14930 => conv_std_logic_vector(4756, 16),
14931 => conv_std_logic_vector(4814, 16),
14932 => conv_std_logic_vector(4872, 16),
14933 => conv_std_logic_vector(4930, 16),
14934 => conv_std_logic_vector(4988, 16),
14935 => conv_std_logic_vector(5046, 16),
14936 => conv_std_logic_vector(5104, 16),
14937 => conv_std_logic_vector(5162, 16),
14938 => conv_std_logic_vector(5220, 16),
14939 => conv_std_logic_vector(5278, 16),
14940 => conv_std_logic_vector(5336, 16),
14941 => conv_std_logic_vector(5394, 16),
14942 => conv_std_logic_vector(5452, 16),
14943 => conv_std_logic_vector(5510, 16),
14944 => conv_std_logic_vector(5568, 16),
14945 => conv_std_logic_vector(5626, 16),
14946 => conv_std_logic_vector(5684, 16),
14947 => conv_std_logic_vector(5742, 16),
14948 => conv_std_logic_vector(5800, 16),
14949 => conv_std_logic_vector(5858, 16),
14950 => conv_std_logic_vector(5916, 16),
14951 => conv_std_logic_vector(5974, 16),
14952 => conv_std_logic_vector(6032, 16),
14953 => conv_std_logic_vector(6090, 16),
14954 => conv_std_logic_vector(6148, 16),
14955 => conv_std_logic_vector(6206, 16),
14956 => conv_std_logic_vector(6264, 16),
14957 => conv_std_logic_vector(6322, 16),
14958 => conv_std_logic_vector(6380, 16),
14959 => conv_std_logic_vector(6438, 16),
14960 => conv_std_logic_vector(6496, 16),
14961 => conv_std_logic_vector(6554, 16),
14962 => conv_std_logic_vector(6612, 16),
14963 => conv_std_logic_vector(6670, 16),
14964 => conv_std_logic_vector(6728, 16),
14965 => conv_std_logic_vector(6786, 16),
14966 => conv_std_logic_vector(6844, 16),
14967 => conv_std_logic_vector(6902, 16),
14968 => conv_std_logic_vector(6960, 16),
14969 => conv_std_logic_vector(7018, 16),
14970 => conv_std_logic_vector(7076, 16),
14971 => conv_std_logic_vector(7134, 16),
14972 => conv_std_logic_vector(7192, 16),
14973 => conv_std_logic_vector(7250, 16),
14974 => conv_std_logic_vector(7308, 16),
14975 => conv_std_logic_vector(7366, 16),
14976 => conv_std_logic_vector(7424, 16),
14977 => conv_std_logic_vector(7482, 16),
14978 => conv_std_logic_vector(7540, 16),
14979 => conv_std_logic_vector(7598, 16),
14980 => conv_std_logic_vector(7656, 16),
14981 => conv_std_logic_vector(7714, 16),
14982 => conv_std_logic_vector(7772, 16),
14983 => conv_std_logic_vector(7830, 16),
14984 => conv_std_logic_vector(7888, 16),
14985 => conv_std_logic_vector(7946, 16),
14986 => conv_std_logic_vector(8004, 16),
14987 => conv_std_logic_vector(8062, 16),
14988 => conv_std_logic_vector(8120, 16),
14989 => conv_std_logic_vector(8178, 16),
14990 => conv_std_logic_vector(8236, 16),
14991 => conv_std_logic_vector(8294, 16),
14992 => conv_std_logic_vector(8352, 16),
14993 => conv_std_logic_vector(8410, 16),
14994 => conv_std_logic_vector(8468, 16),
14995 => conv_std_logic_vector(8526, 16),
14996 => conv_std_logic_vector(8584, 16),
14997 => conv_std_logic_vector(8642, 16),
14998 => conv_std_logic_vector(8700, 16),
14999 => conv_std_logic_vector(8758, 16),
15000 => conv_std_logic_vector(8816, 16),
15001 => conv_std_logic_vector(8874, 16),
15002 => conv_std_logic_vector(8932, 16),
15003 => conv_std_logic_vector(8990, 16),
15004 => conv_std_logic_vector(9048, 16),
15005 => conv_std_logic_vector(9106, 16),
15006 => conv_std_logic_vector(9164, 16),
15007 => conv_std_logic_vector(9222, 16),
15008 => conv_std_logic_vector(9280, 16),
15009 => conv_std_logic_vector(9338, 16),
15010 => conv_std_logic_vector(9396, 16),
15011 => conv_std_logic_vector(9454, 16),
15012 => conv_std_logic_vector(9512, 16),
15013 => conv_std_logic_vector(9570, 16),
15014 => conv_std_logic_vector(9628, 16),
15015 => conv_std_logic_vector(9686, 16),
15016 => conv_std_logic_vector(9744, 16),
15017 => conv_std_logic_vector(9802, 16),
15018 => conv_std_logic_vector(9860, 16),
15019 => conv_std_logic_vector(9918, 16),
15020 => conv_std_logic_vector(9976, 16),
15021 => conv_std_logic_vector(10034, 16),
15022 => conv_std_logic_vector(10092, 16),
15023 => conv_std_logic_vector(10150, 16),
15024 => conv_std_logic_vector(10208, 16),
15025 => conv_std_logic_vector(10266, 16),
15026 => conv_std_logic_vector(10324, 16),
15027 => conv_std_logic_vector(10382, 16),
15028 => conv_std_logic_vector(10440, 16),
15029 => conv_std_logic_vector(10498, 16),
15030 => conv_std_logic_vector(10556, 16),
15031 => conv_std_logic_vector(10614, 16),
15032 => conv_std_logic_vector(10672, 16),
15033 => conv_std_logic_vector(10730, 16),
15034 => conv_std_logic_vector(10788, 16),
15035 => conv_std_logic_vector(10846, 16),
15036 => conv_std_logic_vector(10904, 16),
15037 => conv_std_logic_vector(10962, 16),
15038 => conv_std_logic_vector(11020, 16),
15039 => conv_std_logic_vector(11078, 16),
15040 => conv_std_logic_vector(11136, 16),
15041 => conv_std_logic_vector(11194, 16),
15042 => conv_std_logic_vector(11252, 16),
15043 => conv_std_logic_vector(11310, 16),
15044 => conv_std_logic_vector(11368, 16),
15045 => conv_std_logic_vector(11426, 16),
15046 => conv_std_logic_vector(11484, 16),
15047 => conv_std_logic_vector(11542, 16),
15048 => conv_std_logic_vector(11600, 16),
15049 => conv_std_logic_vector(11658, 16),
15050 => conv_std_logic_vector(11716, 16),
15051 => conv_std_logic_vector(11774, 16),
15052 => conv_std_logic_vector(11832, 16),
15053 => conv_std_logic_vector(11890, 16),
15054 => conv_std_logic_vector(11948, 16),
15055 => conv_std_logic_vector(12006, 16),
15056 => conv_std_logic_vector(12064, 16),
15057 => conv_std_logic_vector(12122, 16),
15058 => conv_std_logic_vector(12180, 16),
15059 => conv_std_logic_vector(12238, 16),
15060 => conv_std_logic_vector(12296, 16),
15061 => conv_std_logic_vector(12354, 16),
15062 => conv_std_logic_vector(12412, 16),
15063 => conv_std_logic_vector(12470, 16),
15064 => conv_std_logic_vector(12528, 16),
15065 => conv_std_logic_vector(12586, 16),
15066 => conv_std_logic_vector(12644, 16),
15067 => conv_std_logic_vector(12702, 16),
15068 => conv_std_logic_vector(12760, 16),
15069 => conv_std_logic_vector(12818, 16),
15070 => conv_std_logic_vector(12876, 16),
15071 => conv_std_logic_vector(12934, 16),
15072 => conv_std_logic_vector(12992, 16),
15073 => conv_std_logic_vector(13050, 16),
15074 => conv_std_logic_vector(13108, 16),
15075 => conv_std_logic_vector(13166, 16),
15076 => conv_std_logic_vector(13224, 16),
15077 => conv_std_logic_vector(13282, 16),
15078 => conv_std_logic_vector(13340, 16),
15079 => conv_std_logic_vector(13398, 16),
15080 => conv_std_logic_vector(13456, 16),
15081 => conv_std_logic_vector(13514, 16),
15082 => conv_std_logic_vector(13572, 16),
15083 => conv_std_logic_vector(13630, 16),
15084 => conv_std_logic_vector(13688, 16),
15085 => conv_std_logic_vector(13746, 16),
15086 => conv_std_logic_vector(13804, 16),
15087 => conv_std_logic_vector(13862, 16),
15088 => conv_std_logic_vector(13920, 16),
15089 => conv_std_logic_vector(13978, 16),
15090 => conv_std_logic_vector(14036, 16),
15091 => conv_std_logic_vector(14094, 16),
15092 => conv_std_logic_vector(14152, 16),
15093 => conv_std_logic_vector(14210, 16),
15094 => conv_std_logic_vector(14268, 16),
15095 => conv_std_logic_vector(14326, 16),
15096 => conv_std_logic_vector(14384, 16),
15097 => conv_std_logic_vector(14442, 16),
15098 => conv_std_logic_vector(14500, 16),
15099 => conv_std_logic_vector(14558, 16),
15100 => conv_std_logic_vector(14616, 16),
15101 => conv_std_logic_vector(14674, 16),
15102 => conv_std_logic_vector(14732, 16),
15103 => conv_std_logic_vector(14790, 16),
15104 => conv_std_logic_vector(0, 16),
15105 => conv_std_logic_vector(59, 16),
15106 => conv_std_logic_vector(118, 16),
15107 => conv_std_logic_vector(177, 16),
15108 => conv_std_logic_vector(236, 16),
15109 => conv_std_logic_vector(295, 16),
15110 => conv_std_logic_vector(354, 16),
15111 => conv_std_logic_vector(413, 16),
15112 => conv_std_logic_vector(472, 16),
15113 => conv_std_logic_vector(531, 16),
15114 => conv_std_logic_vector(590, 16),
15115 => conv_std_logic_vector(649, 16),
15116 => conv_std_logic_vector(708, 16),
15117 => conv_std_logic_vector(767, 16),
15118 => conv_std_logic_vector(826, 16),
15119 => conv_std_logic_vector(885, 16),
15120 => conv_std_logic_vector(944, 16),
15121 => conv_std_logic_vector(1003, 16),
15122 => conv_std_logic_vector(1062, 16),
15123 => conv_std_logic_vector(1121, 16),
15124 => conv_std_logic_vector(1180, 16),
15125 => conv_std_logic_vector(1239, 16),
15126 => conv_std_logic_vector(1298, 16),
15127 => conv_std_logic_vector(1357, 16),
15128 => conv_std_logic_vector(1416, 16),
15129 => conv_std_logic_vector(1475, 16),
15130 => conv_std_logic_vector(1534, 16),
15131 => conv_std_logic_vector(1593, 16),
15132 => conv_std_logic_vector(1652, 16),
15133 => conv_std_logic_vector(1711, 16),
15134 => conv_std_logic_vector(1770, 16),
15135 => conv_std_logic_vector(1829, 16),
15136 => conv_std_logic_vector(1888, 16),
15137 => conv_std_logic_vector(1947, 16),
15138 => conv_std_logic_vector(2006, 16),
15139 => conv_std_logic_vector(2065, 16),
15140 => conv_std_logic_vector(2124, 16),
15141 => conv_std_logic_vector(2183, 16),
15142 => conv_std_logic_vector(2242, 16),
15143 => conv_std_logic_vector(2301, 16),
15144 => conv_std_logic_vector(2360, 16),
15145 => conv_std_logic_vector(2419, 16),
15146 => conv_std_logic_vector(2478, 16),
15147 => conv_std_logic_vector(2537, 16),
15148 => conv_std_logic_vector(2596, 16),
15149 => conv_std_logic_vector(2655, 16),
15150 => conv_std_logic_vector(2714, 16),
15151 => conv_std_logic_vector(2773, 16),
15152 => conv_std_logic_vector(2832, 16),
15153 => conv_std_logic_vector(2891, 16),
15154 => conv_std_logic_vector(2950, 16),
15155 => conv_std_logic_vector(3009, 16),
15156 => conv_std_logic_vector(3068, 16),
15157 => conv_std_logic_vector(3127, 16),
15158 => conv_std_logic_vector(3186, 16),
15159 => conv_std_logic_vector(3245, 16),
15160 => conv_std_logic_vector(3304, 16),
15161 => conv_std_logic_vector(3363, 16),
15162 => conv_std_logic_vector(3422, 16),
15163 => conv_std_logic_vector(3481, 16),
15164 => conv_std_logic_vector(3540, 16),
15165 => conv_std_logic_vector(3599, 16),
15166 => conv_std_logic_vector(3658, 16),
15167 => conv_std_logic_vector(3717, 16),
15168 => conv_std_logic_vector(3776, 16),
15169 => conv_std_logic_vector(3835, 16),
15170 => conv_std_logic_vector(3894, 16),
15171 => conv_std_logic_vector(3953, 16),
15172 => conv_std_logic_vector(4012, 16),
15173 => conv_std_logic_vector(4071, 16),
15174 => conv_std_logic_vector(4130, 16),
15175 => conv_std_logic_vector(4189, 16),
15176 => conv_std_logic_vector(4248, 16),
15177 => conv_std_logic_vector(4307, 16),
15178 => conv_std_logic_vector(4366, 16),
15179 => conv_std_logic_vector(4425, 16),
15180 => conv_std_logic_vector(4484, 16),
15181 => conv_std_logic_vector(4543, 16),
15182 => conv_std_logic_vector(4602, 16),
15183 => conv_std_logic_vector(4661, 16),
15184 => conv_std_logic_vector(4720, 16),
15185 => conv_std_logic_vector(4779, 16),
15186 => conv_std_logic_vector(4838, 16),
15187 => conv_std_logic_vector(4897, 16),
15188 => conv_std_logic_vector(4956, 16),
15189 => conv_std_logic_vector(5015, 16),
15190 => conv_std_logic_vector(5074, 16),
15191 => conv_std_logic_vector(5133, 16),
15192 => conv_std_logic_vector(5192, 16),
15193 => conv_std_logic_vector(5251, 16),
15194 => conv_std_logic_vector(5310, 16),
15195 => conv_std_logic_vector(5369, 16),
15196 => conv_std_logic_vector(5428, 16),
15197 => conv_std_logic_vector(5487, 16),
15198 => conv_std_logic_vector(5546, 16),
15199 => conv_std_logic_vector(5605, 16),
15200 => conv_std_logic_vector(5664, 16),
15201 => conv_std_logic_vector(5723, 16),
15202 => conv_std_logic_vector(5782, 16),
15203 => conv_std_logic_vector(5841, 16),
15204 => conv_std_logic_vector(5900, 16),
15205 => conv_std_logic_vector(5959, 16),
15206 => conv_std_logic_vector(6018, 16),
15207 => conv_std_logic_vector(6077, 16),
15208 => conv_std_logic_vector(6136, 16),
15209 => conv_std_logic_vector(6195, 16),
15210 => conv_std_logic_vector(6254, 16),
15211 => conv_std_logic_vector(6313, 16),
15212 => conv_std_logic_vector(6372, 16),
15213 => conv_std_logic_vector(6431, 16),
15214 => conv_std_logic_vector(6490, 16),
15215 => conv_std_logic_vector(6549, 16),
15216 => conv_std_logic_vector(6608, 16),
15217 => conv_std_logic_vector(6667, 16),
15218 => conv_std_logic_vector(6726, 16),
15219 => conv_std_logic_vector(6785, 16),
15220 => conv_std_logic_vector(6844, 16),
15221 => conv_std_logic_vector(6903, 16),
15222 => conv_std_logic_vector(6962, 16),
15223 => conv_std_logic_vector(7021, 16),
15224 => conv_std_logic_vector(7080, 16),
15225 => conv_std_logic_vector(7139, 16),
15226 => conv_std_logic_vector(7198, 16),
15227 => conv_std_logic_vector(7257, 16),
15228 => conv_std_logic_vector(7316, 16),
15229 => conv_std_logic_vector(7375, 16),
15230 => conv_std_logic_vector(7434, 16),
15231 => conv_std_logic_vector(7493, 16),
15232 => conv_std_logic_vector(7552, 16),
15233 => conv_std_logic_vector(7611, 16),
15234 => conv_std_logic_vector(7670, 16),
15235 => conv_std_logic_vector(7729, 16),
15236 => conv_std_logic_vector(7788, 16),
15237 => conv_std_logic_vector(7847, 16),
15238 => conv_std_logic_vector(7906, 16),
15239 => conv_std_logic_vector(7965, 16),
15240 => conv_std_logic_vector(8024, 16),
15241 => conv_std_logic_vector(8083, 16),
15242 => conv_std_logic_vector(8142, 16),
15243 => conv_std_logic_vector(8201, 16),
15244 => conv_std_logic_vector(8260, 16),
15245 => conv_std_logic_vector(8319, 16),
15246 => conv_std_logic_vector(8378, 16),
15247 => conv_std_logic_vector(8437, 16),
15248 => conv_std_logic_vector(8496, 16),
15249 => conv_std_logic_vector(8555, 16),
15250 => conv_std_logic_vector(8614, 16),
15251 => conv_std_logic_vector(8673, 16),
15252 => conv_std_logic_vector(8732, 16),
15253 => conv_std_logic_vector(8791, 16),
15254 => conv_std_logic_vector(8850, 16),
15255 => conv_std_logic_vector(8909, 16),
15256 => conv_std_logic_vector(8968, 16),
15257 => conv_std_logic_vector(9027, 16),
15258 => conv_std_logic_vector(9086, 16),
15259 => conv_std_logic_vector(9145, 16),
15260 => conv_std_logic_vector(9204, 16),
15261 => conv_std_logic_vector(9263, 16),
15262 => conv_std_logic_vector(9322, 16),
15263 => conv_std_logic_vector(9381, 16),
15264 => conv_std_logic_vector(9440, 16),
15265 => conv_std_logic_vector(9499, 16),
15266 => conv_std_logic_vector(9558, 16),
15267 => conv_std_logic_vector(9617, 16),
15268 => conv_std_logic_vector(9676, 16),
15269 => conv_std_logic_vector(9735, 16),
15270 => conv_std_logic_vector(9794, 16),
15271 => conv_std_logic_vector(9853, 16),
15272 => conv_std_logic_vector(9912, 16),
15273 => conv_std_logic_vector(9971, 16),
15274 => conv_std_logic_vector(10030, 16),
15275 => conv_std_logic_vector(10089, 16),
15276 => conv_std_logic_vector(10148, 16),
15277 => conv_std_logic_vector(10207, 16),
15278 => conv_std_logic_vector(10266, 16),
15279 => conv_std_logic_vector(10325, 16),
15280 => conv_std_logic_vector(10384, 16),
15281 => conv_std_logic_vector(10443, 16),
15282 => conv_std_logic_vector(10502, 16),
15283 => conv_std_logic_vector(10561, 16),
15284 => conv_std_logic_vector(10620, 16),
15285 => conv_std_logic_vector(10679, 16),
15286 => conv_std_logic_vector(10738, 16),
15287 => conv_std_logic_vector(10797, 16),
15288 => conv_std_logic_vector(10856, 16),
15289 => conv_std_logic_vector(10915, 16),
15290 => conv_std_logic_vector(10974, 16),
15291 => conv_std_logic_vector(11033, 16),
15292 => conv_std_logic_vector(11092, 16),
15293 => conv_std_logic_vector(11151, 16),
15294 => conv_std_logic_vector(11210, 16),
15295 => conv_std_logic_vector(11269, 16),
15296 => conv_std_logic_vector(11328, 16),
15297 => conv_std_logic_vector(11387, 16),
15298 => conv_std_logic_vector(11446, 16),
15299 => conv_std_logic_vector(11505, 16),
15300 => conv_std_logic_vector(11564, 16),
15301 => conv_std_logic_vector(11623, 16),
15302 => conv_std_logic_vector(11682, 16),
15303 => conv_std_logic_vector(11741, 16),
15304 => conv_std_logic_vector(11800, 16),
15305 => conv_std_logic_vector(11859, 16),
15306 => conv_std_logic_vector(11918, 16),
15307 => conv_std_logic_vector(11977, 16),
15308 => conv_std_logic_vector(12036, 16),
15309 => conv_std_logic_vector(12095, 16),
15310 => conv_std_logic_vector(12154, 16),
15311 => conv_std_logic_vector(12213, 16),
15312 => conv_std_logic_vector(12272, 16),
15313 => conv_std_logic_vector(12331, 16),
15314 => conv_std_logic_vector(12390, 16),
15315 => conv_std_logic_vector(12449, 16),
15316 => conv_std_logic_vector(12508, 16),
15317 => conv_std_logic_vector(12567, 16),
15318 => conv_std_logic_vector(12626, 16),
15319 => conv_std_logic_vector(12685, 16),
15320 => conv_std_logic_vector(12744, 16),
15321 => conv_std_logic_vector(12803, 16),
15322 => conv_std_logic_vector(12862, 16),
15323 => conv_std_logic_vector(12921, 16),
15324 => conv_std_logic_vector(12980, 16),
15325 => conv_std_logic_vector(13039, 16),
15326 => conv_std_logic_vector(13098, 16),
15327 => conv_std_logic_vector(13157, 16),
15328 => conv_std_logic_vector(13216, 16),
15329 => conv_std_logic_vector(13275, 16),
15330 => conv_std_logic_vector(13334, 16),
15331 => conv_std_logic_vector(13393, 16),
15332 => conv_std_logic_vector(13452, 16),
15333 => conv_std_logic_vector(13511, 16),
15334 => conv_std_logic_vector(13570, 16),
15335 => conv_std_logic_vector(13629, 16),
15336 => conv_std_logic_vector(13688, 16),
15337 => conv_std_logic_vector(13747, 16),
15338 => conv_std_logic_vector(13806, 16),
15339 => conv_std_logic_vector(13865, 16),
15340 => conv_std_logic_vector(13924, 16),
15341 => conv_std_logic_vector(13983, 16),
15342 => conv_std_logic_vector(14042, 16),
15343 => conv_std_logic_vector(14101, 16),
15344 => conv_std_logic_vector(14160, 16),
15345 => conv_std_logic_vector(14219, 16),
15346 => conv_std_logic_vector(14278, 16),
15347 => conv_std_logic_vector(14337, 16),
15348 => conv_std_logic_vector(14396, 16),
15349 => conv_std_logic_vector(14455, 16),
15350 => conv_std_logic_vector(14514, 16),
15351 => conv_std_logic_vector(14573, 16),
15352 => conv_std_logic_vector(14632, 16),
15353 => conv_std_logic_vector(14691, 16),
15354 => conv_std_logic_vector(14750, 16),
15355 => conv_std_logic_vector(14809, 16),
15356 => conv_std_logic_vector(14868, 16),
15357 => conv_std_logic_vector(14927, 16),
15358 => conv_std_logic_vector(14986, 16),
15359 => conv_std_logic_vector(15045, 16),
15360 => conv_std_logic_vector(0, 16),
15361 => conv_std_logic_vector(60, 16),
15362 => conv_std_logic_vector(120, 16),
15363 => conv_std_logic_vector(180, 16),
15364 => conv_std_logic_vector(240, 16),
15365 => conv_std_logic_vector(300, 16),
15366 => conv_std_logic_vector(360, 16),
15367 => conv_std_logic_vector(420, 16),
15368 => conv_std_logic_vector(480, 16),
15369 => conv_std_logic_vector(540, 16),
15370 => conv_std_logic_vector(600, 16),
15371 => conv_std_logic_vector(660, 16),
15372 => conv_std_logic_vector(720, 16),
15373 => conv_std_logic_vector(780, 16),
15374 => conv_std_logic_vector(840, 16),
15375 => conv_std_logic_vector(900, 16),
15376 => conv_std_logic_vector(960, 16),
15377 => conv_std_logic_vector(1020, 16),
15378 => conv_std_logic_vector(1080, 16),
15379 => conv_std_logic_vector(1140, 16),
15380 => conv_std_logic_vector(1200, 16),
15381 => conv_std_logic_vector(1260, 16),
15382 => conv_std_logic_vector(1320, 16),
15383 => conv_std_logic_vector(1380, 16),
15384 => conv_std_logic_vector(1440, 16),
15385 => conv_std_logic_vector(1500, 16),
15386 => conv_std_logic_vector(1560, 16),
15387 => conv_std_logic_vector(1620, 16),
15388 => conv_std_logic_vector(1680, 16),
15389 => conv_std_logic_vector(1740, 16),
15390 => conv_std_logic_vector(1800, 16),
15391 => conv_std_logic_vector(1860, 16),
15392 => conv_std_logic_vector(1920, 16),
15393 => conv_std_logic_vector(1980, 16),
15394 => conv_std_logic_vector(2040, 16),
15395 => conv_std_logic_vector(2100, 16),
15396 => conv_std_logic_vector(2160, 16),
15397 => conv_std_logic_vector(2220, 16),
15398 => conv_std_logic_vector(2280, 16),
15399 => conv_std_logic_vector(2340, 16),
15400 => conv_std_logic_vector(2400, 16),
15401 => conv_std_logic_vector(2460, 16),
15402 => conv_std_logic_vector(2520, 16),
15403 => conv_std_logic_vector(2580, 16),
15404 => conv_std_logic_vector(2640, 16),
15405 => conv_std_logic_vector(2700, 16),
15406 => conv_std_logic_vector(2760, 16),
15407 => conv_std_logic_vector(2820, 16),
15408 => conv_std_logic_vector(2880, 16),
15409 => conv_std_logic_vector(2940, 16),
15410 => conv_std_logic_vector(3000, 16),
15411 => conv_std_logic_vector(3060, 16),
15412 => conv_std_logic_vector(3120, 16),
15413 => conv_std_logic_vector(3180, 16),
15414 => conv_std_logic_vector(3240, 16),
15415 => conv_std_logic_vector(3300, 16),
15416 => conv_std_logic_vector(3360, 16),
15417 => conv_std_logic_vector(3420, 16),
15418 => conv_std_logic_vector(3480, 16),
15419 => conv_std_logic_vector(3540, 16),
15420 => conv_std_logic_vector(3600, 16),
15421 => conv_std_logic_vector(3660, 16),
15422 => conv_std_logic_vector(3720, 16),
15423 => conv_std_logic_vector(3780, 16),
15424 => conv_std_logic_vector(3840, 16),
15425 => conv_std_logic_vector(3900, 16),
15426 => conv_std_logic_vector(3960, 16),
15427 => conv_std_logic_vector(4020, 16),
15428 => conv_std_logic_vector(4080, 16),
15429 => conv_std_logic_vector(4140, 16),
15430 => conv_std_logic_vector(4200, 16),
15431 => conv_std_logic_vector(4260, 16),
15432 => conv_std_logic_vector(4320, 16),
15433 => conv_std_logic_vector(4380, 16),
15434 => conv_std_logic_vector(4440, 16),
15435 => conv_std_logic_vector(4500, 16),
15436 => conv_std_logic_vector(4560, 16),
15437 => conv_std_logic_vector(4620, 16),
15438 => conv_std_logic_vector(4680, 16),
15439 => conv_std_logic_vector(4740, 16),
15440 => conv_std_logic_vector(4800, 16),
15441 => conv_std_logic_vector(4860, 16),
15442 => conv_std_logic_vector(4920, 16),
15443 => conv_std_logic_vector(4980, 16),
15444 => conv_std_logic_vector(5040, 16),
15445 => conv_std_logic_vector(5100, 16),
15446 => conv_std_logic_vector(5160, 16),
15447 => conv_std_logic_vector(5220, 16),
15448 => conv_std_logic_vector(5280, 16),
15449 => conv_std_logic_vector(5340, 16),
15450 => conv_std_logic_vector(5400, 16),
15451 => conv_std_logic_vector(5460, 16),
15452 => conv_std_logic_vector(5520, 16),
15453 => conv_std_logic_vector(5580, 16),
15454 => conv_std_logic_vector(5640, 16),
15455 => conv_std_logic_vector(5700, 16),
15456 => conv_std_logic_vector(5760, 16),
15457 => conv_std_logic_vector(5820, 16),
15458 => conv_std_logic_vector(5880, 16),
15459 => conv_std_logic_vector(5940, 16),
15460 => conv_std_logic_vector(6000, 16),
15461 => conv_std_logic_vector(6060, 16),
15462 => conv_std_logic_vector(6120, 16),
15463 => conv_std_logic_vector(6180, 16),
15464 => conv_std_logic_vector(6240, 16),
15465 => conv_std_logic_vector(6300, 16),
15466 => conv_std_logic_vector(6360, 16),
15467 => conv_std_logic_vector(6420, 16),
15468 => conv_std_logic_vector(6480, 16),
15469 => conv_std_logic_vector(6540, 16),
15470 => conv_std_logic_vector(6600, 16),
15471 => conv_std_logic_vector(6660, 16),
15472 => conv_std_logic_vector(6720, 16),
15473 => conv_std_logic_vector(6780, 16),
15474 => conv_std_logic_vector(6840, 16),
15475 => conv_std_logic_vector(6900, 16),
15476 => conv_std_logic_vector(6960, 16),
15477 => conv_std_logic_vector(7020, 16),
15478 => conv_std_logic_vector(7080, 16),
15479 => conv_std_logic_vector(7140, 16),
15480 => conv_std_logic_vector(7200, 16),
15481 => conv_std_logic_vector(7260, 16),
15482 => conv_std_logic_vector(7320, 16),
15483 => conv_std_logic_vector(7380, 16),
15484 => conv_std_logic_vector(7440, 16),
15485 => conv_std_logic_vector(7500, 16),
15486 => conv_std_logic_vector(7560, 16),
15487 => conv_std_logic_vector(7620, 16),
15488 => conv_std_logic_vector(7680, 16),
15489 => conv_std_logic_vector(7740, 16),
15490 => conv_std_logic_vector(7800, 16),
15491 => conv_std_logic_vector(7860, 16),
15492 => conv_std_logic_vector(7920, 16),
15493 => conv_std_logic_vector(7980, 16),
15494 => conv_std_logic_vector(8040, 16),
15495 => conv_std_logic_vector(8100, 16),
15496 => conv_std_logic_vector(8160, 16),
15497 => conv_std_logic_vector(8220, 16),
15498 => conv_std_logic_vector(8280, 16),
15499 => conv_std_logic_vector(8340, 16),
15500 => conv_std_logic_vector(8400, 16),
15501 => conv_std_logic_vector(8460, 16),
15502 => conv_std_logic_vector(8520, 16),
15503 => conv_std_logic_vector(8580, 16),
15504 => conv_std_logic_vector(8640, 16),
15505 => conv_std_logic_vector(8700, 16),
15506 => conv_std_logic_vector(8760, 16),
15507 => conv_std_logic_vector(8820, 16),
15508 => conv_std_logic_vector(8880, 16),
15509 => conv_std_logic_vector(8940, 16),
15510 => conv_std_logic_vector(9000, 16),
15511 => conv_std_logic_vector(9060, 16),
15512 => conv_std_logic_vector(9120, 16),
15513 => conv_std_logic_vector(9180, 16),
15514 => conv_std_logic_vector(9240, 16),
15515 => conv_std_logic_vector(9300, 16),
15516 => conv_std_logic_vector(9360, 16),
15517 => conv_std_logic_vector(9420, 16),
15518 => conv_std_logic_vector(9480, 16),
15519 => conv_std_logic_vector(9540, 16),
15520 => conv_std_logic_vector(9600, 16),
15521 => conv_std_logic_vector(9660, 16),
15522 => conv_std_logic_vector(9720, 16),
15523 => conv_std_logic_vector(9780, 16),
15524 => conv_std_logic_vector(9840, 16),
15525 => conv_std_logic_vector(9900, 16),
15526 => conv_std_logic_vector(9960, 16),
15527 => conv_std_logic_vector(10020, 16),
15528 => conv_std_logic_vector(10080, 16),
15529 => conv_std_logic_vector(10140, 16),
15530 => conv_std_logic_vector(10200, 16),
15531 => conv_std_logic_vector(10260, 16),
15532 => conv_std_logic_vector(10320, 16),
15533 => conv_std_logic_vector(10380, 16),
15534 => conv_std_logic_vector(10440, 16),
15535 => conv_std_logic_vector(10500, 16),
15536 => conv_std_logic_vector(10560, 16),
15537 => conv_std_logic_vector(10620, 16),
15538 => conv_std_logic_vector(10680, 16),
15539 => conv_std_logic_vector(10740, 16),
15540 => conv_std_logic_vector(10800, 16),
15541 => conv_std_logic_vector(10860, 16),
15542 => conv_std_logic_vector(10920, 16),
15543 => conv_std_logic_vector(10980, 16),
15544 => conv_std_logic_vector(11040, 16),
15545 => conv_std_logic_vector(11100, 16),
15546 => conv_std_logic_vector(11160, 16),
15547 => conv_std_logic_vector(11220, 16),
15548 => conv_std_logic_vector(11280, 16),
15549 => conv_std_logic_vector(11340, 16),
15550 => conv_std_logic_vector(11400, 16),
15551 => conv_std_logic_vector(11460, 16),
15552 => conv_std_logic_vector(11520, 16),
15553 => conv_std_logic_vector(11580, 16),
15554 => conv_std_logic_vector(11640, 16),
15555 => conv_std_logic_vector(11700, 16),
15556 => conv_std_logic_vector(11760, 16),
15557 => conv_std_logic_vector(11820, 16),
15558 => conv_std_logic_vector(11880, 16),
15559 => conv_std_logic_vector(11940, 16),
15560 => conv_std_logic_vector(12000, 16),
15561 => conv_std_logic_vector(12060, 16),
15562 => conv_std_logic_vector(12120, 16),
15563 => conv_std_logic_vector(12180, 16),
15564 => conv_std_logic_vector(12240, 16),
15565 => conv_std_logic_vector(12300, 16),
15566 => conv_std_logic_vector(12360, 16),
15567 => conv_std_logic_vector(12420, 16),
15568 => conv_std_logic_vector(12480, 16),
15569 => conv_std_logic_vector(12540, 16),
15570 => conv_std_logic_vector(12600, 16),
15571 => conv_std_logic_vector(12660, 16),
15572 => conv_std_logic_vector(12720, 16),
15573 => conv_std_logic_vector(12780, 16),
15574 => conv_std_logic_vector(12840, 16),
15575 => conv_std_logic_vector(12900, 16),
15576 => conv_std_logic_vector(12960, 16),
15577 => conv_std_logic_vector(13020, 16),
15578 => conv_std_logic_vector(13080, 16),
15579 => conv_std_logic_vector(13140, 16),
15580 => conv_std_logic_vector(13200, 16),
15581 => conv_std_logic_vector(13260, 16),
15582 => conv_std_logic_vector(13320, 16),
15583 => conv_std_logic_vector(13380, 16),
15584 => conv_std_logic_vector(13440, 16),
15585 => conv_std_logic_vector(13500, 16),
15586 => conv_std_logic_vector(13560, 16),
15587 => conv_std_logic_vector(13620, 16),
15588 => conv_std_logic_vector(13680, 16),
15589 => conv_std_logic_vector(13740, 16),
15590 => conv_std_logic_vector(13800, 16),
15591 => conv_std_logic_vector(13860, 16),
15592 => conv_std_logic_vector(13920, 16),
15593 => conv_std_logic_vector(13980, 16),
15594 => conv_std_logic_vector(14040, 16),
15595 => conv_std_logic_vector(14100, 16),
15596 => conv_std_logic_vector(14160, 16),
15597 => conv_std_logic_vector(14220, 16),
15598 => conv_std_logic_vector(14280, 16),
15599 => conv_std_logic_vector(14340, 16),
15600 => conv_std_logic_vector(14400, 16),
15601 => conv_std_logic_vector(14460, 16),
15602 => conv_std_logic_vector(14520, 16),
15603 => conv_std_logic_vector(14580, 16),
15604 => conv_std_logic_vector(14640, 16),
15605 => conv_std_logic_vector(14700, 16),
15606 => conv_std_logic_vector(14760, 16),
15607 => conv_std_logic_vector(14820, 16),
15608 => conv_std_logic_vector(14880, 16),
15609 => conv_std_logic_vector(14940, 16),
15610 => conv_std_logic_vector(15000, 16),
15611 => conv_std_logic_vector(15060, 16),
15612 => conv_std_logic_vector(15120, 16),
15613 => conv_std_logic_vector(15180, 16),
15614 => conv_std_logic_vector(15240, 16),
15615 => conv_std_logic_vector(15300, 16),
15616 => conv_std_logic_vector(0, 16),
15617 => conv_std_logic_vector(61, 16),
15618 => conv_std_logic_vector(122, 16),
15619 => conv_std_logic_vector(183, 16),
15620 => conv_std_logic_vector(244, 16),
15621 => conv_std_logic_vector(305, 16),
15622 => conv_std_logic_vector(366, 16),
15623 => conv_std_logic_vector(427, 16),
15624 => conv_std_logic_vector(488, 16),
15625 => conv_std_logic_vector(549, 16),
15626 => conv_std_logic_vector(610, 16),
15627 => conv_std_logic_vector(671, 16),
15628 => conv_std_logic_vector(732, 16),
15629 => conv_std_logic_vector(793, 16),
15630 => conv_std_logic_vector(854, 16),
15631 => conv_std_logic_vector(915, 16),
15632 => conv_std_logic_vector(976, 16),
15633 => conv_std_logic_vector(1037, 16),
15634 => conv_std_logic_vector(1098, 16),
15635 => conv_std_logic_vector(1159, 16),
15636 => conv_std_logic_vector(1220, 16),
15637 => conv_std_logic_vector(1281, 16),
15638 => conv_std_logic_vector(1342, 16),
15639 => conv_std_logic_vector(1403, 16),
15640 => conv_std_logic_vector(1464, 16),
15641 => conv_std_logic_vector(1525, 16),
15642 => conv_std_logic_vector(1586, 16),
15643 => conv_std_logic_vector(1647, 16),
15644 => conv_std_logic_vector(1708, 16),
15645 => conv_std_logic_vector(1769, 16),
15646 => conv_std_logic_vector(1830, 16),
15647 => conv_std_logic_vector(1891, 16),
15648 => conv_std_logic_vector(1952, 16),
15649 => conv_std_logic_vector(2013, 16),
15650 => conv_std_logic_vector(2074, 16),
15651 => conv_std_logic_vector(2135, 16),
15652 => conv_std_logic_vector(2196, 16),
15653 => conv_std_logic_vector(2257, 16),
15654 => conv_std_logic_vector(2318, 16),
15655 => conv_std_logic_vector(2379, 16),
15656 => conv_std_logic_vector(2440, 16),
15657 => conv_std_logic_vector(2501, 16),
15658 => conv_std_logic_vector(2562, 16),
15659 => conv_std_logic_vector(2623, 16),
15660 => conv_std_logic_vector(2684, 16),
15661 => conv_std_logic_vector(2745, 16),
15662 => conv_std_logic_vector(2806, 16),
15663 => conv_std_logic_vector(2867, 16),
15664 => conv_std_logic_vector(2928, 16),
15665 => conv_std_logic_vector(2989, 16),
15666 => conv_std_logic_vector(3050, 16),
15667 => conv_std_logic_vector(3111, 16),
15668 => conv_std_logic_vector(3172, 16),
15669 => conv_std_logic_vector(3233, 16),
15670 => conv_std_logic_vector(3294, 16),
15671 => conv_std_logic_vector(3355, 16),
15672 => conv_std_logic_vector(3416, 16),
15673 => conv_std_logic_vector(3477, 16),
15674 => conv_std_logic_vector(3538, 16),
15675 => conv_std_logic_vector(3599, 16),
15676 => conv_std_logic_vector(3660, 16),
15677 => conv_std_logic_vector(3721, 16),
15678 => conv_std_logic_vector(3782, 16),
15679 => conv_std_logic_vector(3843, 16),
15680 => conv_std_logic_vector(3904, 16),
15681 => conv_std_logic_vector(3965, 16),
15682 => conv_std_logic_vector(4026, 16),
15683 => conv_std_logic_vector(4087, 16),
15684 => conv_std_logic_vector(4148, 16),
15685 => conv_std_logic_vector(4209, 16),
15686 => conv_std_logic_vector(4270, 16),
15687 => conv_std_logic_vector(4331, 16),
15688 => conv_std_logic_vector(4392, 16),
15689 => conv_std_logic_vector(4453, 16),
15690 => conv_std_logic_vector(4514, 16),
15691 => conv_std_logic_vector(4575, 16),
15692 => conv_std_logic_vector(4636, 16),
15693 => conv_std_logic_vector(4697, 16),
15694 => conv_std_logic_vector(4758, 16),
15695 => conv_std_logic_vector(4819, 16),
15696 => conv_std_logic_vector(4880, 16),
15697 => conv_std_logic_vector(4941, 16),
15698 => conv_std_logic_vector(5002, 16),
15699 => conv_std_logic_vector(5063, 16),
15700 => conv_std_logic_vector(5124, 16),
15701 => conv_std_logic_vector(5185, 16),
15702 => conv_std_logic_vector(5246, 16),
15703 => conv_std_logic_vector(5307, 16),
15704 => conv_std_logic_vector(5368, 16),
15705 => conv_std_logic_vector(5429, 16),
15706 => conv_std_logic_vector(5490, 16),
15707 => conv_std_logic_vector(5551, 16),
15708 => conv_std_logic_vector(5612, 16),
15709 => conv_std_logic_vector(5673, 16),
15710 => conv_std_logic_vector(5734, 16),
15711 => conv_std_logic_vector(5795, 16),
15712 => conv_std_logic_vector(5856, 16),
15713 => conv_std_logic_vector(5917, 16),
15714 => conv_std_logic_vector(5978, 16),
15715 => conv_std_logic_vector(6039, 16),
15716 => conv_std_logic_vector(6100, 16),
15717 => conv_std_logic_vector(6161, 16),
15718 => conv_std_logic_vector(6222, 16),
15719 => conv_std_logic_vector(6283, 16),
15720 => conv_std_logic_vector(6344, 16),
15721 => conv_std_logic_vector(6405, 16),
15722 => conv_std_logic_vector(6466, 16),
15723 => conv_std_logic_vector(6527, 16),
15724 => conv_std_logic_vector(6588, 16),
15725 => conv_std_logic_vector(6649, 16),
15726 => conv_std_logic_vector(6710, 16),
15727 => conv_std_logic_vector(6771, 16),
15728 => conv_std_logic_vector(6832, 16),
15729 => conv_std_logic_vector(6893, 16),
15730 => conv_std_logic_vector(6954, 16),
15731 => conv_std_logic_vector(7015, 16),
15732 => conv_std_logic_vector(7076, 16),
15733 => conv_std_logic_vector(7137, 16),
15734 => conv_std_logic_vector(7198, 16),
15735 => conv_std_logic_vector(7259, 16),
15736 => conv_std_logic_vector(7320, 16),
15737 => conv_std_logic_vector(7381, 16),
15738 => conv_std_logic_vector(7442, 16),
15739 => conv_std_logic_vector(7503, 16),
15740 => conv_std_logic_vector(7564, 16),
15741 => conv_std_logic_vector(7625, 16),
15742 => conv_std_logic_vector(7686, 16),
15743 => conv_std_logic_vector(7747, 16),
15744 => conv_std_logic_vector(7808, 16),
15745 => conv_std_logic_vector(7869, 16),
15746 => conv_std_logic_vector(7930, 16),
15747 => conv_std_logic_vector(7991, 16),
15748 => conv_std_logic_vector(8052, 16),
15749 => conv_std_logic_vector(8113, 16),
15750 => conv_std_logic_vector(8174, 16),
15751 => conv_std_logic_vector(8235, 16),
15752 => conv_std_logic_vector(8296, 16),
15753 => conv_std_logic_vector(8357, 16),
15754 => conv_std_logic_vector(8418, 16),
15755 => conv_std_logic_vector(8479, 16),
15756 => conv_std_logic_vector(8540, 16),
15757 => conv_std_logic_vector(8601, 16),
15758 => conv_std_logic_vector(8662, 16),
15759 => conv_std_logic_vector(8723, 16),
15760 => conv_std_logic_vector(8784, 16),
15761 => conv_std_logic_vector(8845, 16),
15762 => conv_std_logic_vector(8906, 16),
15763 => conv_std_logic_vector(8967, 16),
15764 => conv_std_logic_vector(9028, 16),
15765 => conv_std_logic_vector(9089, 16),
15766 => conv_std_logic_vector(9150, 16),
15767 => conv_std_logic_vector(9211, 16),
15768 => conv_std_logic_vector(9272, 16),
15769 => conv_std_logic_vector(9333, 16),
15770 => conv_std_logic_vector(9394, 16),
15771 => conv_std_logic_vector(9455, 16),
15772 => conv_std_logic_vector(9516, 16),
15773 => conv_std_logic_vector(9577, 16),
15774 => conv_std_logic_vector(9638, 16),
15775 => conv_std_logic_vector(9699, 16),
15776 => conv_std_logic_vector(9760, 16),
15777 => conv_std_logic_vector(9821, 16),
15778 => conv_std_logic_vector(9882, 16),
15779 => conv_std_logic_vector(9943, 16),
15780 => conv_std_logic_vector(10004, 16),
15781 => conv_std_logic_vector(10065, 16),
15782 => conv_std_logic_vector(10126, 16),
15783 => conv_std_logic_vector(10187, 16),
15784 => conv_std_logic_vector(10248, 16),
15785 => conv_std_logic_vector(10309, 16),
15786 => conv_std_logic_vector(10370, 16),
15787 => conv_std_logic_vector(10431, 16),
15788 => conv_std_logic_vector(10492, 16),
15789 => conv_std_logic_vector(10553, 16),
15790 => conv_std_logic_vector(10614, 16),
15791 => conv_std_logic_vector(10675, 16),
15792 => conv_std_logic_vector(10736, 16),
15793 => conv_std_logic_vector(10797, 16),
15794 => conv_std_logic_vector(10858, 16),
15795 => conv_std_logic_vector(10919, 16),
15796 => conv_std_logic_vector(10980, 16),
15797 => conv_std_logic_vector(11041, 16),
15798 => conv_std_logic_vector(11102, 16),
15799 => conv_std_logic_vector(11163, 16),
15800 => conv_std_logic_vector(11224, 16),
15801 => conv_std_logic_vector(11285, 16),
15802 => conv_std_logic_vector(11346, 16),
15803 => conv_std_logic_vector(11407, 16),
15804 => conv_std_logic_vector(11468, 16),
15805 => conv_std_logic_vector(11529, 16),
15806 => conv_std_logic_vector(11590, 16),
15807 => conv_std_logic_vector(11651, 16),
15808 => conv_std_logic_vector(11712, 16),
15809 => conv_std_logic_vector(11773, 16),
15810 => conv_std_logic_vector(11834, 16),
15811 => conv_std_logic_vector(11895, 16),
15812 => conv_std_logic_vector(11956, 16),
15813 => conv_std_logic_vector(12017, 16),
15814 => conv_std_logic_vector(12078, 16),
15815 => conv_std_logic_vector(12139, 16),
15816 => conv_std_logic_vector(12200, 16),
15817 => conv_std_logic_vector(12261, 16),
15818 => conv_std_logic_vector(12322, 16),
15819 => conv_std_logic_vector(12383, 16),
15820 => conv_std_logic_vector(12444, 16),
15821 => conv_std_logic_vector(12505, 16),
15822 => conv_std_logic_vector(12566, 16),
15823 => conv_std_logic_vector(12627, 16),
15824 => conv_std_logic_vector(12688, 16),
15825 => conv_std_logic_vector(12749, 16),
15826 => conv_std_logic_vector(12810, 16),
15827 => conv_std_logic_vector(12871, 16),
15828 => conv_std_logic_vector(12932, 16),
15829 => conv_std_logic_vector(12993, 16),
15830 => conv_std_logic_vector(13054, 16),
15831 => conv_std_logic_vector(13115, 16),
15832 => conv_std_logic_vector(13176, 16),
15833 => conv_std_logic_vector(13237, 16),
15834 => conv_std_logic_vector(13298, 16),
15835 => conv_std_logic_vector(13359, 16),
15836 => conv_std_logic_vector(13420, 16),
15837 => conv_std_logic_vector(13481, 16),
15838 => conv_std_logic_vector(13542, 16),
15839 => conv_std_logic_vector(13603, 16),
15840 => conv_std_logic_vector(13664, 16),
15841 => conv_std_logic_vector(13725, 16),
15842 => conv_std_logic_vector(13786, 16),
15843 => conv_std_logic_vector(13847, 16),
15844 => conv_std_logic_vector(13908, 16),
15845 => conv_std_logic_vector(13969, 16),
15846 => conv_std_logic_vector(14030, 16),
15847 => conv_std_logic_vector(14091, 16),
15848 => conv_std_logic_vector(14152, 16),
15849 => conv_std_logic_vector(14213, 16),
15850 => conv_std_logic_vector(14274, 16),
15851 => conv_std_logic_vector(14335, 16),
15852 => conv_std_logic_vector(14396, 16),
15853 => conv_std_logic_vector(14457, 16),
15854 => conv_std_logic_vector(14518, 16),
15855 => conv_std_logic_vector(14579, 16),
15856 => conv_std_logic_vector(14640, 16),
15857 => conv_std_logic_vector(14701, 16),
15858 => conv_std_logic_vector(14762, 16),
15859 => conv_std_logic_vector(14823, 16),
15860 => conv_std_logic_vector(14884, 16),
15861 => conv_std_logic_vector(14945, 16),
15862 => conv_std_logic_vector(15006, 16),
15863 => conv_std_logic_vector(15067, 16),
15864 => conv_std_logic_vector(15128, 16),
15865 => conv_std_logic_vector(15189, 16),
15866 => conv_std_logic_vector(15250, 16),
15867 => conv_std_logic_vector(15311, 16),
15868 => conv_std_logic_vector(15372, 16),
15869 => conv_std_logic_vector(15433, 16),
15870 => conv_std_logic_vector(15494, 16),
15871 => conv_std_logic_vector(15555, 16),
15872 => conv_std_logic_vector(0, 16),
15873 => conv_std_logic_vector(62, 16),
15874 => conv_std_logic_vector(124, 16),
15875 => conv_std_logic_vector(186, 16),
15876 => conv_std_logic_vector(248, 16),
15877 => conv_std_logic_vector(310, 16),
15878 => conv_std_logic_vector(372, 16),
15879 => conv_std_logic_vector(434, 16),
15880 => conv_std_logic_vector(496, 16),
15881 => conv_std_logic_vector(558, 16),
15882 => conv_std_logic_vector(620, 16),
15883 => conv_std_logic_vector(682, 16),
15884 => conv_std_logic_vector(744, 16),
15885 => conv_std_logic_vector(806, 16),
15886 => conv_std_logic_vector(868, 16),
15887 => conv_std_logic_vector(930, 16),
15888 => conv_std_logic_vector(992, 16),
15889 => conv_std_logic_vector(1054, 16),
15890 => conv_std_logic_vector(1116, 16),
15891 => conv_std_logic_vector(1178, 16),
15892 => conv_std_logic_vector(1240, 16),
15893 => conv_std_logic_vector(1302, 16),
15894 => conv_std_logic_vector(1364, 16),
15895 => conv_std_logic_vector(1426, 16),
15896 => conv_std_logic_vector(1488, 16),
15897 => conv_std_logic_vector(1550, 16),
15898 => conv_std_logic_vector(1612, 16),
15899 => conv_std_logic_vector(1674, 16),
15900 => conv_std_logic_vector(1736, 16),
15901 => conv_std_logic_vector(1798, 16),
15902 => conv_std_logic_vector(1860, 16),
15903 => conv_std_logic_vector(1922, 16),
15904 => conv_std_logic_vector(1984, 16),
15905 => conv_std_logic_vector(2046, 16),
15906 => conv_std_logic_vector(2108, 16),
15907 => conv_std_logic_vector(2170, 16),
15908 => conv_std_logic_vector(2232, 16),
15909 => conv_std_logic_vector(2294, 16),
15910 => conv_std_logic_vector(2356, 16),
15911 => conv_std_logic_vector(2418, 16),
15912 => conv_std_logic_vector(2480, 16),
15913 => conv_std_logic_vector(2542, 16),
15914 => conv_std_logic_vector(2604, 16),
15915 => conv_std_logic_vector(2666, 16),
15916 => conv_std_logic_vector(2728, 16),
15917 => conv_std_logic_vector(2790, 16),
15918 => conv_std_logic_vector(2852, 16),
15919 => conv_std_logic_vector(2914, 16),
15920 => conv_std_logic_vector(2976, 16),
15921 => conv_std_logic_vector(3038, 16),
15922 => conv_std_logic_vector(3100, 16),
15923 => conv_std_logic_vector(3162, 16),
15924 => conv_std_logic_vector(3224, 16),
15925 => conv_std_logic_vector(3286, 16),
15926 => conv_std_logic_vector(3348, 16),
15927 => conv_std_logic_vector(3410, 16),
15928 => conv_std_logic_vector(3472, 16),
15929 => conv_std_logic_vector(3534, 16),
15930 => conv_std_logic_vector(3596, 16),
15931 => conv_std_logic_vector(3658, 16),
15932 => conv_std_logic_vector(3720, 16),
15933 => conv_std_logic_vector(3782, 16),
15934 => conv_std_logic_vector(3844, 16),
15935 => conv_std_logic_vector(3906, 16),
15936 => conv_std_logic_vector(3968, 16),
15937 => conv_std_logic_vector(4030, 16),
15938 => conv_std_logic_vector(4092, 16),
15939 => conv_std_logic_vector(4154, 16),
15940 => conv_std_logic_vector(4216, 16),
15941 => conv_std_logic_vector(4278, 16),
15942 => conv_std_logic_vector(4340, 16),
15943 => conv_std_logic_vector(4402, 16),
15944 => conv_std_logic_vector(4464, 16),
15945 => conv_std_logic_vector(4526, 16),
15946 => conv_std_logic_vector(4588, 16),
15947 => conv_std_logic_vector(4650, 16),
15948 => conv_std_logic_vector(4712, 16),
15949 => conv_std_logic_vector(4774, 16),
15950 => conv_std_logic_vector(4836, 16),
15951 => conv_std_logic_vector(4898, 16),
15952 => conv_std_logic_vector(4960, 16),
15953 => conv_std_logic_vector(5022, 16),
15954 => conv_std_logic_vector(5084, 16),
15955 => conv_std_logic_vector(5146, 16),
15956 => conv_std_logic_vector(5208, 16),
15957 => conv_std_logic_vector(5270, 16),
15958 => conv_std_logic_vector(5332, 16),
15959 => conv_std_logic_vector(5394, 16),
15960 => conv_std_logic_vector(5456, 16),
15961 => conv_std_logic_vector(5518, 16),
15962 => conv_std_logic_vector(5580, 16),
15963 => conv_std_logic_vector(5642, 16),
15964 => conv_std_logic_vector(5704, 16),
15965 => conv_std_logic_vector(5766, 16),
15966 => conv_std_logic_vector(5828, 16),
15967 => conv_std_logic_vector(5890, 16),
15968 => conv_std_logic_vector(5952, 16),
15969 => conv_std_logic_vector(6014, 16),
15970 => conv_std_logic_vector(6076, 16),
15971 => conv_std_logic_vector(6138, 16),
15972 => conv_std_logic_vector(6200, 16),
15973 => conv_std_logic_vector(6262, 16),
15974 => conv_std_logic_vector(6324, 16),
15975 => conv_std_logic_vector(6386, 16),
15976 => conv_std_logic_vector(6448, 16),
15977 => conv_std_logic_vector(6510, 16),
15978 => conv_std_logic_vector(6572, 16),
15979 => conv_std_logic_vector(6634, 16),
15980 => conv_std_logic_vector(6696, 16),
15981 => conv_std_logic_vector(6758, 16),
15982 => conv_std_logic_vector(6820, 16),
15983 => conv_std_logic_vector(6882, 16),
15984 => conv_std_logic_vector(6944, 16),
15985 => conv_std_logic_vector(7006, 16),
15986 => conv_std_logic_vector(7068, 16),
15987 => conv_std_logic_vector(7130, 16),
15988 => conv_std_logic_vector(7192, 16),
15989 => conv_std_logic_vector(7254, 16),
15990 => conv_std_logic_vector(7316, 16),
15991 => conv_std_logic_vector(7378, 16),
15992 => conv_std_logic_vector(7440, 16),
15993 => conv_std_logic_vector(7502, 16),
15994 => conv_std_logic_vector(7564, 16),
15995 => conv_std_logic_vector(7626, 16),
15996 => conv_std_logic_vector(7688, 16),
15997 => conv_std_logic_vector(7750, 16),
15998 => conv_std_logic_vector(7812, 16),
15999 => conv_std_logic_vector(7874, 16),
16000 => conv_std_logic_vector(7936, 16),
16001 => conv_std_logic_vector(7998, 16),
16002 => conv_std_logic_vector(8060, 16),
16003 => conv_std_logic_vector(8122, 16),
16004 => conv_std_logic_vector(8184, 16),
16005 => conv_std_logic_vector(8246, 16),
16006 => conv_std_logic_vector(8308, 16),
16007 => conv_std_logic_vector(8370, 16),
16008 => conv_std_logic_vector(8432, 16),
16009 => conv_std_logic_vector(8494, 16),
16010 => conv_std_logic_vector(8556, 16),
16011 => conv_std_logic_vector(8618, 16),
16012 => conv_std_logic_vector(8680, 16),
16013 => conv_std_logic_vector(8742, 16),
16014 => conv_std_logic_vector(8804, 16),
16015 => conv_std_logic_vector(8866, 16),
16016 => conv_std_logic_vector(8928, 16),
16017 => conv_std_logic_vector(8990, 16),
16018 => conv_std_logic_vector(9052, 16),
16019 => conv_std_logic_vector(9114, 16),
16020 => conv_std_logic_vector(9176, 16),
16021 => conv_std_logic_vector(9238, 16),
16022 => conv_std_logic_vector(9300, 16),
16023 => conv_std_logic_vector(9362, 16),
16024 => conv_std_logic_vector(9424, 16),
16025 => conv_std_logic_vector(9486, 16),
16026 => conv_std_logic_vector(9548, 16),
16027 => conv_std_logic_vector(9610, 16),
16028 => conv_std_logic_vector(9672, 16),
16029 => conv_std_logic_vector(9734, 16),
16030 => conv_std_logic_vector(9796, 16),
16031 => conv_std_logic_vector(9858, 16),
16032 => conv_std_logic_vector(9920, 16),
16033 => conv_std_logic_vector(9982, 16),
16034 => conv_std_logic_vector(10044, 16),
16035 => conv_std_logic_vector(10106, 16),
16036 => conv_std_logic_vector(10168, 16),
16037 => conv_std_logic_vector(10230, 16),
16038 => conv_std_logic_vector(10292, 16),
16039 => conv_std_logic_vector(10354, 16),
16040 => conv_std_logic_vector(10416, 16),
16041 => conv_std_logic_vector(10478, 16),
16042 => conv_std_logic_vector(10540, 16),
16043 => conv_std_logic_vector(10602, 16),
16044 => conv_std_logic_vector(10664, 16),
16045 => conv_std_logic_vector(10726, 16),
16046 => conv_std_logic_vector(10788, 16),
16047 => conv_std_logic_vector(10850, 16),
16048 => conv_std_logic_vector(10912, 16),
16049 => conv_std_logic_vector(10974, 16),
16050 => conv_std_logic_vector(11036, 16),
16051 => conv_std_logic_vector(11098, 16),
16052 => conv_std_logic_vector(11160, 16),
16053 => conv_std_logic_vector(11222, 16),
16054 => conv_std_logic_vector(11284, 16),
16055 => conv_std_logic_vector(11346, 16),
16056 => conv_std_logic_vector(11408, 16),
16057 => conv_std_logic_vector(11470, 16),
16058 => conv_std_logic_vector(11532, 16),
16059 => conv_std_logic_vector(11594, 16),
16060 => conv_std_logic_vector(11656, 16),
16061 => conv_std_logic_vector(11718, 16),
16062 => conv_std_logic_vector(11780, 16),
16063 => conv_std_logic_vector(11842, 16),
16064 => conv_std_logic_vector(11904, 16),
16065 => conv_std_logic_vector(11966, 16),
16066 => conv_std_logic_vector(12028, 16),
16067 => conv_std_logic_vector(12090, 16),
16068 => conv_std_logic_vector(12152, 16),
16069 => conv_std_logic_vector(12214, 16),
16070 => conv_std_logic_vector(12276, 16),
16071 => conv_std_logic_vector(12338, 16),
16072 => conv_std_logic_vector(12400, 16),
16073 => conv_std_logic_vector(12462, 16),
16074 => conv_std_logic_vector(12524, 16),
16075 => conv_std_logic_vector(12586, 16),
16076 => conv_std_logic_vector(12648, 16),
16077 => conv_std_logic_vector(12710, 16),
16078 => conv_std_logic_vector(12772, 16),
16079 => conv_std_logic_vector(12834, 16),
16080 => conv_std_logic_vector(12896, 16),
16081 => conv_std_logic_vector(12958, 16),
16082 => conv_std_logic_vector(13020, 16),
16083 => conv_std_logic_vector(13082, 16),
16084 => conv_std_logic_vector(13144, 16),
16085 => conv_std_logic_vector(13206, 16),
16086 => conv_std_logic_vector(13268, 16),
16087 => conv_std_logic_vector(13330, 16),
16088 => conv_std_logic_vector(13392, 16),
16089 => conv_std_logic_vector(13454, 16),
16090 => conv_std_logic_vector(13516, 16),
16091 => conv_std_logic_vector(13578, 16),
16092 => conv_std_logic_vector(13640, 16),
16093 => conv_std_logic_vector(13702, 16),
16094 => conv_std_logic_vector(13764, 16),
16095 => conv_std_logic_vector(13826, 16),
16096 => conv_std_logic_vector(13888, 16),
16097 => conv_std_logic_vector(13950, 16),
16098 => conv_std_logic_vector(14012, 16),
16099 => conv_std_logic_vector(14074, 16),
16100 => conv_std_logic_vector(14136, 16),
16101 => conv_std_logic_vector(14198, 16),
16102 => conv_std_logic_vector(14260, 16),
16103 => conv_std_logic_vector(14322, 16),
16104 => conv_std_logic_vector(14384, 16),
16105 => conv_std_logic_vector(14446, 16),
16106 => conv_std_logic_vector(14508, 16),
16107 => conv_std_logic_vector(14570, 16),
16108 => conv_std_logic_vector(14632, 16),
16109 => conv_std_logic_vector(14694, 16),
16110 => conv_std_logic_vector(14756, 16),
16111 => conv_std_logic_vector(14818, 16),
16112 => conv_std_logic_vector(14880, 16),
16113 => conv_std_logic_vector(14942, 16),
16114 => conv_std_logic_vector(15004, 16),
16115 => conv_std_logic_vector(15066, 16),
16116 => conv_std_logic_vector(15128, 16),
16117 => conv_std_logic_vector(15190, 16),
16118 => conv_std_logic_vector(15252, 16),
16119 => conv_std_logic_vector(15314, 16),
16120 => conv_std_logic_vector(15376, 16),
16121 => conv_std_logic_vector(15438, 16),
16122 => conv_std_logic_vector(15500, 16),
16123 => conv_std_logic_vector(15562, 16),
16124 => conv_std_logic_vector(15624, 16),
16125 => conv_std_logic_vector(15686, 16),
16126 => conv_std_logic_vector(15748, 16),
16127 => conv_std_logic_vector(15810, 16),
16128 => conv_std_logic_vector(0, 16),
16129 => conv_std_logic_vector(63, 16),
16130 => conv_std_logic_vector(126, 16),
16131 => conv_std_logic_vector(189, 16),
16132 => conv_std_logic_vector(252, 16),
16133 => conv_std_logic_vector(315, 16),
16134 => conv_std_logic_vector(378, 16),
16135 => conv_std_logic_vector(441, 16),
16136 => conv_std_logic_vector(504, 16),
16137 => conv_std_logic_vector(567, 16),
16138 => conv_std_logic_vector(630, 16),
16139 => conv_std_logic_vector(693, 16),
16140 => conv_std_logic_vector(756, 16),
16141 => conv_std_logic_vector(819, 16),
16142 => conv_std_logic_vector(882, 16),
16143 => conv_std_logic_vector(945, 16),
16144 => conv_std_logic_vector(1008, 16),
16145 => conv_std_logic_vector(1071, 16),
16146 => conv_std_logic_vector(1134, 16),
16147 => conv_std_logic_vector(1197, 16),
16148 => conv_std_logic_vector(1260, 16),
16149 => conv_std_logic_vector(1323, 16),
16150 => conv_std_logic_vector(1386, 16),
16151 => conv_std_logic_vector(1449, 16),
16152 => conv_std_logic_vector(1512, 16),
16153 => conv_std_logic_vector(1575, 16),
16154 => conv_std_logic_vector(1638, 16),
16155 => conv_std_logic_vector(1701, 16),
16156 => conv_std_logic_vector(1764, 16),
16157 => conv_std_logic_vector(1827, 16),
16158 => conv_std_logic_vector(1890, 16),
16159 => conv_std_logic_vector(1953, 16),
16160 => conv_std_logic_vector(2016, 16),
16161 => conv_std_logic_vector(2079, 16),
16162 => conv_std_logic_vector(2142, 16),
16163 => conv_std_logic_vector(2205, 16),
16164 => conv_std_logic_vector(2268, 16),
16165 => conv_std_logic_vector(2331, 16),
16166 => conv_std_logic_vector(2394, 16),
16167 => conv_std_logic_vector(2457, 16),
16168 => conv_std_logic_vector(2520, 16),
16169 => conv_std_logic_vector(2583, 16),
16170 => conv_std_logic_vector(2646, 16),
16171 => conv_std_logic_vector(2709, 16),
16172 => conv_std_logic_vector(2772, 16),
16173 => conv_std_logic_vector(2835, 16),
16174 => conv_std_logic_vector(2898, 16),
16175 => conv_std_logic_vector(2961, 16),
16176 => conv_std_logic_vector(3024, 16),
16177 => conv_std_logic_vector(3087, 16),
16178 => conv_std_logic_vector(3150, 16),
16179 => conv_std_logic_vector(3213, 16),
16180 => conv_std_logic_vector(3276, 16),
16181 => conv_std_logic_vector(3339, 16),
16182 => conv_std_logic_vector(3402, 16),
16183 => conv_std_logic_vector(3465, 16),
16184 => conv_std_logic_vector(3528, 16),
16185 => conv_std_logic_vector(3591, 16),
16186 => conv_std_logic_vector(3654, 16),
16187 => conv_std_logic_vector(3717, 16),
16188 => conv_std_logic_vector(3780, 16),
16189 => conv_std_logic_vector(3843, 16),
16190 => conv_std_logic_vector(3906, 16),
16191 => conv_std_logic_vector(3969, 16),
16192 => conv_std_logic_vector(4032, 16),
16193 => conv_std_logic_vector(4095, 16),
16194 => conv_std_logic_vector(4158, 16),
16195 => conv_std_logic_vector(4221, 16),
16196 => conv_std_logic_vector(4284, 16),
16197 => conv_std_logic_vector(4347, 16),
16198 => conv_std_logic_vector(4410, 16),
16199 => conv_std_logic_vector(4473, 16),
16200 => conv_std_logic_vector(4536, 16),
16201 => conv_std_logic_vector(4599, 16),
16202 => conv_std_logic_vector(4662, 16),
16203 => conv_std_logic_vector(4725, 16),
16204 => conv_std_logic_vector(4788, 16),
16205 => conv_std_logic_vector(4851, 16),
16206 => conv_std_logic_vector(4914, 16),
16207 => conv_std_logic_vector(4977, 16),
16208 => conv_std_logic_vector(5040, 16),
16209 => conv_std_logic_vector(5103, 16),
16210 => conv_std_logic_vector(5166, 16),
16211 => conv_std_logic_vector(5229, 16),
16212 => conv_std_logic_vector(5292, 16),
16213 => conv_std_logic_vector(5355, 16),
16214 => conv_std_logic_vector(5418, 16),
16215 => conv_std_logic_vector(5481, 16),
16216 => conv_std_logic_vector(5544, 16),
16217 => conv_std_logic_vector(5607, 16),
16218 => conv_std_logic_vector(5670, 16),
16219 => conv_std_logic_vector(5733, 16),
16220 => conv_std_logic_vector(5796, 16),
16221 => conv_std_logic_vector(5859, 16),
16222 => conv_std_logic_vector(5922, 16),
16223 => conv_std_logic_vector(5985, 16),
16224 => conv_std_logic_vector(6048, 16),
16225 => conv_std_logic_vector(6111, 16),
16226 => conv_std_logic_vector(6174, 16),
16227 => conv_std_logic_vector(6237, 16),
16228 => conv_std_logic_vector(6300, 16),
16229 => conv_std_logic_vector(6363, 16),
16230 => conv_std_logic_vector(6426, 16),
16231 => conv_std_logic_vector(6489, 16),
16232 => conv_std_logic_vector(6552, 16),
16233 => conv_std_logic_vector(6615, 16),
16234 => conv_std_logic_vector(6678, 16),
16235 => conv_std_logic_vector(6741, 16),
16236 => conv_std_logic_vector(6804, 16),
16237 => conv_std_logic_vector(6867, 16),
16238 => conv_std_logic_vector(6930, 16),
16239 => conv_std_logic_vector(6993, 16),
16240 => conv_std_logic_vector(7056, 16),
16241 => conv_std_logic_vector(7119, 16),
16242 => conv_std_logic_vector(7182, 16),
16243 => conv_std_logic_vector(7245, 16),
16244 => conv_std_logic_vector(7308, 16),
16245 => conv_std_logic_vector(7371, 16),
16246 => conv_std_logic_vector(7434, 16),
16247 => conv_std_logic_vector(7497, 16),
16248 => conv_std_logic_vector(7560, 16),
16249 => conv_std_logic_vector(7623, 16),
16250 => conv_std_logic_vector(7686, 16),
16251 => conv_std_logic_vector(7749, 16),
16252 => conv_std_logic_vector(7812, 16),
16253 => conv_std_logic_vector(7875, 16),
16254 => conv_std_logic_vector(7938, 16),
16255 => conv_std_logic_vector(8001, 16),
16256 => conv_std_logic_vector(8064, 16),
16257 => conv_std_logic_vector(8127, 16),
16258 => conv_std_logic_vector(8190, 16),
16259 => conv_std_logic_vector(8253, 16),
16260 => conv_std_logic_vector(8316, 16),
16261 => conv_std_logic_vector(8379, 16),
16262 => conv_std_logic_vector(8442, 16),
16263 => conv_std_logic_vector(8505, 16),
16264 => conv_std_logic_vector(8568, 16),
16265 => conv_std_logic_vector(8631, 16),
16266 => conv_std_logic_vector(8694, 16),
16267 => conv_std_logic_vector(8757, 16),
16268 => conv_std_logic_vector(8820, 16),
16269 => conv_std_logic_vector(8883, 16),
16270 => conv_std_logic_vector(8946, 16),
16271 => conv_std_logic_vector(9009, 16),
16272 => conv_std_logic_vector(9072, 16),
16273 => conv_std_logic_vector(9135, 16),
16274 => conv_std_logic_vector(9198, 16),
16275 => conv_std_logic_vector(9261, 16),
16276 => conv_std_logic_vector(9324, 16),
16277 => conv_std_logic_vector(9387, 16),
16278 => conv_std_logic_vector(9450, 16),
16279 => conv_std_logic_vector(9513, 16),
16280 => conv_std_logic_vector(9576, 16),
16281 => conv_std_logic_vector(9639, 16),
16282 => conv_std_logic_vector(9702, 16),
16283 => conv_std_logic_vector(9765, 16),
16284 => conv_std_logic_vector(9828, 16),
16285 => conv_std_logic_vector(9891, 16),
16286 => conv_std_logic_vector(9954, 16),
16287 => conv_std_logic_vector(10017, 16),
16288 => conv_std_logic_vector(10080, 16),
16289 => conv_std_logic_vector(10143, 16),
16290 => conv_std_logic_vector(10206, 16),
16291 => conv_std_logic_vector(10269, 16),
16292 => conv_std_logic_vector(10332, 16),
16293 => conv_std_logic_vector(10395, 16),
16294 => conv_std_logic_vector(10458, 16),
16295 => conv_std_logic_vector(10521, 16),
16296 => conv_std_logic_vector(10584, 16),
16297 => conv_std_logic_vector(10647, 16),
16298 => conv_std_logic_vector(10710, 16),
16299 => conv_std_logic_vector(10773, 16),
16300 => conv_std_logic_vector(10836, 16),
16301 => conv_std_logic_vector(10899, 16),
16302 => conv_std_logic_vector(10962, 16),
16303 => conv_std_logic_vector(11025, 16),
16304 => conv_std_logic_vector(11088, 16),
16305 => conv_std_logic_vector(11151, 16),
16306 => conv_std_logic_vector(11214, 16),
16307 => conv_std_logic_vector(11277, 16),
16308 => conv_std_logic_vector(11340, 16),
16309 => conv_std_logic_vector(11403, 16),
16310 => conv_std_logic_vector(11466, 16),
16311 => conv_std_logic_vector(11529, 16),
16312 => conv_std_logic_vector(11592, 16),
16313 => conv_std_logic_vector(11655, 16),
16314 => conv_std_logic_vector(11718, 16),
16315 => conv_std_logic_vector(11781, 16),
16316 => conv_std_logic_vector(11844, 16),
16317 => conv_std_logic_vector(11907, 16),
16318 => conv_std_logic_vector(11970, 16),
16319 => conv_std_logic_vector(12033, 16),
16320 => conv_std_logic_vector(12096, 16),
16321 => conv_std_logic_vector(12159, 16),
16322 => conv_std_logic_vector(12222, 16),
16323 => conv_std_logic_vector(12285, 16),
16324 => conv_std_logic_vector(12348, 16),
16325 => conv_std_logic_vector(12411, 16),
16326 => conv_std_logic_vector(12474, 16),
16327 => conv_std_logic_vector(12537, 16),
16328 => conv_std_logic_vector(12600, 16),
16329 => conv_std_logic_vector(12663, 16),
16330 => conv_std_logic_vector(12726, 16),
16331 => conv_std_logic_vector(12789, 16),
16332 => conv_std_logic_vector(12852, 16),
16333 => conv_std_logic_vector(12915, 16),
16334 => conv_std_logic_vector(12978, 16),
16335 => conv_std_logic_vector(13041, 16),
16336 => conv_std_logic_vector(13104, 16),
16337 => conv_std_logic_vector(13167, 16),
16338 => conv_std_logic_vector(13230, 16),
16339 => conv_std_logic_vector(13293, 16),
16340 => conv_std_logic_vector(13356, 16),
16341 => conv_std_logic_vector(13419, 16),
16342 => conv_std_logic_vector(13482, 16),
16343 => conv_std_logic_vector(13545, 16),
16344 => conv_std_logic_vector(13608, 16),
16345 => conv_std_logic_vector(13671, 16),
16346 => conv_std_logic_vector(13734, 16),
16347 => conv_std_logic_vector(13797, 16),
16348 => conv_std_logic_vector(13860, 16),
16349 => conv_std_logic_vector(13923, 16),
16350 => conv_std_logic_vector(13986, 16),
16351 => conv_std_logic_vector(14049, 16),
16352 => conv_std_logic_vector(14112, 16),
16353 => conv_std_logic_vector(14175, 16),
16354 => conv_std_logic_vector(14238, 16),
16355 => conv_std_logic_vector(14301, 16),
16356 => conv_std_logic_vector(14364, 16),
16357 => conv_std_logic_vector(14427, 16),
16358 => conv_std_logic_vector(14490, 16),
16359 => conv_std_logic_vector(14553, 16),
16360 => conv_std_logic_vector(14616, 16),
16361 => conv_std_logic_vector(14679, 16),
16362 => conv_std_logic_vector(14742, 16),
16363 => conv_std_logic_vector(14805, 16),
16364 => conv_std_logic_vector(14868, 16),
16365 => conv_std_logic_vector(14931, 16),
16366 => conv_std_logic_vector(14994, 16),
16367 => conv_std_logic_vector(15057, 16),
16368 => conv_std_logic_vector(15120, 16),
16369 => conv_std_logic_vector(15183, 16),
16370 => conv_std_logic_vector(15246, 16),
16371 => conv_std_logic_vector(15309, 16),
16372 => conv_std_logic_vector(15372, 16),
16373 => conv_std_logic_vector(15435, 16),
16374 => conv_std_logic_vector(15498, 16),
16375 => conv_std_logic_vector(15561, 16),
16376 => conv_std_logic_vector(15624, 16),
16377 => conv_std_logic_vector(15687, 16),
16378 => conv_std_logic_vector(15750, 16),
16379 => conv_std_logic_vector(15813, 16),
16380 => conv_std_logic_vector(15876, 16),
16381 => conv_std_logic_vector(15939, 16),
16382 => conv_std_logic_vector(16002, 16),
16383 => conv_std_logic_vector(16065, 16),
16384 => conv_std_logic_vector(0, 16),
16385 => conv_std_logic_vector(64, 16),
16386 => conv_std_logic_vector(128, 16),
16387 => conv_std_logic_vector(192, 16),
16388 => conv_std_logic_vector(256, 16),
16389 => conv_std_logic_vector(320, 16),
16390 => conv_std_logic_vector(384, 16),
16391 => conv_std_logic_vector(448, 16),
16392 => conv_std_logic_vector(512, 16),
16393 => conv_std_logic_vector(576, 16),
16394 => conv_std_logic_vector(640, 16),
16395 => conv_std_logic_vector(704, 16),
16396 => conv_std_logic_vector(768, 16),
16397 => conv_std_logic_vector(832, 16),
16398 => conv_std_logic_vector(896, 16),
16399 => conv_std_logic_vector(960, 16),
16400 => conv_std_logic_vector(1024, 16),
16401 => conv_std_logic_vector(1088, 16),
16402 => conv_std_logic_vector(1152, 16),
16403 => conv_std_logic_vector(1216, 16),
16404 => conv_std_logic_vector(1280, 16),
16405 => conv_std_logic_vector(1344, 16),
16406 => conv_std_logic_vector(1408, 16),
16407 => conv_std_logic_vector(1472, 16),
16408 => conv_std_logic_vector(1536, 16),
16409 => conv_std_logic_vector(1600, 16),
16410 => conv_std_logic_vector(1664, 16),
16411 => conv_std_logic_vector(1728, 16),
16412 => conv_std_logic_vector(1792, 16),
16413 => conv_std_logic_vector(1856, 16),
16414 => conv_std_logic_vector(1920, 16),
16415 => conv_std_logic_vector(1984, 16),
16416 => conv_std_logic_vector(2048, 16),
16417 => conv_std_logic_vector(2112, 16),
16418 => conv_std_logic_vector(2176, 16),
16419 => conv_std_logic_vector(2240, 16),
16420 => conv_std_logic_vector(2304, 16),
16421 => conv_std_logic_vector(2368, 16),
16422 => conv_std_logic_vector(2432, 16),
16423 => conv_std_logic_vector(2496, 16),
16424 => conv_std_logic_vector(2560, 16),
16425 => conv_std_logic_vector(2624, 16),
16426 => conv_std_logic_vector(2688, 16),
16427 => conv_std_logic_vector(2752, 16),
16428 => conv_std_logic_vector(2816, 16),
16429 => conv_std_logic_vector(2880, 16),
16430 => conv_std_logic_vector(2944, 16),
16431 => conv_std_logic_vector(3008, 16),
16432 => conv_std_logic_vector(3072, 16),
16433 => conv_std_logic_vector(3136, 16),
16434 => conv_std_logic_vector(3200, 16),
16435 => conv_std_logic_vector(3264, 16),
16436 => conv_std_logic_vector(3328, 16),
16437 => conv_std_logic_vector(3392, 16),
16438 => conv_std_logic_vector(3456, 16),
16439 => conv_std_logic_vector(3520, 16),
16440 => conv_std_logic_vector(3584, 16),
16441 => conv_std_logic_vector(3648, 16),
16442 => conv_std_logic_vector(3712, 16),
16443 => conv_std_logic_vector(3776, 16),
16444 => conv_std_logic_vector(3840, 16),
16445 => conv_std_logic_vector(3904, 16),
16446 => conv_std_logic_vector(3968, 16),
16447 => conv_std_logic_vector(4032, 16),
16448 => conv_std_logic_vector(4096, 16),
16449 => conv_std_logic_vector(4160, 16),
16450 => conv_std_logic_vector(4224, 16),
16451 => conv_std_logic_vector(4288, 16),
16452 => conv_std_logic_vector(4352, 16),
16453 => conv_std_logic_vector(4416, 16),
16454 => conv_std_logic_vector(4480, 16),
16455 => conv_std_logic_vector(4544, 16),
16456 => conv_std_logic_vector(4608, 16),
16457 => conv_std_logic_vector(4672, 16),
16458 => conv_std_logic_vector(4736, 16),
16459 => conv_std_logic_vector(4800, 16),
16460 => conv_std_logic_vector(4864, 16),
16461 => conv_std_logic_vector(4928, 16),
16462 => conv_std_logic_vector(4992, 16),
16463 => conv_std_logic_vector(5056, 16),
16464 => conv_std_logic_vector(5120, 16),
16465 => conv_std_logic_vector(5184, 16),
16466 => conv_std_logic_vector(5248, 16),
16467 => conv_std_logic_vector(5312, 16),
16468 => conv_std_logic_vector(5376, 16),
16469 => conv_std_logic_vector(5440, 16),
16470 => conv_std_logic_vector(5504, 16),
16471 => conv_std_logic_vector(5568, 16),
16472 => conv_std_logic_vector(5632, 16),
16473 => conv_std_logic_vector(5696, 16),
16474 => conv_std_logic_vector(5760, 16),
16475 => conv_std_logic_vector(5824, 16),
16476 => conv_std_logic_vector(5888, 16),
16477 => conv_std_logic_vector(5952, 16),
16478 => conv_std_logic_vector(6016, 16),
16479 => conv_std_logic_vector(6080, 16),
16480 => conv_std_logic_vector(6144, 16),
16481 => conv_std_logic_vector(6208, 16),
16482 => conv_std_logic_vector(6272, 16),
16483 => conv_std_logic_vector(6336, 16),
16484 => conv_std_logic_vector(6400, 16),
16485 => conv_std_logic_vector(6464, 16),
16486 => conv_std_logic_vector(6528, 16),
16487 => conv_std_logic_vector(6592, 16),
16488 => conv_std_logic_vector(6656, 16),
16489 => conv_std_logic_vector(6720, 16),
16490 => conv_std_logic_vector(6784, 16),
16491 => conv_std_logic_vector(6848, 16),
16492 => conv_std_logic_vector(6912, 16),
16493 => conv_std_logic_vector(6976, 16),
16494 => conv_std_logic_vector(7040, 16),
16495 => conv_std_logic_vector(7104, 16),
16496 => conv_std_logic_vector(7168, 16),
16497 => conv_std_logic_vector(7232, 16),
16498 => conv_std_logic_vector(7296, 16),
16499 => conv_std_logic_vector(7360, 16),
16500 => conv_std_logic_vector(7424, 16),
16501 => conv_std_logic_vector(7488, 16),
16502 => conv_std_logic_vector(7552, 16),
16503 => conv_std_logic_vector(7616, 16),
16504 => conv_std_logic_vector(7680, 16),
16505 => conv_std_logic_vector(7744, 16),
16506 => conv_std_logic_vector(7808, 16),
16507 => conv_std_logic_vector(7872, 16),
16508 => conv_std_logic_vector(7936, 16),
16509 => conv_std_logic_vector(8000, 16),
16510 => conv_std_logic_vector(8064, 16),
16511 => conv_std_logic_vector(8128, 16),
16512 => conv_std_logic_vector(8192, 16),
16513 => conv_std_logic_vector(8256, 16),
16514 => conv_std_logic_vector(8320, 16),
16515 => conv_std_logic_vector(8384, 16),
16516 => conv_std_logic_vector(8448, 16),
16517 => conv_std_logic_vector(8512, 16),
16518 => conv_std_logic_vector(8576, 16),
16519 => conv_std_logic_vector(8640, 16),
16520 => conv_std_logic_vector(8704, 16),
16521 => conv_std_logic_vector(8768, 16),
16522 => conv_std_logic_vector(8832, 16),
16523 => conv_std_logic_vector(8896, 16),
16524 => conv_std_logic_vector(8960, 16),
16525 => conv_std_logic_vector(9024, 16),
16526 => conv_std_logic_vector(9088, 16),
16527 => conv_std_logic_vector(9152, 16),
16528 => conv_std_logic_vector(9216, 16),
16529 => conv_std_logic_vector(9280, 16),
16530 => conv_std_logic_vector(9344, 16),
16531 => conv_std_logic_vector(9408, 16),
16532 => conv_std_logic_vector(9472, 16),
16533 => conv_std_logic_vector(9536, 16),
16534 => conv_std_logic_vector(9600, 16),
16535 => conv_std_logic_vector(9664, 16),
16536 => conv_std_logic_vector(9728, 16),
16537 => conv_std_logic_vector(9792, 16),
16538 => conv_std_logic_vector(9856, 16),
16539 => conv_std_logic_vector(9920, 16),
16540 => conv_std_logic_vector(9984, 16),
16541 => conv_std_logic_vector(10048, 16),
16542 => conv_std_logic_vector(10112, 16),
16543 => conv_std_logic_vector(10176, 16),
16544 => conv_std_logic_vector(10240, 16),
16545 => conv_std_logic_vector(10304, 16),
16546 => conv_std_logic_vector(10368, 16),
16547 => conv_std_logic_vector(10432, 16),
16548 => conv_std_logic_vector(10496, 16),
16549 => conv_std_logic_vector(10560, 16),
16550 => conv_std_logic_vector(10624, 16),
16551 => conv_std_logic_vector(10688, 16),
16552 => conv_std_logic_vector(10752, 16),
16553 => conv_std_logic_vector(10816, 16),
16554 => conv_std_logic_vector(10880, 16),
16555 => conv_std_logic_vector(10944, 16),
16556 => conv_std_logic_vector(11008, 16),
16557 => conv_std_logic_vector(11072, 16),
16558 => conv_std_logic_vector(11136, 16),
16559 => conv_std_logic_vector(11200, 16),
16560 => conv_std_logic_vector(11264, 16),
16561 => conv_std_logic_vector(11328, 16),
16562 => conv_std_logic_vector(11392, 16),
16563 => conv_std_logic_vector(11456, 16),
16564 => conv_std_logic_vector(11520, 16),
16565 => conv_std_logic_vector(11584, 16),
16566 => conv_std_logic_vector(11648, 16),
16567 => conv_std_logic_vector(11712, 16),
16568 => conv_std_logic_vector(11776, 16),
16569 => conv_std_logic_vector(11840, 16),
16570 => conv_std_logic_vector(11904, 16),
16571 => conv_std_logic_vector(11968, 16),
16572 => conv_std_logic_vector(12032, 16),
16573 => conv_std_logic_vector(12096, 16),
16574 => conv_std_logic_vector(12160, 16),
16575 => conv_std_logic_vector(12224, 16),
16576 => conv_std_logic_vector(12288, 16),
16577 => conv_std_logic_vector(12352, 16),
16578 => conv_std_logic_vector(12416, 16),
16579 => conv_std_logic_vector(12480, 16),
16580 => conv_std_logic_vector(12544, 16),
16581 => conv_std_logic_vector(12608, 16),
16582 => conv_std_logic_vector(12672, 16),
16583 => conv_std_logic_vector(12736, 16),
16584 => conv_std_logic_vector(12800, 16),
16585 => conv_std_logic_vector(12864, 16),
16586 => conv_std_logic_vector(12928, 16),
16587 => conv_std_logic_vector(12992, 16),
16588 => conv_std_logic_vector(13056, 16),
16589 => conv_std_logic_vector(13120, 16),
16590 => conv_std_logic_vector(13184, 16),
16591 => conv_std_logic_vector(13248, 16),
16592 => conv_std_logic_vector(13312, 16),
16593 => conv_std_logic_vector(13376, 16),
16594 => conv_std_logic_vector(13440, 16),
16595 => conv_std_logic_vector(13504, 16),
16596 => conv_std_logic_vector(13568, 16),
16597 => conv_std_logic_vector(13632, 16),
16598 => conv_std_logic_vector(13696, 16),
16599 => conv_std_logic_vector(13760, 16),
16600 => conv_std_logic_vector(13824, 16),
16601 => conv_std_logic_vector(13888, 16),
16602 => conv_std_logic_vector(13952, 16),
16603 => conv_std_logic_vector(14016, 16),
16604 => conv_std_logic_vector(14080, 16),
16605 => conv_std_logic_vector(14144, 16),
16606 => conv_std_logic_vector(14208, 16),
16607 => conv_std_logic_vector(14272, 16),
16608 => conv_std_logic_vector(14336, 16),
16609 => conv_std_logic_vector(14400, 16),
16610 => conv_std_logic_vector(14464, 16),
16611 => conv_std_logic_vector(14528, 16),
16612 => conv_std_logic_vector(14592, 16),
16613 => conv_std_logic_vector(14656, 16),
16614 => conv_std_logic_vector(14720, 16),
16615 => conv_std_logic_vector(14784, 16),
16616 => conv_std_logic_vector(14848, 16),
16617 => conv_std_logic_vector(14912, 16),
16618 => conv_std_logic_vector(14976, 16),
16619 => conv_std_logic_vector(15040, 16),
16620 => conv_std_logic_vector(15104, 16),
16621 => conv_std_logic_vector(15168, 16),
16622 => conv_std_logic_vector(15232, 16),
16623 => conv_std_logic_vector(15296, 16),
16624 => conv_std_logic_vector(15360, 16),
16625 => conv_std_logic_vector(15424, 16),
16626 => conv_std_logic_vector(15488, 16),
16627 => conv_std_logic_vector(15552, 16),
16628 => conv_std_logic_vector(15616, 16),
16629 => conv_std_logic_vector(15680, 16),
16630 => conv_std_logic_vector(15744, 16),
16631 => conv_std_logic_vector(15808, 16),
16632 => conv_std_logic_vector(15872, 16),
16633 => conv_std_logic_vector(15936, 16),
16634 => conv_std_logic_vector(16000, 16),
16635 => conv_std_logic_vector(16064, 16),
16636 => conv_std_logic_vector(16128, 16),
16637 => conv_std_logic_vector(16192, 16),
16638 => conv_std_logic_vector(16256, 16),
16639 => conv_std_logic_vector(16320, 16),
16640 => conv_std_logic_vector(0, 16),
16641 => conv_std_logic_vector(65, 16),
16642 => conv_std_logic_vector(130, 16),
16643 => conv_std_logic_vector(195, 16),
16644 => conv_std_logic_vector(260, 16),
16645 => conv_std_logic_vector(325, 16),
16646 => conv_std_logic_vector(390, 16),
16647 => conv_std_logic_vector(455, 16),
16648 => conv_std_logic_vector(520, 16),
16649 => conv_std_logic_vector(585, 16),
16650 => conv_std_logic_vector(650, 16),
16651 => conv_std_logic_vector(715, 16),
16652 => conv_std_logic_vector(780, 16),
16653 => conv_std_logic_vector(845, 16),
16654 => conv_std_logic_vector(910, 16),
16655 => conv_std_logic_vector(975, 16),
16656 => conv_std_logic_vector(1040, 16),
16657 => conv_std_logic_vector(1105, 16),
16658 => conv_std_logic_vector(1170, 16),
16659 => conv_std_logic_vector(1235, 16),
16660 => conv_std_logic_vector(1300, 16),
16661 => conv_std_logic_vector(1365, 16),
16662 => conv_std_logic_vector(1430, 16),
16663 => conv_std_logic_vector(1495, 16),
16664 => conv_std_logic_vector(1560, 16),
16665 => conv_std_logic_vector(1625, 16),
16666 => conv_std_logic_vector(1690, 16),
16667 => conv_std_logic_vector(1755, 16),
16668 => conv_std_logic_vector(1820, 16),
16669 => conv_std_logic_vector(1885, 16),
16670 => conv_std_logic_vector(1950, 16),
16671 => conv_std_logic_vector(2015, 16),
16672 => conv_std_logic_vector(2080, 16),
16673 => conv_std_logic_vector(2145, 16),
16674 => conv_std_logic_vector(2210, 16),
16675 => conv_std_logic_vector(2275, 16),
16676 => conv_std_logic_vector(2340, 16),
16677 => conv_std_logic_vector(2405, 16),
16678 => conv_std_logic_vector(2470, 16),
16679 => conv_std_logic_vector(2535, 16),
16680 => conv_std_logic_vector(2600, 16),
16681 => conv_std_logic_vector(2665, 16),
16682 => conv_std_logic_vector(2730, 16),
16683 => conv_std_logic_vector(2795, 16),
16684 => conv_std_logic_vector(2860, 16),
16685 => conv_std_logic_vector(2925, 16),
16686 => conv_std_logic_vector(2990, 16),
16687 => conv_std_logic_vector(3055, 16),
16688 => conv_std_logic_vector(3120, 16),
16689 => conv_std_logic_vector(3185, 16),
16690 => conv_std_logic_vector(3250, 16),
16691 => conv_std_logic_vector(3315, 16),
16692 => conv_std_logic_vector(3380, 16),
16693 => conv_std_logic_vector(3445, 16),
16694 => conv_std_logic_vector(3510, 16),
16695 => conv_std_logic_vector(3575, 16),
16696 => conv_std_logic_vector(3640, 16),
16697 => conv_std_logic_vector(3705, 16),
16698 => conv_std_logic_vector(3770, 16),
16699 => conv_std_logic_vector(3835, 16),
16700 => conv_std_logic_vector(3900, 16),
16701 => conv_std_logic_vector(3965, 16),
16702 => conv_std_logic_vector(4030, 16),
16703 => conv_std_logic_vector(4095, 16),
16704 => conv_std_logic_vector(4160, 16),
16705 => conv_std_logic_vector(4225, 16),
16706 => conv_std_logic_vector(4290, 16),
16707 => conv_std_logic_vector(4355, 16),
16708 => conv_std_logic_vector(4420, 16),
16709 => conv_std_logic_vector(4485, 16),
16710 => conv_std_logic_vector(4550, 16),
16711 => conv_std_logic_vector(4615, 16),
16712 => conv_std_logic_vector(4680, 16),
16713 => conv_std_logic_vector(4745, 16),
16714 => conv_std_logic_vector(4810, 16),
16715 => conv_std_logic_vector(4875, 16),
16716 => conv_std_logic_vector(4940, 16),
16717 => conv_std_logic_vector(5005, 16),
16718 => conv_std_logic_vector(5070, 16),
16719 => conv_std_logic_vector(5135, 16),
16720 => conv_std_logic_vector(5200, 16),
16721 => conv_std_logic_vector(5265, 16),
16722 => conv_std_logic_vector(5330, 16),
16723 => conv_std_logic_vector(5395, 16),
16724 => conv_std_logic_vector(5460, 16),
16725 => conv_std_logic_vector(5525, 16),
16726 => conv_std_logic_vector(5590, 16),
16727 => conv_std_logic_vector(5655, 16),
16728 => conv_std_logic_vector(5720, 16),
16729 => conv_std_logic_vector(5785, 16),
16730 => conv_std_logic_vector(5850, 16),
16731 => conv_std_logic_vector(5915, 16),
16732 => conv_std_logic_vector(5980, 16),
16733 => conv_std_logic_vector(6045, 16),
16734 => conv_std_logic_vector(6110, 16),
16735 => conv_std_logic_vector(6175, 16),
16736 => conv_std_logic_vector(6240, 16),
16737 => conv_std_logic_vector(6305, 16),
16738 => conv_std_logic_vector(6370, 16),
16739 => conv_std_logic_vector(6435, 16),
16740 => conv_std_logic_vector(6500, 16),
16741 => conv_std_logic_vector(6565, 16),
16742 => conv_std_logic_vector(6630, 16),
16743 => conv_std_logic_vector(6695, 16),
16744 => conv_std_logic_vector(6760, 16),
16745 => conv_std_logic_vector(6825, 16),
16746 => conv_std_logic_vector(6890, 16),
16747 => conv_std_logic_vector(6955, 16),
16748 => conv_std_logic_vector(7020, 16),
16749 => conv_std_logic_vector(7085, 16),
16750 => conv_std_logic_vector(7150, 16),
16751 => conv_std_logic_vector(7215, 16),
16752 => conv_std_logic_vector(7280, 16),
16753 => conv_std_logic_vector(7345, 16),
16754 => conv_std_logic_vector(7410, 16),
16755 => conv_std_logic_vector(7475, 16),
16756 => conv_std_logic_vector(7540, 16),
16757 => conv_std_logic_vector(7605, 16),
16758 => conv_std_logic_vector(7670, 16),
16759 => conv_std_logic_vector(7735, 16),
16760 => conv_std_logic_vector(7800, 16),
16761 => conv_std_logic_vector(7865, 16),
16762 => conv_std_logic_vector(7930, 16),
16763 => conv_std_logic_vector(7995, 16),
16764 => conv_std_logic_vector(8060, 16),
16765 => conv_std_logic_vector(8125, 16),
16766 => conv_std_logic_vector(8190, 16),
16767 => conv_std_logic_vector(8255, 16),
16768 => conv_std_logic_vector(8320, 16),
16769 => conv_std_logic_vector(8385, 16),
16770 => conv_std_logic_vector(8450, 16),
16771 => conv_std_logic_vector(8515, 16),
16772 => conv_std_logic_vector(8580, 16),
16773 => conv_std_logic_vector(8645, 16),
16774 => conv_std_logic_vector(8710, 16),
16775 => conv_std_logic_vector(8775, 16),
16776 => conv_std_logic_vector(8840, 16),
16777 => conv_std_logic_vector(8905, 16),
16778 => conv_std_logic_vector(8970, 16),
16779 => conv_std_logic_vector(9035, 16),
16780 => conv_std_logic_vector(9100, 16),
16781 => conv_std_logic_vector(9165, 16),
16782 => conv_std_logic_vector(9230, 16),
16783 => conv_std_logic_vector(9295, 16),
16784 => conv_std_logic_vector(9360, 16),
16785 => conv_std_logic_vector(9425, 16),
16786 => conv_std_logic_vector(9490, 16),
16787 => conv_std_logic_vector(9555, 16),
16788 => conv_std_logic_vector(9620, 16),
16789 => conv_std_logic_vector(9685, 16),
16790 => conv_std_logic_vector(9750, 16),
16791 => conv_std_logic_vector(9815, 16),
16792 => conv_std_logic_vector(9880, 16),
16793 => conv_std_logic_vector(9945, 16),
16794 => conv_std_logic_vector(10010, 16),
16795 => conv_std_logic_vector(10075, 16),
16796 => conv_std_logic_vector(10140, 16),
16797 => conv_std_logic_vector(10205, 16),
16798 => conv_std_logic_vector(10270, 16),
16799 => conv_std_logic_vector(10335, 16),
16800 => conv_std_logic_vector(10400, 16),
16801 => conv_std_logic_vector(10465, 16),
16802 => conv_std_logic_vector(10530, 16),
16803 => conv_std_logic_vector(10595, 16),
16804 => conv_std_logic_vector(10660, 16),
16805 => conv_std_logic_vector(10725, 16),
16806 => conv_std_logic_vector(10790, 16),
16807 => conv_std_logic_vector(10855, 16),
16808 => conv_std_logic_vector(10920, 16),
16809 => conv_std_logic_vector(10985, 16),
16810 => conv_std_logic_vector(11050, 16),
16811 => conv_std_logic_vector(11115, 16),
16812 => conv_std_logic_vector(11180, 16),
16813 => conv_std_logic_vector(11245, 16),
16814 => conv_std_logic_vector(11310, 16),
16815 => conv_std_logic_vector(11375, 16),
16816 => conv_std_logic_vector(11440, 16),
16817 => conv_std_logic_vector(11505, 16),
16818 => conv_std_logic_vector(11570, 16),
16819 => conv_std_logic_vector(11635, 16),
16820 => conv_std_logic_vector(11700, 16),
16821 => conv_std_logic_vector(11765, 16),
16822 => conv_std_logic_vector(11830, 16),
16823 => conv_std_logic_vector(11895, 16),
16824 => conv_std_logic_vector(11960, 16),
16825 => conv_std_logic_vector(12025, 16),
16826 => conv_std_logic_vector(12090, 16),
16827 => conv_std_logic_vector(12155, 16),
16828 => conv_std_logic_vector(12220, 16),
16829 => conv_std_logic_vector(12285, 16),
16830 => conv_std_logic_vector(12350, 16),
16831 => conv_std_logic_vector(12415, 16),
16832 => conv_std_logic_vector(12480, 16),
16833 => conv_std_logic_vector(12545, 16),
16834 => conv_std_logic_vector(12610, 16),
16835 => conv_std_logic_vector(12675, 16),
16836 => conv_std_logic_vector(12740, 16),
16837 => conv_std_logic_vector(12805, 16),
16838 => conv_std_logic_vector(12870, 16),
16839 => conv_std_logic_vector(12935, 16),
16840 => conv_std_logic_vector(13000, 16),
16841 => conv_std_logic_vector(13065, 16),
16842 => conv_std_logic_vector(13130, 16),
16843 => conv_std_logic_vector(13195, 16),
16844 => conv_std_logic_vector(13260, 16),
16845 => conv_std_logic_vector(13325, 16),
16846 => conv_std_logic_vector(13390, 16),
16847 => conv_std_logic_vector(13455, 16),
16848 => conv_std_logic_vector(13520, 16),
16849 => conv_std_logic_vector(13585, 16),
16850 => conv_std_logic_vector(13650, 16),
16851 => conv_std_logic_vector(13715, 16),
16852 => conv_std_logic_vector(13780, 16),
16853 => conv_std_logic_vector(13845, 16),
16854 => conv_std_logic_vector(13910, 16),
16855 => conv_std_logic_vector(13975, 16),
16856 => conv_std_logic_vector(14040, 16),
16857 => conv_std_logic_vector(14105, 16),
16858 => conv_std_logic_vector(14170, 16),
16859 => conv_std_logic_vector(14235, 16),
16860 => conv_std_logic_vector(14300, 16),
16861 => conv_std_logic_vector(14365, 16),
16862 => conv_std_logic_vector(14430, 16),
16863 => conv_std_logic_vector(14495, 16),
16864 => conv_std_logic_vector(14560, 16),
16865 => conv_std_logic_vector(14625, 16),
16866 => conv_std_logic_vector(14690, 16),
16867 => conv_std_logic_vector(14755, 16),
16868 => conv_std_logic_vector(14820, 16),
16869 => conv_std_logic_vector(14885, 16),
16870 => conv_std_logic_vector(14950, 16),
16871 => conv_std_logic_vector(15015, 16),
16872 => conv_std_logic_vector(15080, 16),
16873 => conv_std_logic_vector(15145, 16),
16874 => conv_std_logic_vector(15210, 16),
16875 => conv_std_logic_vector(15275, 16),
16876 => conv_std_logic_vector(15340, 16),
16877 => conv_std_logic_vector(15405, 16),
16878 => conv_std_logic_vector(15470, 16),
16879 => conv_std_logic_vector(15535, 16),
16880 => conv_std_logic_vector(15600, 16),
16881 => conv_std_logic_vector(15665, 16),
16882 => conv_std_logic_vector(15730, 16),
16883 => conv_std_logic_vector(15795, 16),
16884 => conv_std_logic_vector(15860, 16),
16885 => conv_std_logic_vector(15925, 16),
16886 => conv_std_logic_vector(15990, 16),
16887 => conv_std_logic_vector(16055, 16),
16888 => conv_std_logic_vector(16120, 16),
16889 => conv_std_logic_vector(16185, 16),
16890 => conv_std_logic_vector(16250, 16),
16891 => conv_std_logic_vector(16315, 16),
16892 => conv_std_logic_vector(16380, 16),
16893 => conv_std_logic_vector(16445, 16),
16894 => conv_std_logic_vector(16510, 16),
16895 => conv_std_logic_vector(16575, 16),
16896 => conv_std_logic_vector(0, 16),
16897 => conv_std_logic_vector(66, 16),
16898 => conv_std_logic_vector(132, 16),
16899 => conv_std_logic_vector(198, 16),
16900 => conv_std_logic_vector(264, 16),
16901 => conv_std_logic_vector(330, 16),
16902 => conv_std_logic_vector(396, 16),
16903 => conv_std_logic_vector(462, 16),
16904 => conv_std_logic_vector(528, 16),
16905 => conv_std_logic_vector(594, 16),
16906 => conv_std_logic_vector(660, 16),
16907 => conv_std_logic_vector(726, 16),
16908 => conv_std_logic_vector(792, 16),
16909 => conv_std_logic_vector(858, 16),
16910 => conv_std_logic_vector(924, 16),
16911 => conv_std_logic_vector(990, 16),
16912 => conv_std_logic_vector(1056, 16),
16913 => conv_std_logic_vector(1122, 16),
16914 => conv_std_logic_vector(1188, 16),
16915 => conv_std_logic_vector(1254, 16),
16916 => conv_std_logic_vector(1320, 16),
16917 => conv_std_logic_vector(1386, 16),
16918 => conv_std_logic_vector(1452, 16),
16919 => conv_std_logic_vector(1518, 16),
16920 => conv_std_logic_vector(1584, 16),
16921 => conv_std_logic_vector(1650, 16),
16922 => conv_std_logic_vector(1716, 16),
16923 => conv_std_logic_vector(1782, 16),
16924 => conv_std_logic_vector(1848, 16),
16925 => conv_std_logic_vector(1914, 16),
16926 => conv_std_logic_vector(1980, 16),
16927 => conv_std_logic_vector(2046, 16),
16928 => conv_std_logic_vector(2112, 16),
16929 => conv_std_logic_vector(2178, 16),
16930 => conv_std_logic_vector(2244, 16),
16931 => conv_std_logic_vector(2310, 16),
16932 => conv_std_logic_vector(2376, 16),
16933 => conv_std_logic_vector(2442, 16),
16934 => conv_std_logic_vector(2508, 16),
16935 => conv_std_logic_vector(2574, 16),
16936 => conv_std_logic_vector(2640, 16),
16937 => conv_std_logic_vector(2706, 16),
16938 => conv_std_logic_vector(2772, 16),
16939 => conv_std_logic_vector(2838, 16),
16940 => conv_std_logic_vector(2904, 16),
16941 => conv_std_logic_vector(2970, 16),
16942 => conv_std_logic_vector(3036, 16),
16943 => conv_std_logic_vector(3102, 16),
16944 => conv_std_logic_vector(3168, 16),
16945 => conv_std_logic_vector(3234, 16),
16946 => conv_std_logic_vector(3300, 16),
16947 => conv_std_logic_vector(3366, 16),
16948 => conv_std_logic_vector(3432, 16),
16949 => conv_std_logic_vector(3498, 16),
16950 => conv_std_logic_vector(3564, 16),
16951 => conv_std_logic_vector(3630, 16),
16952 => conv_std_logic_vector(3696, 16),
16953 => conv_std_logic_vector(3762, 16),
16954 => conv_std_logic_vector(3828, 16),
16955 => conv_std_logic_vector(3894, 16),
16956 => conv_std_logic_vector(3960, 16),
16957 => conv_std_logic_vector(4026, 16),
16958 => conv_std_logic_vector(4092, 16),
16959 => conv_std_logic_vector(4158, 16),
16960 => conv_std_logic_vector(4224, 16),
16961 => conv_std_logic_vector(4290, 16),
16962 => conv_std_logic_vector(4356, 16),
16963 => conv_std_logic_vector(4422, 16),
16964 => conv_std_logic_vector(4488, 16),
16965 => conv_std_logic_vector(4554, 16),
16966 => conv_std_logic_vector(4620, 16),
16967 => conv_std_logic_vector(4686, 16),
16968 => conv_std_logic_vector(4752, 16),
16969 => conv_std_logic_vector(4818, 16),
16970 => conv_std_logic_vector(4884, 16),
16971 => conv_std_logic_vector(4950, 16),
16972 => conv_std_logic_vector(5016, 16),
16973 => conv_std_logic_vector(5082, 16),
16974 => conv_std_logic_vector(5148, 16),
16975 => conv_std_logic_vector(5214, 16),
16976 => conv_std_logic_vector(5280, 16),
16977 => conv_std_logic_vector(5346, 16),
16978 => conv_std_logic_vector(5412, 16),
16979 => conv_std_logic_vector(5478, 16),
16980 => conv_std_logic_vector(5544, 16),
16981 => conv_std_logic_vector(5610, 16),
16982 => conv_std_logic_vector(5676, 16),
16983 => conv_std_logic_vector(5742, 16),
16984 => conv_std_logic_vector(5808, 16),
16985 => conv_std_logic_vector(5874, 16),
16986 => conv_std_logic_vector(5940, 16),
16987 => conv_std_logic_vector(6006, 16),
16988 => conv_std_logic_vector(6072, 16),
16989 => conv_std_logic_vector(6138, 16),
16990 => conv_std_logic_vector(6204, 16),
16991 => conv_std_logic_vector(6270, 16),
16992 => conv_std_logic_vector(6336, 16),
16993 => conv_std_logic_vector(6402, 16),
16994 => conv_std_logic_vector(6468, 16),
16995 => conv_std_logic_vector(6534, 16),
16996 => conv_std_logic_vector(6600, 16),
16997 => conv_std_logic_vector(6666, 16),
16998 => conv_std_logic_vector(6732, 16),
16999 => conv_std_logic_vector(6798, 16),
17000 => conv_std_logic_vector(6864, 16),
17001 => conv_std_logic_vector(6930, 16),
17002 => conv_std_logic_vector(6996, 16),
17003 => conv_std_logic_vector(7062, 16),
17004 => conv_std_logic_vector(7128, 16),
17005 => conv_std_logic_vector(7194, 16),
17006 => conv_std_logic_vector(7260, 16),
17007 => conv_std_logic_vector(7326, 16),
17008 => conv_std_logic_vector(7392, 16),
17009 => conv_std_logic_vector(7458, 16),
17010 => conv_std_logic_vector(7524, 16),
17011 => conv_std_logic_vector(7590, 16),
17012 => conv_std_logic_vector(7656, 16),
17013 => conv_std_logic_vector(7722, 16),
17014 => conv_std_logic_vector(7788, 16),
17015 => conv_std_logic_vector(7854, 16),
17016 => conv_std_logic_vector(7920, 16),
17017 => conv_std_logic_vector(7986, 16),
17018 => conv_std_logic_vector(8052, 16),
17019 => conv_std_logic_vector(8118, 16),
17020 => conv_std_logic_vector(8184, 16),
17021 => conv_std_logic_vector(8250, 16),
17022 => conv_std_logic_vector(8316, 16),
17023 => conv_std_logic_vector(8382, 16),
17024 => conv_std_logic_vector(8448, 16),
17025 => conv_std_logic_vector(8514, 16),
17026 => conv_std_logic_vector(8580, 16),
17027 => conv_std_logic_vector(8646, 16),
17028 => conv_std_logic_vector(8712, 16),
17029 => conv_std_logic_vector(8778, 16),
17030 => conv_std_logic_vector(8844, 16),
17031 => conv_std_logic_vector(8910, 16),
17032 => conv_std_logic_vector(8976, 16),
17033 => conv_std_logic_vector(9042, 16),
17034 => conv_std_logic_vector(9108, 16),
17035 => conv_std_logic_vector(9174, 16),
17036 => conv_std_logic_vector(9240, 16),
17037 => conv_std_logic_vector(9306, 16),
17038 => conv_std_logic_vector(9372, 16),
17039 => conv_std_logic_vector(9438, 16),
17040 => conv_std_logic_vector(9504, 16),
17041 => conv_std_logic_vector(9570, 16),
17042 => conv_std_logic_vector(9636, 16),
17043 => conv_std_logic_vector(9702, 16),
17044 => conv_std_logic_vector(9768, 16),
17045 => conv_std_logic_vector(9834, 16),
17046 => conv_std_logic_vector(9900, 16),
17047 => conv_std_logic_vector(9966, 16),
17048 => conv_std_logic_vector(10032, 16),
17049 => conv_std_logic_vector(10098, 16),
17050 => conv_std_logic_vector(10164, 16),
17051 => conv_std_logic_vector(10230, 16),
17052 => conv_std_logic_vector(10296, 16),
17053 => conv_std_logic_vector(10362, 16),
17054 => conv_std_logic_vector(10428, 16),
17055 => conv_std_logic_vector(10494, 16),
17056 => conv_std_logic_vector(10560, 16),
17057 => conv_std_logic_vector(10626, 16),
17058 => conv_std_logic_vector(10692, 16),
17059 => conv_std_logic_vector(10758, 16),
17060 => conv_std_logic_vector(10824, 16),
17061 => conv_std_logic_vector(10890, 16),
17062 => conv_std_logic_vector(10956, 16),
17063 => conv_std_logic_vector(11022, 16),
17064 => conv_std_logic_vector(11088, 16),
17065 => conv_std_logic_vector(11154, 16),
17066 => conv_std_logic_vector(11220, 16),
17067 => conv_std_logic_vector(11286, 16),
17068 => conv_std_logic_vector(11352, 16),
17069 => conv_std_logic_vector(11418, 16),
17070 => conv_std_logic_vector(11484, 16),
17071 => conv_std_logic_vector(11550, 16),
17072 => conv_std_logic_vector(11616, 16),
17073 => conv_std_logic_vector(11682, 16),
17074 => conv_std_logic_vector(11748, 16),
17075 => conv_std_logic_vector(11814, 16),
17076 => conv_std_logic_vector(11880, 16),
17077 => conv_std_logic_vector(11946, 16),
17078 => conv_std_logic_vector(12012, 16),
17079 => conv_std_logic_vector(12078, 16),
17080 => conv_std_logic_vector(12144, 16),
17081 => conv_std_logic_vector(12210, 16),
17082 => conv_std_logic_vector(12276, 16),
17083 => conv_std_logic_vector(12342, 16),
17084 => conv_std_logic_vector(12408, 16),
17085 => conv_std_logic_vector(12474, 16),
17086 => conv_std_logic_vector(12540, 16),
17087 => conv_std_logic_vector(12606, 16),
17088 => conv_std_logic_vector(12672, 16),
17089 => conv_std_logic_vector(12738, 16),
17090 => conv_std_logic_vector(12804, 16),
17091 => conv_std_logic_vector(12870, 16),
17092 => conv_std_logic_vector(12936, 16),
17093 => conv_std_logic_vector(13002, 16),
17094 => conv_std_logic_vector(13068, 16),
17095 => conv_std_logic_vector(13134, 16),
17096 => conv_std_logic_vector(13200, 16),
17097 => conv_std_logic_vector(13266, 16),
17098 => conv_std_logic_vector(13332, 16),
17099 => conv_std_logic_vector(13398, 16),
17100 => conv_std_logic_vector(13464, 16),
17101 => conv_std_logic_vector(13530, 16),
17102 => conv_std_logic_vector(13596, 16),
17103 => conv_std_logic_vector(13662, 16),
17104 => conv_std_logic_vector(13728, 16),
17105 => conv_std_logic_vector(13794, 16),
17106 => conv_std_logic_vector(13860, 16),
17107 => conv_std_logic_vector(13926, 16),
17108 => conv_std_logic_vector(13992, 16),
17109 => conv_std_logic_vector(14058, 16),
17110 => conv_std_logic_vector(14124, 16),
17111 => conv_std_logic_vector(14190, 16),
17112 => conv_std_logic_vector(14256, 16),
17113 => conv_std_logic_vector(14322, 16),
17114 => conv_std_logic_vector(14388, 16),
17115 => conv_std_logic_vector(14454, 16),
17116 => conv_std_logic_vector(14520, 16),
17117 => conv_std_logic_vector(14586, 16),
17118 => conv_std_logic_vector(14652, 16),
17119 => conv_std_logic_vector(14718, 16),
17120 => conv_std_logic_vector(14784, 16),
17121 => conv_std_logic_vector(14850, 16),
17122 => conv_std_logic_vector(14916, 16),
17123 => conv_std_logic_vector(14982, 16),
17124 => conv_std_logic_vector(15048, 16),
17125 => conv_std_logic_vector(15114, 16),
17126 => conv_std_logic_vector(15180, 16),
17127 => conv_std_logic_vector(15246, 16),
17128 => conv_std_logic_vector(15312, 16),
17129 => conv_std_logic_vector(15378, 16),
17130 => conv_std_logic_vector(15444, 16),
17131 => conv_std_logic_vector(15510, 16),
17132 => conv_std_logic_vector(15576, 16),
17133 => conv_std_logic_vector(15642, 16),
17134 => conv_std_logic_vector(15708, 16),
17135 => conv_std_logic_vector(15774, 16),
17136 => conv_std_logic_vector(15840, 16),
17137 => conv_std_logic_vector(15906, 16),
17138 => conv_std_logic_vector(15972, 16),
17139 => conv_std_logic_vector(16038, 16),
17140 => conv_std_logic_vector(16104, 16),
17141 => conv_std_logic_vector(16170, 16),
17142 => conv_std_logic_vector(16236, 16),
17143 => conv_std_logic_vector(16302, 16),
17144 => conv_std_logic_vector(16368, 16),
17145 => conv_std_logic_vector(16434, 16),
17146 => conv_std_logic_vector(16500, 16),
17147 => conv_std_logic_vector(16566, 16),
17148 => conv_std_logic_vector(16632, 16),
17149 => conv_std_logic_vector(16698, 16),
17150 => conv_std_logic_vector(16764, 16),
17151 => conv_std_logic_vector(16830, 16),
17152 => conv_std_logic_vector(0, 16),
17153 => conv_std_logic_vector(67, 16),
17154 => conv_std_logic_vector(134, 16),
17155 => conv_std_logic_vector(201, 16),
17156 => conv_std_logic_vector(268, 16),
17157 => conv_std_logic_vector(335, 16),
17158 => conv_std_logic_vector(402, 16),
17159 => conv_std_logic_vector(469, 16),
17160 => conv_std_logic_vector(536, 16),
17161 => conv_std_logic_vector(603, 16),
17162 => conv_std_logic_vector(670, 16),
17163 => conv_std_logic_vector(737, 16),
17164 => conv_std_logic_vector(804, 16),
17165 => conv_std_logic_vector(871, 16),
17166 => conv_std_logic_vector(938, 16),
17167 => conv_std_logic_vector(1005, 16),
17168 => conv_std_logic_vector(1072, 16),
17169 => conv_std_logic_vector(1139, 16),
17170 => conv_std_logic_vector(1206, 16),
17171 => conv_std_logic_vector(1273, 16),
17172 => conv_std_logic_vector(1340, 16),
17173 => conv_std_logic_vector(1407, 16),
17174 => conv_std_logic_vector(1474, 16),
17175 => conv_std_logic_vector(1541, 16),
17176 => conv_std_logic_vector(1608, 16),
17177 => conv_std_logic_vector(1675, 16),
17178 => conv_std_logic_vector(1742, 16),
17179 => conv_std_logic_vector(1809, 16),
17180 => conv_std_logic_vector(1876, 16),
17181 => conv_std_logic_vector(1943, 16),
17182 => conv_std_logic_vector(2010, 16),
17183 => conv_std_logic_vector(2077, 16),
17184 => conv_std_logic_vector(2144, 16),
17185 => conv_std_logic_vector(2211, 16),
17186 => conv_std_logic_vector(2278, 16),
17187 => conv_std_logic_vector(2345, 16),
17188 => conv_std_logic_vector(2412, 16),
17189 => conv_std_logic_vector(2479, 16),
17190 => conv_std_logic_vector(2546, 16),
17191 => conv_std_logic_vector(2613, 16),
17192 => conv_std_logic_vector(2680, 16),
17193 => conv_std_logic_vector(2747, 16),
17194 => conv_std_logic_vector(2814, 16),
17195 => conv_std_logic_vector(2881, 16),
17196 => conv_std_logic_vector(2948, 16),
17197 => conv_std_logic_vector(3015, 16),
17198 => conv_std_logic_vector(3082, 16),
17199 => conv_std_logic_vector(3149, 16),
17200 => conv_std_logic_vector(3216, 16),
17201 => conv_std_logic_vector(3283, 16),
17202 => conv_std_logic_vector(3350, 16),
17203 => conv_std_logic_vector(3417, 16),
17204 => conv_std_logic_vector(3484, 16),
17205 => conv_std_logic_vector(3551, 16),
17206 => conv_std_logic_vector(3618, 16),
17207 => conv_std_logic_vector(3685, 16),
17208 => conv_std_logic_vector(3752, 16),
17209 => conv_std_logic_vector(3819, 16),
17210 => conv_std_logic_vector(3886, 16),
17211 => conv_std_logic_vector(3953, 16),
17212 => conv_std_logic_vector(4020, 16),
17213 => conv_std_logic_vector(4087, 16),
17214 => conv_std_logic_vector(4154, 16),
17215 => conv_std_logic_vector(4221, 16),
17216 => conv_std_logic_vector(4288, 16),
17217 => conv_std_logic_vector(4355, 16),
17218 => conv_std_logic_vector(4422, 16),
17219 => conv_std_logic_vector(4489, 16),
17220 => conv_std_logic_vector(4556, 16),
17221 => conv_std_logic_vector(4623, 16),
17222 => conv_std_logic_vector(4690, 16),
17223 => conv_std_logic_vector(4757, 16),
17224 => conv_std_logic_vector(4824, 16),
17225 => conv_std_logic_vector(4891, 16),
17226 => conv_std_logic_vector(4958, 16),
17227 => conv_std_logic_vector(5025, 16),
17228 => conv_std_logic_vector(5092, 16),
17229 => conv_std_logic_vector(5159, 16),
17230 => conv_std_logic_vector(5226, 16),
17231 => conv_std_logic_vector(5293, 16),
17232 => conv_std_logic_vector(5360, 16),
17233 => conv_std_logic_vector(5427, 16),
17234 => conv_std_logic_vector(5494, 16),
17235 => conv_std_logic_vector(5561, 16),
17236 => conv_std_logic_vector(5628, 16),
17237 => conv_std_logic_vector(5695, 16),
17238 => conv_std_logic_vector(5762, 16),
17239 => conv_std_logic_vector(5829, 16),
17240 => conv_std_logic_vector(5896, 16),
17241 => conv_std_logic_vector(5963, 16),
17242 => conv_std_logic_vector(6030, 16),
17243 => conv_std_logic_vector(6097, 16),
17244 => conv_std_logic_vector(6164, 16),
17245 => conv_std_logic_vector(6231, 16),
17246 => conv_std_logic_vector(6298, 16),
17247 => conv_std_logic_vector(6365, 16),
17248 => conv_std_logic_vector(6432, 16),
17249 => conv_std_logic_vector(6499, 16),
17250 => conv_std_logic_vector(6566, 16),
17251 => conv_std_logic_vector(6633, 16),
17252 => conv_std_logic_vector(6700, 16),
17253 => conv_std_logic_vector(6767, 16),
17254 => conv_std_logic_vector(6834, 16),
17255 => conv_std_logic_vector(6901, 16),
17256 => conv_std_logic_vector(6968, 16),
17257 => conv_std_logic_vector(7035, 16),
17258 => conv_std_logic_vector(7102, 16),
17259 => conv_std_logic_vector(7169, 16),
17260 => conv_std_logic_vector(7236, 16),
17261 => conv_std_logic_vector(7303, 16),
17262 => conv_std_logic_vector(7370, 16),
17263 => conv_std_logic_vector(7437, 16),
17264 => conv_std_logic_vector(7504, 16),
17265 => conv_std_logic_vector(7571, 16),
17266 => conv_std_logic_vector(7638, 16),
17267 => conv_std_logic_vector(7705, 16),
17268 => conv_std_logic_vector(7772, 16),
17269 => conv_std_logic_vector(7839, 16),
17270 => conv_std_logic_vector(7906, 16),
17271 => conv_std_logic_vector(7973, 16),
17272 => conv_std_logic_vector(8040, 16),
17273 => conv_std_logic_vector(8107, 16),
17274 => conv_std_logic_vector(8174, 16),
17275 => conv_std_logic_vector(8241, 16),
17276 => conv_std_logic_vector(8308, 16),
17277 => conv_std_logic_vector(8375, 16),
17278 => conv_std_logic_vector(8442, 16),
17279 => conv_std_logic_vector(8509, 16),
17280 => conv_std_logic_vector(8576, 16),
17281 => conv_std_logic_vector(8643, 16),
17282 => conv_std_logic_vector(8710, 16),
17283 => conv_std_logic_vector(8777, 16),
17284 => conv_std_logic_vector(8844, 16),
17285 => conv_std_logic_vector(8911, 16),
17286 => conv_std_logic_vector(8978, 16),
17287 => conv_std_logic_vector(9045, 16),
17288 => conv_std_logic_vector(9112, 16),
17289 => conv_std_logic_vector(9179, 16),
17290 => conv_std_logic_vector(9246, 16),
17291 => conv_std_logic_vector(9313, 16),
17292 => conv_std_logic_vector(9380, 16),
17293 => conv_std_logic_vector(9447, 16),
17294 => conv_std_logic_vector(9514, 16),
17295 => conv_std_logic_vector(9581, 16),
17296 => conv_std_logic_vector(9648, 16),
17297 => conv_std_logic_vector(9715, 16),
17298 => conv_std_logic_vector(9782, 16),
17299 => conv_std_logic_vector(9849, 16),
17300 => conv_std_logic_vector(9916, 16),
17301 => conv_std_logic_vector(9983, 16),
17302 => conv_std_logic_vector(10050, 16),
17303 => conv_std_logic_vector(10117, 16),
17304 => conv_std_logic_vector(10184, 16),
17305 => conv_std_logic_vector(10251, 16),
17306 => conv_std_logic_vector(10318, 16),
17307 => conv_std_logic_vector(10385, 16),
17308 => conv_std_logic_vector(10452, 16),
17309 => conv_std_logic_vector(10519, 16),
17310 => conv_std_logic_vector(10586, 16),
17311 => conv_std_logic_vector(10653, 16),
17312 => conv_std_logic_vector(10720, 16),
17313 => conv_std_logic_vector(10787, 16),
17314 => conv_std_logic_vector(10854, 16),
17315 => conv_std_logic_vector(10921, 16),
17316 => conv_std_logic_vector(10988, 16),
17317 => conv_std_logic_vector(11055, 16),
17318 => conv_std_logic_vector(11122, 16),
17319 => conv_std_logic_vector(11189, 16),
17320 => conv_std_logic_vector(11256, 16),
17321 => conv_std_logic_vector(11323, 16),
17322 => conv_std_logic_vector(11390, 16),
17323 => conv_std_logic_vector(11457, 16),
17324 => conv_std_logic_vector(11524, 16),
17325 => conv_std_logic_vector(11591, 16),
17326 => conv_std_logic_vector(11658, 16),
17327 => conv_std_logic_vector(11725, 16),
17328 => conv_std_logic_vector(11792, 16),
17329 => conv_std_logic_vector(11859, 16),
17330 => conv_std_logic_vector(11926, 16),
17331 => conv_std_logic_vector(11993, 16),
17332 => conv_std_logic_vector(12060, 16),
17333 => conv_std_logic_vector(12127, 16),
17334 => conv_std_logic_vector(12194, 16),
17335 => conv_std_logic_vector(12261, 16),
17336 => conv_std_logic_vector(12328, 16),
17337 => conv_std_logic_vector(12395, 16),
17338 => conv_std_logic_vector(12462, 16),
17339 => conv_std_logic_vector(12529, 16),
17340 => conv_std_logic_vector(12596, 16),
17341 => conv_std_logic_vector(12663, 16),
17342 => conv_std_logic_vector(12730, 16),
17343 => conv_std_logic_vector(12797, 16),
17344 => conv_std_logic_vector(12864, 16),
17345 => conv_std_logic_vector(12931, 16),
17346 => conv_std_logic_vector(12998, 16),
17347 => conv_std_logic_vector(13065, 16),
17348 => conv_std_logic_vector(13132, 16),
17349 => conv_std_logic_vector(13199, 16),
17350 => conv_std_logic_vector(13266, 16),
17351 => conv_std_logic_vector(13333, 16),
17352 => conv_std_logic_vector(13400, 16),
17353 => conv_std_logic_vector(13467, 16),
17354 => conv_std_logic_vector(13534, 16),
17355 => conv_std_logic_vector(13601, 16),
17356 => conv_std_logic_vector(13668, 16),
17357 => conv_std_logic_vector(13735, 16),
17358 => conv_std_logic_vector(13802, 16),
17359 => conv_std_logic_vector(13869, 16),
17360 => conv_std_logic_vector(13936, 16),
17361 => conv_std_logic_vector(14003, 16),
17362 => conv_std_logic_vector(14070, 16),
17363 => conv_std_logic_vector(14137, 16),
17364 => conv_std_logic_vector(14204, 16),
17365 => conv_std_logic_vector(14271, 16),
17366 => conv_std_logic_vector(14338, 16),
17367 => conv_std_logic_vector(14405, 16),
17368 => conv_std_logic_vector(14472, 16),
17369 => conv_std_logic_vector(14539, 16),
17370 => conv_std_logic_vector(14606, 16),
17371 => conv_std_logic_vector(14673, 16),
17372 => conv_std_logic_vector(14740, 16),
17373 => conv_std_logic_vector(14807, 16),
17374 => conv_std_logic_vector(14874, 16),
17375 => conv_std_logic_vector(14941, 16),
17376 => conv_std_logic_vector(15008, 16),
17377 => conv_std_logic_vector(15075, 16),
17378 => conv_std_logic_vector(15142, 16),
17379 => conv_std_logic_vector(15209, 16),
17380 => conv_std_logic_vector(15276, 16),
17381 => conv_std_logic_vector(15343, 16),
17382 => conv_std_logic_vector(15410, 16),
17383 => conv_std_logic_vector(15477, 16),
17384 => conv_std_logic_vector(15544, 16),
17385 => conv_std_logic_vector(15611, 16),
17386 => conv_std_logic_vector(15678, 16),
17387 => conv_std_logic_vector(15745, 16),
17388 => conv_std_logic_vector(15812, 16),
17389 => conv_std_logic_vector(15879, 16),
17390 => conv_std_logic_vector(15946, 16),
17391 => conv_std_logic_vector(16013, 16),
17392 => conv_std_logic_vector(16080, 16),
17393 => conv_std_logic_vector(16147, 16),
17394 => conv_std_logic_vector(16214, 16),
17395 => conv_std_logic_vector(16281, 16),
17396 => conv_std_logic_vector(16348, 16),
17397 => conv_std_logic_vector(16415, 16),
17398 => conv_std_logic_vector(16482, 16),
17399 => conv_std_logic_vector(16549, 16),
17400 => conv_std_logic_vector(16616, 16),
17401 => conv_std_logic_vector(16683, 16),
17402 => conv_std_logic_vector(16750, 16),
17403 => conv_std_logic_vector(16817, 16),
17404 => conv_std_logic_vector(16884, 16),
17405 => conv_std_logic_vector(16951, 16),
17406 => conv_std_logic_vector(17018, 16),
17407 => conv_std_logic_vector(17085, 16),
17408 => conv_std_logic_vector(0, 16),
17409 => conv_std_logic_vector(68, 16),
17410 => conv_std_logic_vector(136, 16),
17411 => conv_std_logic_vector(204, 16),
17412 => conv_std_logic_vector(272, 16),
17413 => conv_std_logic_vector(340, 16),
17414 => conv_std_logic_vector(408, 16),
17415 => conv_std_logic_vector(476, 16),
17416 => conv_std_logic_vector(544, 16),
17417 => conv_std_logic_vector(612, 16),
17418 => conv_std_logic_vector(680, 16),
17419 => conv_std_logic_vector(748, 16),
17420 => conv_std_logic_vector(816, 16),
17421 => conv_std_logic_vector(884, 16),
17422 => conv_std_logic_vector(952, 16),
17423 => conv_std_logic_vector(1020, 16),
17424 => conv_std_logic_vector(1088, 16),
17425 => conv_std_logic_vector(1156, 16),
17426 => conv_std_logic_vector(1224, 16),
17427 => conv_std_logic_vector(1292, 16),
17428 => conv_std_logic_vector(1360, 16),
17429 => conv_std_logic_vector(1428, 16),
17430 => conv_std_logic_vector(1496, 16),
17431 => conv_std_logic_vector(1564, 16),
17432 => conv_std_logic_vector(1632, 16),
17433 => conv_std_logic_vector(1700, 16),
17434 => conv_std_logic_vector(1768, 16),
17435 => conv_std_logic_vector(1836, 16),
17436 => conv_std_logic_vector(1904, 16),
17437 => conv_std_logic_vector(1972, 16),
17438 => conv_std_logic_vector(2040, 16),
17439 => conv_std_logic_vector(2108, 16),
17440 => conv_std_logic_vector(2176, 16),
17441 => conv_std_logic_vector(2244, 16),
17442 => conv_std_logic_vector(2312, 16),
17443 => conv_std_logic_vector(2380, 16),
17444 => conv_std_logic_vector(2448, 16),
17445 => conv_std_logic_vector(2516, 16),
17446 => conv_std_logic_vector(2584, 16),
17447 => conv_std_logic_vector(2652, 16),
17448 => conv_std_logic_vector(2720, 16),
17449 => conv_std_logic_vector(2788, 16),
17450 => conv_std_logic_vector(2856, 16),
17451 => conv_std_logic_vector(2924, 16),
17452 => conv_std_logic_vector(2992, 16),
17453 => conv_std_logic_vector(3060, 16),
17454 => conv_std_logic_vector(3128, 16),
17455 => conv_std_logic_vector(3196, 16),
17456 => conv_std_logic_vector(3264, 16),
17457 => conv_std_logic_vector(3332, 16),
17458 => conv_std_logic_vector(3400, 16),
17459 => conv_std_logic_vector(3468, 16),
17460 => conv_std_logic_vector(3536, 16),
17461 => conv_std_logic_vector(3604, 16),
17462 => conv_std_logic_vector(3672, 16),
17463 => conv_std_logic_vector(3740, 16),
17464 => conv_std_logic_vector(3808, 16),
17465 => conv_std_logic_vector(3876, 16),
17466 => conv_std_logic_vector(3944, 16),
17467 => conv_std_logic_vector(4012, 16),
17468 => conv_std_logic_vector(4080, 16),
17469 => conv_std_logic_vector(4148, 16),
17470 => conv_std_logic_vector(4216, 16),
17471 => conv_std_logic_vector(4284, 16),
17472 => conv_std_logic_vector(4352, 16),
17473 => conv_std_logic_vector(4420, 16),
17474 => conv_std_logic_vector(4488, 16),
17475 => conv_std_logic_vector(4556, 16),
17476 => conv_std_logic_vector(4624, 16),
17477 => conv_std_logic_vector(4692, 16),
17478 => conv_std_logic_vector(4760, 16),
17479 => conv_std_logic_vector(4828, 16),
17480 => conv_std_logic_vector(4896, 16),
17481 => conv_std_logic_vector(4964, 16),
17482 => conv_std_logic_vector(5032, 16),
17483 => conv_std_logic_vector(5100, 16),
17484 => conv_std_logic_vector(5168, 16),
17485 => conv_std_logic_vector(5236, 16),
17486 => conv_std_logic_vector(5304, 16),
17487 => conv_std_logic_vector(5372, 16),
17488 => conv_std_logic_vector(5440, 16),
17489 => conv_std_logic_vector(5508, 16),
17490 => conv_std_logic_vector(5576, 16),
17491 => conv_std_logic_vector(5644, 16),
17492 => conv_std_logic_vector(5712, 16),
17493 => conv_std_logic_vector(5780, 16),
17494 => conv_std_logic_vector(5848, 16),
17495 => conv_std_logic_vector(5916, 16),
17496 => conv_std_logic_vector(5984, 16),
17497 => conv_std_logic_vector(6052, 16),
17498 => conv_std_logic_vector(6120, 16),
17499 => conv_std_logic_vector(6188, 16),
17500 => conv_std_logic_vector(6256, 16),
17501 => conv_std_logic_vector(6324, 16),
17502 => conv_std_logic_vector(6392, 16),
17503 => conv_std_logic_vector(6460, 16),
17504 => conv_std_logic_vector(6528, 16),
17505 => conv_std_logic_vector(6596, 16),
17506 => conv_std_logic_vector(6664, 16),
17507 => conv_std_logic_vector(6732, 16),
17508 => conv_std_logic_vector(6800, 16),
17509 => conv_std_logic_vector(6868, 16),
17510 => conv_std_logic_vector(6936, 16),
17511 => conv_std_logic_vector(7004, 16),
17512 => conv_std_logic_vector(7072, 16),
17513 => conv_std_logic_vector(7140, 16),
17514 => conv_std_logic_vector(7208, 16),
17515 => conv_std_logic_vector(7276, 16),
17516 => conv_std_logic_vector(7344, 16),
17517 => conv_std_logic_vector(7412, 16),
17518 => conv_std_logic_vector(7480, 16),
17519 => conv_std_logic_vector(7548, 16),
17520 => conv_std_logic_vector(7616, 16),
17521 => conv_std_logic_vector(7684, 16),
17522 => conv_std_logic_vector(7752, 16),
17523 => conv_std_logic_vector(7820, 16),
17524 => conv_std_logic_vector(7888, 16),
17525 => conv_std_logic_vector(7956, 16),
17526 => conv_std_logic_vector(8024, 16),
17527 => conv_std_logic_vector(8092, 16),
17528 => conv_std_logic_vector(8160, 16),
17529 => conv_std_logic_vector(8228, 16),
17530 => conv_std_logic_vector(8296, 16),
17531 => conv_std_logic_vector(8364, 16),
17532 => conv_std_logic_vector(8432, 16),
17533 => conv_std_logic_vector(8500, 16),
17534 => conv_std_logic_vector(8568, 16),
17535 => conv_std_logic_vector(8636, 16),
17536 => conv_std_logic_vector(8704, 16),
17537 => conv_std_logic_vector(8772, 16),
17538 => conv_std_logic_vector(8840, 16),
17539 => conv_std_logic_vector(8908, 16),
17540 => conv_std_logic_vector(8976, 16),
17541 => conv_std_logic_vector(9044, 16),
17542 => conv_std_logic_vector(9112, 16),
17543 => conv_std_logic_vector(9180, 16),
17544 => conv_std_logic_vector(9248, 16),
17545 => conv_std_logic_vector(9316, 16),
17546 => conv_std_logic_vector(9384, 16),
17547 => conv_std_logic_vector(9452, 16),
17548 => conv_std_logic_vector(9520, 16),
17549 => conv_std_logic_vector(9588, 16),
17550 => conv_std_logic_vector(9656, 16),
17551 => conv_std_logic_vector(9724, 16),
17552 => conv_std_logic_vector(9792, 16),
17553 => conv_std_logic_vector(9860, 16),
17554 => conv_std_logic_vector(9928, 16),
17555 => conv_std_logic_vector(9996, 16),
17556 => conv_std_logic_vector(10064, 16),
17557 => conv_std_logic_vector(10132, 16),
17558 => conv_std_logic_vector(10200, 16),
17559 => conv_std_logic_vector(10268, 16),
17560 => conv_std_logic_vector(10336, 16),
17561 => conv_std_logic_vector(10404, 16),
17562 => conv_std_logic_vector(10472, 16),
17563 => conv_std_logic_vector(10540, 16),
17564 => conv_std_logic_vector(10608, 16),
17565 => conv_std_logic_vector(10676, 16),
17566 => conv_std_logic_vector(10744, 16),
17567 => conv_std_logic_vector(10812, 16),
17568 => conv_std_logic_vector(10880, 16),
17569 => conv_std_logic_vector(10948, 16),
17570 => conv_std_logic_vector(11016, 16),
17571 => conv_std_logic_vector(11084, 16),
17572 => conv_std_logic_vector(11152, 16),
17573 => conv_std_logic_vector(11220, 16),
17574 => conv_std_logic_vector(11288, 16),
17575 => conv_std_logic_vector(11356, 16),
17576 => conv_std_logic_vector(11424, 16),
17577 => conv_std_logic_vector(11492, 16),
17578 => conv_std_logic_vector(11560, 16),
17579 => conv_std_logic_vector(11628, 16),
17580 => conv_std_logic_vector(11696, 16),
17581 => conv_std_logic_vector(11764, 16),
17582 => conv_std_logic_vector(11832, 16),
17583 => conv_std_logic_vector(11900, 16),
17584 => conv_std_logic_vector(11968, 16),
17585 => conv_std_logic_vector(12036, 16),
17586 => conv_std_logic_vector(12104, 16),
17587 => conv_std_logic_vector(12172, 16),
17588 => conv_std_logic_vector(12240, 16),
17589 => conv_std_logic_vector(12308, 16),
17590 => conv_std_logic_vector(12376, 16),
17591 => conv_std_logic_vector(12444, 16),
17592 => conv_std_logic_vector(12512, 16),
17593 => conv_std_logic_vector(12580, 16),
17594 => conv_std_logic_vector(12648, 16),
17595 => conv_std_logic_vector(12716, 16),
17596 => conv_std_logic_vector(12784, 16),
17597 => conv_std_logic_vector(12852, 16),
17598 => conv_std_logic_vector(12920, 16),
17599 => conv_std_logic_vector(12988, 16),
17600 => conv_std_logic_vector(13056, 16),
17601 => conv_std_logic_vector(13124, 16),
17602 => conv_std_logic_vector(13192, 16),
17603 => conv_std_logic_vector(13260, 16),
17604 => conv_std_logic_vector(13328, 16),
17605 => conv_std_logic_vector(13396, 16),
17606 => conv_std_logic_vector(13464, 16),
17607 => conv_std_logic_vector(13532, 16),
17608 => conv_std_logic_vector(13600, 16),
17609 => conv_std_logic_vector(13668, 16),
17610 => conv_std_logic_vector(13736, 16),
17611 => conv_std_logic_vector(13804, 16),
17612 => conv_std_logic_vector(13872, 16),
17613 => conv_std_logic_vector(13940, 16),
17614 => conv_std_logic_vector(14008, 16),
17615 => conv_std_logic_vector(14076, 16),
17616 => conv_std_logic_vector(14144, 16),
17617 => conv_std_logic_vector(14212, 16),
17618 => conv_std_logic_vector(14280, 16),
17619 => conv_std_logic_vector(14348, 16),
17620 => conv_std_logic_vector(14416, 16),
17621 => conv_std_logic_vector(14484, 16),
17622 => conv_std_logic_vector(14552, 16),
17623 => conv_std_logic_vector(14620, 16),
17624 => conv_std_logic_vector(14688, 16),
17625 => conv_std_logic_vector(14756, 16),
17626 => conv_std_logic_vector(14824, 16),
17627 => conv_std_logic_vector(14892, 16),
17628 => conv_std_logic_vector(14960, 16),
17629 => conv_std_logic_vector(15028, 16),
17630 => conv_std_logic_vector(15096, 16),
17631 => conv_std_logic_vector(15164, 16),
17632 => conv_std_logic_vector(15232, 16),
17633 => conv_std_logic_vector(15300, 16),
17634 => conv_std_logic_vector(15368, 16),
17635 => conv_std_logic_vector(15436, 16),
17636 => conv_std_logic_vector(15504, 16),
17637 => conv_std_logic_vector(15572, 16),
17638 => conv_std_logic_vector(15640, 16),
17639 => conv_std_logic_vector(15708, 16),
17640 => conv_std_logic_vector(15776, 16),
17641 => conv_std_logic_vector(15844, 16),
17642 => conv_std_logic_vector(15912, 16),
17643 => conv_std_logic_vector(15980, 16),
17644 => conv_std_logic_vector(16048, 16),
17645 => conv_std_logic_vector(16116, 16),
17646 => conv_std_logic_vector(16184, 16),
17647 => conv_std_logic_vector(16252, 16),
17648 => conv_std_logic_vector(16320, 16),
17649 => conv_std_logic_vector(16388, 16),
17650 => conv_std_logic_vector(16456, 16),
17651 => conv_std_logic_vector(16524, 16),
17652 => conv_std_logic_vector(16592, 16),
17653 => conv_std_logic_vector(16660, 16),
17654 => conv_std_logic_vector(16728, 16),
17655 => conv_std_logic_vector(16796, 16),
17656 => conv_std_logic_vector(16864, 16),
17657 => conv_std_logic_vector(16932, 16),
17658 => conv_std_logic_vector(17000, 16),
17659 => conv_std_logic_vector(17068, 16),
17660 => conv_std_logic_vector(17136, 16),
17661 => conv_std_logic_vector(17204, 16),
17662 => conv_std_logic_vector(17272, 16),
17663 => conv_std_logic_vector(17340, 16),
17664 => conv_std_logic_vector(0, 16),
17665 => conv_std_logic_vector(69, 16),
17666 => conv_std_logic_vector(138, 16),
17667 => conv_std_logic_vector(207, 16),
17668 => conv_std_logic_vector(276, 16),
17669 => conv_std_logic_vector(345, 16),
17670 => conv_std_logic_vector(414, 16),
17671 => conv_std_logic_vector(483, 16),
17672 => conv_std_logic_vector(552, 16),
17673 => conv_std_logic_vector(621, 16),
17674 => conv_std_logic_vector(690, 16),
17675 => conv_std_logic_vector(759, 16),
17676 => conv_std_logic_vector(828, 16),
17677 => conv_std_logic_vector(897, 16),
17678 => conv_std_logic_vector(966, 16),
17679 => conv_std_logic_vector(1035, 16),
17680 => conv_std_logic_vector(1104, 16),
17681 => conv_std_logic_vector(1173, 16),
17682 => conv_std_logic_vector(1242, 16),
17683 => conv_std_logic_vector(1311, 16),
17684 => conv_std_logic_vector(1380, 16),
17685 => conv_std_logic_vector(1449, 16),
17686 => conv_std_logic_vector(1518, 16),
17687 => conv_std_logic_vector(1587, 16),
17688 => conv_std_logic_vector(1656, 16),
17689 => conv_std_logic_vector(1725, 16),
17690 => conv_std_logic_vector(1794, 16),
17691 => conv_std_logic_vector(1863, 16),
17692 => conv_std_logic_vector(1932, 16),
17693 => conv_std_logic_vector(2001, 16),
17694 => conv_std_logic_vector(2070, 16),
17695 => conv_std_logic_vector(2139, 16),
17696 => conv_std_logic_vector(2208, 16),
17697 => conv_std_logic_vector(2277, 16),
17698 => conv_std_logic_vector(2346, 16),
17699 => conv_std_logic_vector(2415, 16),
17700 => conv_std_logic_vector(2484, 16),
17701 => conv_std_logic_vector(2553, 16),
17702 => conv_std_logic_vector(2622, 16),
17703 => conv_std_logic_vector(2691, 16),
17704 => conv_std_logic_vector(2760, 16),
17705 => conv_std_logic_vector(2829, 16),
17706 => conv_std_logic_vector(2898, 16),
17707 => conv_std_logic_vector(2967, 16),
17708 => conv_std_logic_vector(3036, 16),
17709 => conv_std_logic_vector(3105, 16),
17710 => conv_std_logic_vector(3174, 16),
17711 => conv_std_logic_vector(3243, 16),
17712 => conv_std_logic_vector(3312, 16),
17713 => conv_std_logic_vector(3381, 16),
17714 => conv_std_logic_vector(3450, 16),
17715 => conv_std_logic_vector(3519, 16),
17716 => conv_std_logic_vector(3588, 16),
17717 => conv_std_logic_vector(3657, 16),
17718 => conv_std_logic_vector(3726, 16),
17719 => conv_std_logic_vector(3795, 16),
17720 => conv_std_logic_vector(3864, 16),
17721 => conv_std_logic_vector(3933, 16),
17722 => conv_std_logic_vector(4002, 16),
17723 => conv_std_logic_vector(4071, 16),
17724 => conv_std_logic_vector(4140, 16),
17725 => conv_std_logic_vector(4209, 16),
17726 => conv_std_logic_vector(4278, 16),
17727 => conv_std_logic_vector(4347, 16),
17728 => conv_std_logic_vector(4416, 16),
17729 => conv_std_logic_vector(4485, 16),
17730 => conv_std_logic_vector(4554, 16),
17731 => conv_std_logic_vector(4623, 16),
17732 => conv_std_logic_vector(4692, 16),
17733 => conv_std_logic_vector(4761, 16),
17734 => conv_std_logic_vector(4830, 16),
17735 => conv_std_logic_vector(4899, 16),
17736 => conv_std_logic_vector(4968, 16),
17737 => conv_std_logic_vector(5037, 16),
17738 => conv_std_logic_vector(5106, 16),
17739 => conv_std_logic_vector(5175, 16),
17740 => conv_std_logic_vector(5244, 16),
17741 => conv_std_logic_vector(5313, 16),
17742 => conv_std_logic_vector(5382, 16),
17743 => conv_std_logic_vector(5451, 16),
17744 => conv_std_logic_vector(5520, 16),
17745 => conv_std_logic_vector(5589, 16),
17746 => conv_std_logic_vector(5658, 16),
17747 => conv_std_logic_vector(5727, 16),
17748 => conv_std_logic_vector(5796, 16),
17749 => conv_std_logic_vector(5865, 16),
17750 => conv_std_logic_vector(5934, 16),
17751 => conv_std_logic_vector(6003, 16),
17752 => conv_std_logic_vector(6072, 16),
17753 => conv_std_logic_vector(6141, 16),
17754 => conv_std_logic_vector(6210, 16),
17755 => conv_std_logic_vector(6279, 16),
17756 => conv_std_logic_vector(6348, 16),
17757 => conv_std_logic_vector(6417, 16),
17758 => conv_std_logic_vector(6486, 16),
17759 => conv_std_logic_vector(6555, 16),
17760 => conv_std_logic_vector(6624, 16),
17761 => conv_std_logic_vector(6693, 16),
17762 => conv_std_logic_vector(6762, 16),
17763 => conv_std_logic_vector(6831, 16),
17764 => conv_std_logic_vector(6900, 16),
17765 => conv_std_logic_vector(6969, 16),
17766 => conv_std_logic_vector(7038, 16),
17767 => conv_std_logic_vector(7107, 16),
17768 => conv_std_logic_vector(7176, 16),
17769 => conv_std_logic_vector(7245, 16),
17770 => conv_std_logic_vector(7314, 16),
17771 => conv_std_logic_vector(7383, 16),
17772 => conv_std_logic_vector(7452, 16),
17773 => conv_std_logic_vector(7521, 16),
17774 => conv_std_logic_vector(7590, 16),
17775 => conv_std_logic_vector(7659, 16),
17776 => conv_std_logic_vector(7728, 16),
17777 => conv_std_logic_vector(7797, 16),
17778 => conv_std_logic_vector(7866, 16),
17779 => conv_std_logic_vector(7935, 16),
17780 => conv_std_logic_vector(8004, 16),
17781 => conv_std_logic_vector(8073, 16),
17782 => conv_std_logic_vector(8142, 16),
17783 => conv_std_logic_vector(8211, 16),
17784 => conv_std_logic_vector(8280, 16),
17785 => conv_std_logic_vector(8349, 16),
17786 => conv_std_logic_vector(8418, 16),
17787 => conv_std_logic_vector(8487, 16),
17788 => conv_std_logic_vector(8556, 16),
17789 => conv_std_logic_vector(8625, 16),
17790 => conv_std_logic_vector(8694, 16),
17791 => conv_std_logic_vector(8763, 16),
17792 => conv_std_logic_vector(8832, 16),
17793 => conv_std_logic_vector(8901, 16),
17794 => conv_std_logic_vector(8970, 16),
17795 => conv_std_logic_vector(9039, 16),
17796 => conv_std_logic_vector(9108, 16),
17797 => conv_std_logic_vector(9177, 16),
17798 => conv_std_logic_vector(9246, 16),
17799 => conv_std_logic_vector(9315, 16),
17800 => conv_std_logic_vector(9384, 16),
17801 => conv_std_logic_vector(9453, 16),
17802 => conv_std_logic_vector(9522, 16),
17803 => conv_std_logic_vector(9591, 16),
17804 => conv_std_logic_vector(9660, 16),
17805 => conv_std_logic_vector(9729, 16),
17806 => conv_std_logic_vector(9798, 16),
17807 => conv_std_logic_vector(9867, 16),
17808 => conv_std_logic_vector(9936, 16),
17809 => conv_std_logic_vector(10005, 16),
17810 => conv_std_logic_vector(10074, 16),
17811 => conv_std_logic_vector(10143, 16),
17812 => conv_std_logic_vector(10212, 16),
17813 => conv_std_logic_vector(10281, 16),
17814 => conv_std_logic_vector(10350, 16),
17815 => conv_std_logic_vector(10419, 16),
17816 => conv_std_logic_vector(10488, 16),
17817 => conv_std_logic_vector(10557, 16),
17818 => conv_std_logic_vector(10626, 16),
17819 => conv_std_logic_vector(10695, 16),
17820 => conv_std_logic_vector(10764, 16),
17821 => conv_std_logic_vector(10833, 16),
17822 => conv_std_logic_vector(10902, 16),
17823 => conv_std_logic_vector(10971, 16),
17824 => conv_std_logic_vector(11040, 16),
17825 => conv_std_logic_vector(11109, 16),
17826 => conv_std_logic_vector(11178, 16),
17827 => conv_std_logic_vector(11247, 16),
17828 => conv_std_logic_vector(11316, 16),
17829 => conv_std_logic_vector(11385, 16),
17830 => conv_std_logic_vector(11454, 16),
17831 => conv_std_logic_vector(11523, 16),
17832 => conv_std_logic_vector(11592, 16),
17833 => conv_std_logic_vector(11661, 16),
17834 => conv_std_logic_vector(11730, 16),
17835 => conv_std_logic_vector(11799, 16),
17836 => conv_std_logic_vector(11868, 16),
17837 => conv_std_logic_vector(11937, 16),
17838 => conv_std_logic_vector(12006, 16),
17839 => conv_std_logic_vector(12075, 16),
17840 => conv_std_logic_vector(12144, 16),
17841 => conv_std_logic_vector(12213, 16),
17842 => conv_std_logic_vector(12282, 16),
17843 => conv_std_logic_vector(12351, 16),
17844 => conv_std_logic_vector(12420, 16),
17845 => conv_std_logic_vector(12489, 16),
17846 => conv_std_logic_vector(12558, 16),
17847 => conv_std_logic_vector(12627, 16),
17848 => conv_std_logic_vector(12696, 16),
17849 => conv_std_logic_vector(12765, 16),
17850 => conv_std_logic_vector(12834, 16),
17851 => conv_std_logic_vector(12903, 16),
17852 => conv_std_logic_vector(12972, 16),
17853 => conv_std_logic_vector(13041, 16),
17854 => conv_std_logic_vector(13110, 16),
17855 => conv_std_logic_vector(13179, 16),
17856 => conv_std_logic_vector(13248, 16),
17857 => conv_std_logic_vector(13317, 16),
17858 => conv_std_logic_vector(13386, 16),
17859 => conv_std_logic_vector(13455, 16),
17860 => conv_std_logic_vector(13524, 16),
17861 => conv_std_logic_vector(13593, 16),
17862 => conv_std_logic_vector(13662, 16),
17863 => conv_std_logic_vector(13731, 16),
17864 => conv_std_logic_vector(13800, 16),
17865 => conv_std_logic_vector(13869, 16),
17866 => conv_std_logic_vector(13938, 16),
17867 => conv_std_logic_vector(14007, 16),
17868 => conv_std_logic_vector(14076, 16),
17869 => conv_std_logic_vector(14145, 16),
17870 => conv_std_logic_vector(14214, 16),
17871 => conv_std_logic_vector(14283, 16),
17872 => conv_std_logic_vector(14352, 16),
17873 => conv_std_logic_vector(14421, 16),
17874 => conv_std_logic_vector(14490, 16),
17875 => conv_std_logic_vector(14559, 16),
17876 => conv_std_logic_vector(14628, 16),
17877 => conv_std_logic_vector(14697, 16),
17878 => conv_std_logic_vector(14766, 16),
17879 => conv_std_logic_vector(14835, 16),
17880 => conv_std_logic_vector(14904, 16),
17881 => conv_std_logic_vector(14973, 16),
17882 => conv_std_logic_vector(15042, 16),
17883 => conv_std_logic_vector(15111, 16),
17884 => conv_std_logic_vector(15180, 16),
17885 => conv_std_logic_vector(15249, 16),
17886 => conv_std_logic_vector(15318, 16),
17887 => conv_std_logic_vector(15387, 16),
17888 => conv_std_logic_vector(15456, 16),
17889 => conv_std_logic_vector(15525, 16),
17890 => conv_std_logic_vector(15594, 16),
17891 => conv_std_logic_vector(15663, 16),
17892 => conv_std_logic_vector(15732, 16),
17893 => conv_std_logic_vector(15801, 16),
17894 => conv_std_logic_vector(15870, 16),
17895 => conv_std_logic_vector(15939, 16),
17896 => conv_std_logic_vector(16008, 16),
17897 => conv_std_logic_vector(16077, 16),
17898 => conv_std_logic_vector(16146, 16),
17899 => conv_std_logic_vector(16215, 16),
17900 => conv_std_logic_vector(16284, 16),
17901 => conv_std_logic_vector(16353, 16),
17902 => conv_std_logic_vector(16422, 16),
17903 => conv_std_logic_vector(16491, 16),
17904 => conv_std_logic_vector(16560, 16),
17905 => conv_std_logic_vector(16629, 16),
17906 => conv_std_logic_vector(16698, 16),
17907 => conv_std_logic_vector(16767, 16),
17908 => conv_std_logic_vector(16836, 16),
17909 => conv_std_logic_vector(16905, 16),
17910 => conv_std_logic_vector(16974, 16),
17911 => conv_std_logic_vector(17043, 16),
17912 => conv_std_logic_vector(17112, 16),
17913 => conv_std_logic_vector(17181, 16),
17914 => conv_std_logic_vector(17250, 16),
17915 => conv_std_logic_vector(17319, 16),
17916 => conv_std_logic_vector(17388, 16),
17917 => conv_std_logic_vector(17457, 16),
17918 => conv_std_logic_vector(17526, 16),
17919 => conv_std_logic_vector(17595, 16),
17920 => conv_std_logic_vector(0, 16),
17921 => conv_std_logic_vector(70, 16),
17922 => conv_std_logic_vector(140, 16),
17923 => conv_std_logic_vector(210, 16),
17924 => conv_std_logic_vector(280, 16),
17925 => conv_std_logic_vector(350, 16),
17926 => conv_std_logic_vector(420, 16),
17927 => conv_std_logic_vector(490, 16),
17928 => conv_std_logic_vector(560, 16),
17929 => conv_std_logic_vector(630, 16),
17930 => conv_std_logic_vector(700, 16),
17931 => conv_std_logic_vector(770, 16),
17932 => conv_std_logic_vector(840, 16),
17933 => conv_std_logic_vector(910, 16),
17934 => conv_std_logic_vector(980, 16),
17935 => conv_std_logic_vector(1050, 16),
17936 => conv_std_logic_vector(1120, 16),
17937 => conv_std_logic_vector(1190, 16),
17938 => conv_std_logic_vector(1260, 16),
17939 => conv_std_logic_vector(1330, 16),
17940 => conv_std_logic_vector(1400, 16),
17941 => conv_std_logic_vector(1470, 16),
17942 => conv_std_logic_vector(1540, 16),
17943 => conv_std_logic_vector(1610, 16),
17944 => conv_std_logic_vector(1680, 16),
17945 => conv_std_logic_vector(1750, 16),
17946 => conv_std_logic_vector(1820, 16),
17947 => conv_std_logic_vector(1890, 16),
17948 => conv_std_logic_vector(1960, 16),
17949 => conv_std_logic_vector(2030, 16),
17950 => conv_std_logic_vector(2100, 16),
17951 => conv_std_logic_vector(2170, 16),
17952 => conv_std_logic_vector(2240, 16),
17953 => conv_std_logic_vector(2310, 16),
17954 => conv_std_logic_vector(2380, 16),
17955 => conv_std_logic_vector(2450, 16),
17956 => conv_std_logic_vector(2520, 16),
17957 => conv_std_logic_vector(2590, 16),
17958 => conv_std_logic_vector(2660, 16),
17959 => conv_std_logic_vector(2730, 16),
17960 => conv_std_logic_vector(2800, 16),
17961 => conv_std_logic_vector(2870, 16),
17962 => conv_std_logic_vector(2940, 16),
17963 => conv_std_logic_vector(3010, 16),
17964 => conv_std_logic_vector(3080, 16),
17965 => conv_std_logic_vector(3150, 16),
17966 => conv_std_logic_vector(3220, 16),
17967 => conv_std_logic_vector(3290, 16),
17968 => conv_std_logic_vector(3360, 16),
17969 => conv_std_logic_vector(3430, 16),
17970 => conv_std_logic_vector(3500, 16),
17971 => conv_std_logic_vector(3570, 16),
17972 => conv_std_logic_vector(3640, 16),
17973 => conv_std_logic_vector(3710, 16),
17974 => conv_std_logic_vector(3780, 16),
17975 => conv_std_logic_vector(3850, 16),
17976 => conv_std_logic_vector(3920, 16),
17977 => conv_std_logic_vector(3990, 16),
17978 => conv_std_logic_vector(4060, 16),
17979 => conv_std_logic_vector(4130, 16),
17980 => conv_std_logic_vector(4200, 16),
17981 => conv_std_logic_vector(4270, 16),
17982 => conv_std_logic_vector(4340, 16),
17983 => conv_std_logic_vector(4410, 16),
17984 => conv_std_logic_vector(4480, 16),
17985 => conv_std_logic_vector(4550, 16),
17986 => conv_std_logic_vector(4620, 16),
17987 => conv_std_logic_vector(4690, 16),
17988 => conv_std_logic_vector(4760, 16),
17989 => conv_std_logic_vector(4830, 16),
17990 => conv_std_logic_vector(4900, 16),
17991 => conv_std_logic_vector(4970, 16),
17992 => conv_std_logic_vector(5040, 16),
17993 => conv_std_logic_vector(5110, 16),
17994 => conv_std_logic_vector(5180, 16),
17995 => conv_std_logic_vector(5250, 16),
17996 => conv_std_logic_vector(5320, 16),
17997 => conv_std_logic_vector(5390, 16),
17998 => conv_std_logic_vector(5460, 16),
17999 => conv_std_logic_vector(5530, 16),
18000 => conv_std_logic_vector(5600, 16),
18001 => conv_std_logic_vector(5670, 16),
18002 => conv_std_logic_vector(5740, 16),
18003 => conv_std_logic_vector(5810, 16),
18004 => conv_std_logic_vector(5880, 16),
18005 => conv_std_logic_vector(5950, 16),
18006 => conv_std_logic_vector(6020, 16),
18007 => conv_std_logic_vector(6090, 16),
18008 => conv_std_logic_vector(6160, 16),
18009 => conv_std_logic_vector(6230, 16),
18010 => conv_std_logic_vector(6300, 16),
18011 => conv_std_logic_vector(6370, 16),
18012 => conv_std_logic_vector(6440, 16),
18013 => conv_std_logic_vector(6510, 16),
18014 => conv_std_logic_vector(6580, 16),
18015 => conv_std_logic_vector(6650, 16),
18016 => conv_std_logic_vector(6720, 16),
18017 => conv_std_logic_vector(6790, 16),
18018 => conv_std_logic_vector(6860, 16),
18019 => conv_std_logic_vector(6930, 16),
18020 => conv_std_logic_vector(7000, 16),
18021 => conv_std_logic_vector(7070, 16),
18022 => conv_std_logic_vector(7140, 16),
18023 => conv_std_logic_vector(7210, 16),
18024 => conv_std_logic_vector(7280, 16),
18025 => conv_std_logic_vector(7350, 16),
18026 => conv_std_logic_vector(7420, 16),
18027 => conv_std_logic_vector(7490, 16),
18028 => conv_std_logic_vector(7560, 16),
18029 => conv_std_logic_vector(7630, 16),
18030 => conv_std_logic_vector(7700, 16),
18031 => conv_std_logic_vector(7770, 16),
18032 => conv_std_logic_vector(7840, 16),
18033 => conv_std_logic_vector(7910, 16),
18034 => conv_std_logic_vector(7980, 16),
18035 => conv_std_logic_vector(8050, 16),
18036 => conv_std_logic_vector(8120, 16),
18037 => conv_std_logic_vector(8190, 16),
18038 => conv_std_logic_vector(8260, 16),
18039 => conv_std_logic_vector(8330, 16),
18040 => conv_std_logic_vector(8400, 16),
18041 => conv_std_logic_vector(8470, 16),
18042 => conv_std_logic_vector(8540, 16),
18043 => conv_std_logic_vector(8610, 16),
18044 => conv_std_logic_vector(8680, 16),
18045 => conv_std_logic_vector(8750, 16),
18046 => conv_std_logic_vector(8820, 16),
18047 => conv_std_logic_vector(8890, 16),
18048 => conv_std_logic_vector(8960, 16),
18049 => conv_std_logic_vector(9030, 16),
18050 => conv_std_logic_vector(9100, 16),
18051 => conv_std_logic_vector(9170, 16),
18052 => conv_std_logic_vector(9240, 16),
18053 => conv_std_logic_vector(9310, 16),
18054 => conv_std_logic_vector(9380, 16),
18055 => conv_std_logic_vector(9450, 16),
18056 => conv_std_logic_vector(9520, 16),
18057 => conv_std_logic_vector(9590, 16),
18058 => conv_std_logic_vector(9660, 16),
18059 => conv_std_logic_vector(9730, 16),
18060 => conv_std_logic_vector(9800, 16),
18061 => conv_std_logic_vector(9870, 16),
18062 => conv_std_logic_vector(9940, 16),
18063 => conv_std_logic_vector(10010, 16),
18064 => conv_std_logic_vector(10080, 16),
18065 => conv_std_logic_vector(10150, 16),
18066 => conv_std_logic_vector(10220, 16),
18067 => conv_std_logic_vector(10290, 16),
18068 => conv_std_logic_vector(10360, 16),
18069 => conv_std_logic_vector(10430, 16),
18070 => conv_std_logic_vector(10500, 16),
18071 => conv_std_logic_vector(10570, 16),
18072 => conv_std_logic_vector(10640, 16),
18073 => conv_std_logic_vector(10710, 16),
18074 => conv_std_logic_vector(10780, 16),
18075 => conv_std_logic_vector(10850, 16),
18076 => conv_std_logic_vector(10920, 16),
18077 => conv_std_logic_vector(10990, 16),
18078 => conv_std_logic_vector(11060, 16),
18079 => conv_std_logic_vector(11130, 16),
18080 => conv_std_logic_vector(11200, 16),
18081 => conv_std_logic_vector(11270, 16),
18082 => conv_std_logic_vector(11340, 16),
18083 => conv_std_logic_vector(11410, 16),
18084 => conv_std_logic_vector(11480, 16),
18085 => conv_std_logic_vector(11550, 16),
18086 => conv_std_logic_vector(11620, 16),
18087 => conv_std_logic_vector(11690, 16),
18088 => conv_std_logic_vector(11760, 16),
18089 => conv_std_logic_vector(11830, 16),
18090 => conv_std_logic_vector(11900, 16),
18091 => conv_std_logic_vector(11970, 16),
18092 => conv_std_logic_vector(12040, 16),
18093 => conv_std_logic_vector(12110, 16),
18094 => conv_std_logic_vector(12180, 16),
18095 => conv_std_logic_vector(12250, 16),
18096 => conv_std_logic_vector(12320, 16),
18097 => conv_std_logic_vector(12390, 16),
18098 => conv_std_logic_vector(12460, 16),
18099 => conv_std_logic_vector(12530, 16),
18100 => conv_std_logic_vector(12600, 16),
18101 => conv_std_logic_vector(12670, 16),
18102 => conv_std_logic_vector(12740, 16),
18103 => conv_std_logic_vector(12810, 16),
18104 => conv_std_logic_vector(12880, 16),
18105 => conv_std_logic_vector(12950, 16),
18106 => conv_std_logic_vector(13020, 16),
18107 => conv_std_logic_vector(13090, 16),
18108 => conv_std_logic_vector(13160, 16),
18109 => conv_std_logic_vector(13230, 16),
18110 => conv_std_logic_vector(13300, 16),
18111 => conv_std_logic_vector(13370, 16),
18112 => conv_std_logic_vector(13440, 16),
18113 => conv_std_logic_vector(13510, 16),
18114 => conv_std_logic_vector(13580, 16),
18115 => conv_std_logic_vector(13650, 16),
18116 => conv_std_logic_vector(13720, 16),
18117 => conv_std_logic_vector(13790, 16),
18118 => conv_std_logic_vector(13860, 16),
18119 => conv_std_logic_vector(13930, 16),
18120 => conv_std_logic_vector(14000, 16),
18121 => conv_std_logic_vector(14070, 16),
18122 => conv_std_logic_vector(14140, 16),
18123 => conv_std_logic_vector(14210, 16),
18124 => conv_std_logic_vector(14280, 16),
18125 => conv_std_logic_vector(14350, 16),
18126 => conv_std_logic_vector(14420, 16),
18127 => conv_std_logic_vector(14490, 16),
18128 => conv_std_logic_vector(14560, 16),
18129 => conv_std_logic_vector(14630, 16),
18130 => conv_std_logic_vector(14700, 16),
18131 => conv_std_logic_vector(14770, 16),
18132 => conv_std_logic_vector(14840, 16),
18133 => conv_std_logic_vector(14910, 16),
18134 => conv_std_logic_vector(14980, 16),
18135 => conv_std_logic_vector(15050, 16),
18136 => conv_std_logic_vector(15120, 16),
18137 => conv_std_logic_vector(15190, 16),
18138 => conv_std_logic_vector(15260, 16),
18139 => conv_std_logic_vector(15330, 16),
18140 => conv_std_logic_vector(15400, 16),
18141 => conv_std_logic_vector(15470, 16),
18142 => conv_std_logic_vector(15540, 16),
18143 => conv_std_logic_vector(15610, 16),
18144 => conv_std_logic_vector(15680, 16),
18145 => conv_std_logic_vector(15750, 16),
18146 => conv_std_logic_vector(15820, 16),
18147 => conv_std_logic_vector(15890, 16),
18148 => conv_std_logic_vector(15960, 16),
18149 => conv_std_logic_vector(16030, 16),
18150 => conv_std_logic_vector(16100, 16),
18151 => conv_std_logic_vector(16170, 16),
18152 => conv_std_logic_vector(16240, 16),
18153 => conv_std_logic_vector(16310, 16),
18154 => conv_std_logic_vector(16380, 16),
18155 => conv_std_logic_vector(16450, 16),
18156 => conv_std_logic_vector(16520, 16),
18157 => conv_std_logic_vector(16590, 16),
18158 => conv_std_logic_vector(16660, 16),
18159 => conv_std_logic_vector(16730, 16),
18160 => conv_std_logic_vector(16800, 16),
18161 => conv_std_logic_vector(16870, 16),
18162 => conv_std_logic_vector(16940, 16),
18163 => conv_std_logic_vector(17010, 16),
18164 => conv_std_logic_vector(17080, 16),
18165 => conv_std_logic_vector(17150, 16),
18166 => conv_std_logic_vector(17220, 16),
18167 => conv_std_logic_vector(17290, 16),
18168 => conv_std_logic_vector(17360, 16),
18169 => conv_std_logic_vector(17430, 16),
18170 => conv_std_logic_vector(17500, 16),
18171 => conv_std_logic_vector(17570, 16),
18172 => conv_std_logic_vector(17640, 16),
18173 => conv_std_logic_vector(17710, 16),
18174 => conv_std_logic_vector(17780, 16),
18175 => conv_std_logic_vector(17850, 16),
18176 => conv_std_logic_vector(0, 16),
18177 => conv_std_logic_vector(71, 16),
18178 => conv_std_logic_vector(142, 16),
18179 => conv_std_logic_vector(213, 16),
18180 => conv_std_logic_vector(284, 16),
18181 => conv_std_logic_vector(355, 16),
18182 => conv_std_logic_vector(426, 16),
18183 => conv_std_logic_vector(497, 16),
18184 => conv_std_logic_vector(568, 16),
18185 => conv_std_logic_vector(639, 16),
18186 => conv_std_logic_vector(710, 16),
18187 => conv_std_logic_vector(781, 16),
18188 => conv_std_logic_vector(852, 16),
18189 => conv_std_logic_vector(923, 16),
18190 => conv_std_logic_vector(994, 16),
18191 => conv_std_logic_vector(1065, 16),
18192 => conv_std_logic_vector(1136, 16),
18193 => conv_std_logic_vector(1207, 16),
18194 => conv_std_logic_vector(1278, 16),
18195 => conv_std_logic_vector(1349, 16),
18196 => conv_std_logic_vector(1420, 16),
18197 => conv_std_logic_vector(1491, 16),
18198 => conv_std_logic_vector(1562, 16),
18199 => conv_std_logic_vector(1633, 16),
18200 => conv_std_logic_vector(1704, 16),
18201 => conv_std_logic_vector(1775, 16),
18202 => conv_std_logic_vector(1846, 16),
18203 => conv_std_logic_vector(1917, 16),
18204 => conv_std_logic_vector(1988, 16),
18205 => conv_std_logic_vector(2059, 16),
18206 => conv_std_logic_vector(2130, 16),
18207 => conv_std_logic_vector(2201, 16),
18208 => conv_std_logic_vector(2272, 16),
18209 => conv_std_logic_vector(2343, 16),
18210 => conv_std_logic_vector(2414, 16),
18211 => conv_std_logic_vector(2485, 16),
18212 => conv_std_logic_vector(2556, 16),
18213 => conv_std_logic_vector(2627, 16),
18214 => conv_std_logic_vector(2698, 16),
18215 => conv_std_logic_vector(2769, 16),
18216 => conv_std_logic_vector(2840, 16),
18217 => conv_std_logic_vector(2911, 16),
18218 => conv_std_logic_vector(2982, 16),
18219 => conv_std_logic_vector(3053, 16),
18220 => conv_std_logic_vector(3124, 16),
18221 => conv_std_logic_vector(3195, 16),
18222 => conv_std_logic_vector(3266, 16),
18223 => conv_std_logic_vector(3337, 16),
18224 => conv_std_logic_vector(3408, 16),
18225 => conv_std_logic_vector(3479, 16),
18226 => conv_std_logic_vector(3550, 16),
18227 => conv_std_logic_vector(3621, 16),
18228 => conv_std_logic_vector(3692, 16),
18229 => conv_std_logic_vector(3763, 16),
18230 => conv_std_logic_vector(3834, 16),
18231 => conv_std_logic_vector(3905, 16),
18232 => conv_std_logic_vector(3976, 16),
18233 => conv_std_logic_vector(4047, 16),
18234 => conv_std_logic_vector(4118, 16),
18235 => conv_std_logic_vector(4189, 16),
18236 => conv_std_logic_vector(4260, 16),
18237 => conv_std_logic_vector(4331, 16),
18238 => conv_std_logic_vector(4402, 16),
18239 => conv_std_logic_vector(4473, 16),
18240 => conv_std_logic_vector(4544, 16),
18241 => conv_std_logic_vector(4615, 16),
18242 => conv_std_logic_vector(4686, 16),
18243 => conv_std_logic_vector(4757, 16),
18244 => conv_std_logic_vector(4828, 16),
18245 => conv_std_logic_vector(4899, 16),
18246 => conv_std_logic_vector(4970, 16),
18247 => conv_std_logic_vector(5041, 16),
18248 => conv_std_logic_vector(5112, 16),
18249 => conv_std_logic_vector(5183, 16),
18250 => conv_std_logic_vector(5254, 16),
18251 => conv_std_logic_vector(5325, 16),
18252 => conv_std_logic_vector(5396, 16),
18253 => conv_std_logic_vector(5467, 16),
18254 => conv_std_logic_vector(5538, 16),
18255 => conv_std_logic_vector(5609, 16),
18256 => conv_std_logic_vector(5680, 16),
18257 => conv_std_logic_vector(5751, 16),
18258 => conv_std_logic_vector(5822, 16),
18259 => conv_std_logic_vector(5893, 16),
18260 => conv_std_logic_vector(5964, 16),
18261 => conv_std_logic_vector(6035, 16),
18262 => conv_std_logic_vector(6106, 16),
18263 => conv_std_logic_vector(6177, 16),
18264 => conv_std_logic_vector(6248, 16),
18265 => conv_std_logic_vector(6319, 16),
18266 => conv_std_logic_vector(6390, 16),
18267 => conv_std_logic_vector(6461, 16),
18268 => conv_std_logic_vector(6532, 16),
18269 => conv_std_logic_vector(6603, 16),
18270 => conv_std_logic_vector(6674, 16),
18271 => conv_std_logic_vector(6745, 16),
18272 => conv_std_logic_vector(6816, 16),
18273 => conv_std_logic_vector(6887, 16),
18274 => conv_std_logic_vector(6958, 16),
18275 => conv_std_logic_vector(7029, 16),
18276 => conv_std_logic_vector(7100, 16),
18277 => conv_std_logic_vector(7171, 16),
18278 => conv_std_logic_vector(7242, 16),
18279 => conv_std_logic_vector(7313, 16),
18280 => conv_std_logic_vector(7384, 16),
18281 => conv_std_logic_vector(7455, 16),
18282 => conv_std_logic_vector(7526, 16),
18283 => conv_std_logic_vector(7597, 16),
18284 => conv_std_logic_vector(7668, 16),
18285 => conv_std_logic_vector(7739, 16),
18286 => conv_std_logic_vector(7810, 16),
18287 => conv_std_logic_vector(7881, 16),
18288 => conv_std_logic_vector(7952, 16),
18289 => conv_std_logic_vector(8023, 16),
18290 => conv_std_logic_vector(8094, 16),
18291 => conv_std_logic_vector(8165, 16),
18292 => conv_std_logic_vector(8236, 16),
18293 => conv_std_logic_vector(8307, 16),
18294 => conv_std_logic_vector(8378, 16),
18295 => conv_std_logic_vector(8449, 16),
18296 => conv_std_logic_vector(8520, 16),
18297 => conv_std_logic_vector(8591, 16),
18298 => conv_std_logic_vector(8662, 16),
18299 => conv_std_logic_vector(8733, 16),
18300 => conv_std_logic_vector(8804, 16),
18301 => conv_std_logic_vector(8875, 16),
18302 => conv_std_logic_vector(8946, 16),
18303 => conv_std_logic_vector(9017, 16),
18304 => conv_std_logic_vector(9088, 16),
18305 => conv_std_logic_vector(9159, 16),
18306 => conv_std_logic_vector(9230, 16),
18307 => conv_std_logic_vector(9301, 16),
18308 => conv_std_logic_vector(9372, 16),
18309 => conv_std_logic_vector(9443, 16),
18310 => conv_std_logic_vector(9514, 16),
18311 => conv_std_logic_vector(9585, 16),
18312 => conv_std_logic_vector(9656, 16),
18313 => conv_std_logic_vector(9727, 16),
18314 => conv_std_logic_vector(9798, 16),
18315 => conv_std_logic_vector(9869, 16),
18316 => conv_std_logic_vector(9940, 16),
18317 => conv_std_logic_vector(10011, 16),
18318 => conv_std_logic_vector(10082, 16),
18319 => conv_std_logic_vector(10153, 16),
18320 => conv_std_logic_vector(10224, 16),
18321 => conv_std_logic_vector(10295, 16),
18322 => conv_std_logic_vector(10366, 16),
18323 => conv_std_logic_vector(10437, 16),
18324 => conv_std_logic_vector(10508, 16),
18325 => conv_std_logic_vector(10579, 16),
18326 => conv_std_logic_vector(10650, 16),
18327 => conv_std_logic_vector(10721, 16),
18328 => conv_std_logic_vector(10792, 16),
18329 => conv_std_logic_vector(10863, 16),
18330 => conv_std_logic_vector(10934, 16),
18331 => conv_std_logic_vector(11005, 16),
18332 => conv_std_logic_vector(11076, 16),
18333 => conv_std_logic_vector(11147, 16),
18334 => conv_std_logic_vector(11218, 16),
18335 => conv_std_logic_vector(11289, 16),
18336 => conv_std_logic_vector(11360, 16),
18337 => conv_std_logic_vector(11431, 16),
18338 => conv_std_logic_vector(11502, 16),
18339 => conv_std_logic_vector(11573, 16),
18340 => conv_std_logic_vector(11644, 16),
18341 => conv_std_logic_vector(11715, 16),
18342 => conv_std_logic_vector(11786, 16),
18343 => conv_std_logic_vector(11857, 16),
18344 => conv_std_logic_vector(11928, 16),
18345 => conv_std_logic_vector(11999, 16),
18346 => conv_std_logic_vector(12070, 16),
18347 => conv_std_logic_vector(12141, 16),
18348 => conv_std_logic_vector(12212, 16),
18349 => conv_std_logic_vector(12283, 16),
18350 => conv_std_logic_vector(12354, 16),
18351 => conv_std_logic_vector(12425, 16),
18352 => conv_std_logic_vector(12496, 16),
18353 => conv_std_logic_vector(12567, 16),
18354 => conv_std_logic_vector(12638, 16),
18355 => conv_std_logic_vector(12709, 16),
18356 => conv_std_logic_vector(12780, 16),
18357 => conv_std_logic_vector(12851, 16),
18358 => conv_std_logic_vector(12922, 16),
18359 => conv_std_logic_vector(12993, 16),
18360 => conv_std_logic_vector(13064, 16),
18361 => conv_std_logic_vector(13135, 16),
18362 => conv_std_logic_vector(13206, 16),
18363 => conv_std_logic_vector(13277, 16),
18364 => conv_std_logic_vector(13348, 16),
18365 => conv_std_logic_vector(13419, 16),
18366 => conv_std_logic_vector(13490, 16),
18367 => conv_std_logic_vector(13561, 16),
18368 => conv_std_logic_vector(13632, 16),
18369 => conv_std_logic_vector(13703, 16),
18370 => conv_std_logic_vector(13774, 16),
18371 => conv_std_logic_vector(13845, 16),
18372 => conv_std_logic_vector(13916, 16),
18373 => conv_std_logic_vector(13987, 16),
18374 => conv_std_logic_vector(14058, 16),
18375 => conv_std_logic_vector(14129, 16),
18376 => conv_std_logic_vector(14200, 16),
18377 => conv_std_logic_vector(14271, 16),
18378 => conv_std_logic_vector(14342, 16),
18379 => conv_std_logic_vector(14413, 16),
18380 => conv_std_logic_vector(14484, 16),
18381 => conv_std_logic_vector(14555, 16),
18382 => conv_std_logic_vector(14626, 16),
18383 => conv_std_logic_vector(14697, 16),
18384 => conv_std_logic_vector(14768, 16),
18385 => conv_std_logic_vector(14839, 16),
18386 => conv_std_logic_vector(14910, 16),
18387 => conv_std_logic_vector(14981, 16),
18388 => conv_std_logic_vector(15052, 16),
18389 => conv_std_logic_vector(15123, 16),
18390 => conv_std_logic_vector(15194, 16),
18391 => conv_std_logic_vector(15265, 16),
18392 => conv_std_logic_vector(15336, 16),
18393 => conv_std_logic_vector(15407, 16),
18394 => conv_std_logic_vector(15478, 16),
18395 => conv_std_logic_vector(15549, 16),
18396 => conv_std_logic_vector(15620, 16),
18397 => conv_std_logic_vector(15691, 16),
18398 => conv_std_logic_vector(15762, 16),
18399 => conv_std_logic_vector(15833, 16),
18400 => conv_std_logic_vector(15904, 16),
18401 => conv_std_logic_vector(15975, 16),
18402 => conv_std_logic_vector(16046, 16),
18403 => conv_std_logic_vector(16117, 16),
18404 => conv_std_logic_vector(16188, 16),
18405 => conv_std_logic_vector(16259, 16),
18406 => conv_std_logic_vector(16330, 16),
18407 => conv_std_logic_vector(16401, 16),
18408 => conv_std_logic_vector(16472, 16),
18409 => conv_std_logic_vector(16543, 16),
18410 => conv_std_logic_vector(16614, 16),
18411 => conv_std_logic_vector(16685, 16),
18412 => conv_std_logic_vector(16756, 16),
18413 => conv_std_logic_vector(16827, 16),
18414 => conv_std_logic_vector(16898, 16),
18415 => conv_std_logic_vector(16969, 16),
18416 => conv_std_logic_vector(17040, 16),
18417 => conv_std_logic_vector(17111, 16),
18418 => conv_std_logic_vector(17182, 16),
18419 => conv_std_logic_vector(17253, 16),
18420 => conv_std_logic_vector(17324, 16),
18421 => conv_std_logic_vector(17395, 16),
18422 => conv_std_logic_vector(17466, 16),
18423 => conv_std_logic_vector(17537, 16),
18424 => conv_std_logic_vector(17608, 16),
18425 => conv_std_logic_vector(17679, 16),
18426 => conv_std_logic_vector(17750, 16),
18427 => conv_std_logic_vector(17821, 16),
18428 => conv_std_logic_vector(17892, 16),
18429 => conv_std_logic_vector(17963, 16),
18430 => conv_std_logic_vector(18034, 16),
18431 => conv_std_logic_vector(18105, 16),
18432 => conv_std_logic_vector(0, 16),
18433 => conv_std_logic_vector(72, 16),
18434 => conv_std_logic_vector(144, 16),
18435 => conv_std_logic_vector(216, 16),
18436 => conv_std_logic_vector(288, 16),
18437 => conv_std_logic_vector(360, 16),
18438 => conv_std_logic_vector(432, 16),
18439 => conv_std_logic_vector(504, 16),
18440 => conv_std_logic_vector(576, 16),
18441 => conv_std_logic_vector(648, 16),
18442 => conv_std_logic_vector(720, 16),
18443 => conv_std_logic_vector(792, 16),
18444 => conv_std_logic_vector(864, 16),
18445 => conv_std_logic_vector(936, 16),
18446 => conv_std_logic_vector(1008, 16),
18447 => conv_std_logic_vector(1080, 16),
18448 => conv_std_logic_vector(1152, 16),
18449 => conv_std_logic_vector(1224, 16),
18450 => conv_std_logic_vector(1296, 16),
18451 => conv_std_logic_vector(1368, 16),
18452 => conv_std_logic_vector(1440, 16),
18453 => conv_std_logic_vector(1512, 16),
18454 => conv_std_logic_vector(1584, 16),
18455 => conv_std_logic_vector(1656, 16),
18456 => conv_std_logic_vector(1728, 16),
18457 => conv_std_logic_vector(1800, 16),
18458 => conv_std_logic_vector(1872, 16),
18459 => conv_std_logic_vector(1944, 16),
18460 => conv_std_logic_vector(2016, 16),
18461 => conv_std_logic_vector(2088, 16),
18462 => conv_std_logic_vector(2160, 16),
18463 => conv_std_logic_vector(2232, 16),
18464 => conv_std_logic_vector(2304, 16),
18465 => conv_std_logic_vector(2376, 16),
18466 => conv_std_logic_vector(2448, 16),
18467 => conv_std_logic_vector(2520, 16),
18468 => conv_std_logic_vector(2592, 16),
18469 => conv_std_logic_vector(2664, 16),
18470 => conv_std_logic_vector(2736, 16),
18471 => conv_std_logic_vector(2808, 16),
18472 => conv_std_logic_vector(2880, 16),
18473 => conv_std_logic_vector(2952, 16),
18474 => conv_std_logic_vector(3024, 16),
18475 => conv_std_logic_vector(3096, 16),
18476 => conv_std_logic_vector(3168, 16),
18477 => conv_std_logic_vector(3240, 16),
18478 => conv_std_logic_vector(3312, 16),
18479 => conv_std_logic_vector(3384, 16),
18480 => conv_std_logic_vector(3456, 16),
18481 => conv_std_logic_vector(3528, 16),
18482 => conv_std_logic_vector(3600, 16),
18483 => conv_std_logic_vector(3672, 16),
18484 => conv_std_logic_vector(3744, 16),
18485 => conv_std_logic_vector(3816, 16),
18486 => conv_std_logic_vector(3888, 16),
18487 => conv_std_logic_vector(3960, 16),
18488 => conv_std_logic_vector(4032, 16),
18489 => conv_std_logic_vector(4104, 16),
18490 => conv_std_logic_vector(4176, 16),
18491 => conv_std_logic_vector(4248, 16),
18492 => conv_std_logic_vector(4320, 16),
18493 => conv_std_logic_vector(4392, 16),
18494 => conv_std_logic_vector(4464, 16),
18495 => conv_std_logic_vector(4536, 16),
18496 => conv_std_logic_vector(4608, 16),
18497 => conv_std_logic_vector(4680, 16),
18498 => conv_std_logic_vector(4752, 16),
18499 => conv_std_logic_vector(4824, 16),
18500 => conv_std_logic_vector(4896, 16),
18501 => conv_std_logic_vector(4968, 16),
18502 => conv_std_logic_vector(5040, 16),
18503 => conv_std_logic_vector(5112, 16),
18504 => conv_std_logic_vector(5184, 16),
18505 => conv_std_logic_vector(5256, 16),
18506 => conv_std_logic_vector(5328, 16),
18507 => conv_std_logic_vector(5400, 16),
18508 => conv_std_logic_vector(5472, 16),
18509 => conv_std_logic_vector(5544, 16),
18510 => conv_std_logic_vector(5616, 16),
18511 => conv_std_logic_vector(5688, 16),
18512 => conv_std_logic_vector(5760, 16),
18513 => conv_std_logic_vector(5832, 16),
18514 => conv_std_logic_vector(5904, 16),
18515 => conv_std_logic_vector(5976, 16),
18516 => conv_std_logic_vector(6048, 16),
18517 => conv_std_logic_vector(6120, 16),
18518 => conv_std_logic_vector(6192, 16),
18519 => conv_std_logic_vector(6264, 16),
18520 => conv_std_logic_vector(6336, 16),
18521 => conv_std_logic_vector(6408, 16),
18522 => conv_std_logic_vector(6480, 16),
18523 => conv_std_logic_vector(6552, 16),
18524 => conv_std_logic_vector(6624, 16),
18525 => conv_std_logic_vector(6696, 16),
18526 => conv_std_logic_vector(6768, 16),
18527 => conv_std_logic_vector(6840, 16),
18528 => conv_std_logic_vector(6912, 16),
18529 => conv_std_logic_vector(6984, 16),
18530 => conv_std_logic_vector(7056, 16),
18531 => conv_std_logic_vector(7128, 16),
18532 => conv_std_logic_vector(7200, 16),
18533 => conv_std_logic_vector(7272, 16),
18534 => conv_std_logic_vector(7344, 16),
18535 => conv_std_logic_vector(7416, 16),
18536 => conv_std_logic_vector(7488, 16),
18537 => conv_std_logic_vector(7560, 16),
18538 => conv_std_logic_vector(7632, 16),
18539 => conv_std_logic_vector(7704, 16),
18540 => conv_std_logic_vector(7776, 16),
18541 => conv_std_logic_vector(7848, 16),
18542 => conv_std_logic_vector(7920, 16),
18543 => conv_std_logic_vector(7992, 16),
18544 => conv_std_logic_vector(8064, 16),
18545 => conv_std_logic_vector(8136, 16),
18546 => conv_std_logic_vector(8208, 16),
18547 => conv_std_logic_vector(8280, 16),
18548 => conv_std_logic_vector(8352, 16),
18549 => conv_std_logic_vector(8424, 16),
18550 => conv_std_logic_vector(8496, 16),
18551 => conv_std_logic_vector(8568, 16),
18552 => conv_std_logic_vector(8640, 16),
18553 => conv_std_logic_vector(8712, 16),
18554 => conv_std_logic_vector(8784, 16),
18555 => conv_std_logic_vector(8856, 16),
18556 => conv_std_logic_vector(8928, 16),
18557 => conv_std_logic_vector(9000, 16),
18558 => conv_std_logic_vector(9072, 16),
18559 => conv_std_logic_vector(9144, 16),
18560 => conv_std_logic_vector(9216, 16),
18561 => conv_std_logic_vector(9288, 16),
18562 => conv_std_logic_vector(9360, 16),
18563 => conv_std_logic_vector(9432, 16),
18564 => conv_std_logic_vector(9504, 16),
18565 => conv_std_logic_vector(9576, 16),
18566 => conv_std_logic_vector(9648, 16),
18567 => conv_std_logic_vector(9720, 16),
18568 => conv_std_logic_vector(9792, 16),
18569 => conv_std_logic_vector(9864, 16),
18570 => conv_std_logic_vector(9936, 16),
18571 => conv_std_logic_vector(10008, 16),
18572 => conv_std_logic_vector(10080, 16),
18573 => conv_std_logic_vector(10152, 16),
18574 => conv_std_logic_vector(10224, 16),
18575 => conv_std_logic_vector(10296, 16),
18576 => conv_std_logic_vector(10368, 16),
18577 => conv_std_logic_vector(10440, 16),
18578 => conv_std_logic_vector(10512, 16),
18579 => conv_std_logic_vector(10584, 16),
18580 => conv_std_logic_vector(10656, 16),
18581 => conv_std_logic_vector(10728, 16),
18582 => conv_std_logic_vector(10800, 16),
18583 => conv_std_logic_vector(10872, 16),
18584 => conv_std_logic_vector(10944, 16),
18585 => conv_std_logic_vector(11016, 16),
18586 => conv_std_logic_vector(11088, 16),
18587 => conv_std_logic_vector(11160, 16),
18588 => conv_std_logic_vector(11232, 16),
18589 => conv_std_logic_vector(11304, 16),
18590 => conv_std_logic_vector(11376, 16),
18591 => conv_std_logic_vector(11448, 16),
18592 => conv_std_logic_vector(11520, 16),
18593 => conv_std_logic_vector(11592, 16),
18594 => conv_std_logic_vector(11664, 16),
18595 => conv_std_logic_vector(11736, 16),
18596 => conv_std_logic_vector(11808, 16),
18597 => conv_std_logic_vector(11880, 16),
18598 => conv_std_logic_vector(11952, 16),
18599 => conv_std_logic_vector(12024, 16),
18600 => conv_std_logic_vector(12096, 16),
18601 => conv_std_logic_vector(12168, 16),
18602 => conv_std_logic_vector(12240, 16),
18603 => conv_std_logic_vector(12312, 16),
18604 => conv_std_logic_vector(12384, 16),
18605 => conv_std_logic_vector(12456, 16),
18606 => conv_std_logic_vector(12528, 16),
18607 => conv_std_logic_vector(12600, 16),
18608 => conv_std_logic_vector(12672, 16),
18609 => conv_std_logic_vector(12744, 16),
18610 => conv_std_logic_vector(12816, 16),
18611 => conv_std_logic_vector(12888, 16),
18612 => conv_std_logic_vector(12960, 16),
18613 => conv_std_logic_vector(13032, 16),
18614 => conv_std_logic_vector(13104, 16),
18615 => conv_std_logic_vector(13176, 16),
18616 => conv_std_logic_vector(13248, 16),
18617 => conv_std_logic_vector(13320, 16),
18618 => conv_std_logic_vector(13392, 16),
18619 => conv_std_logic_vector(13464, 16),
18620 => conv_std_logic_vector(13536, 16),
18621 => conv_std_logic_vector(13608, 16),
18622 => conv_std_logic_vector(13680, 16),
18623 => conv_std_logic_vector(13752, 16),
18624 => conv_std_logic_vector(13824, 16),
18625 => conv_std_logic_vector(13896, 16),
18626 => conv_std_logic_vector(13968, 16),
18627 => conv_std_logic_vector(14040, 16),
18628 => conv_std_logic_vector(14112, 16),
18629 => conv_std_logic_vector(14184, 16),
18630 => conv_std_logic_vector(14256, 16),
18631 => conv_std_logic_vector(14328, 16),
18632 => conv_std_logic_vector(14400, 16),
18633 => conv_std_logic_vector(14472, 16),
18634 => conv_std_logic_vector(14544, 16),
18635 => conv_std_logic_vector(14616, 16),
18636 => conv_std_logic_vector(14688, 16),
18637 => conv_std_logic_vector(14760, 16),
18638 => conv_std_logic_vector(14832, 16),
18639 => conv_std_logic_vector(14904, 16),
18640 => conv_std_logic_vector(14976, 16),
18641 => conv_std_logic_vector(15048, 16),
18642 => conv_std_logic_vector(15120, 16),
18643 => conv_std_logic_vector(15192, 16),
18644 => conv_std_logic_vector(15264, 16),
18645 => conv_std_logic_vector(15336, 16),
18646 => conv_std_logic_vector(15408, 16),
18647 => conv_std_logic_vector(15480, 16),
18648 => conv_std_logic_vector(15552, 16),
18649 => conv_std_logic_vector(15624, 16),
18650 => conv_std_logic_vector(15696, 16),
18651 => conv_std_logic_vector(15768, 16),
18652 => conv_std_logic_vector(15840, 16),
18653 => conv_std_logic_vector(15912, 16),
18654 => conv_std_logic_vector(15984, 16),
18655 => conv_std_logic_vector(16056, 16),
18656 => conv_std_logic_vector(16128, 16),
18657 => conv_std_logic_vector(16200, 16),
18658 => conv_std_logic_vector(16272, 16),
18659 => conv_std_logic_vector(16344, 16),
18660 => conv_std_logic_vector(16416, 16),
18661 => conv_std_logic_vector(16488, 16),
18662 => conv_std_logic_vector(16560, 16),
18663 => conv_std_logic_vector(16632, 16),
18664 => conv_std_logic_vector(16704, 16),
18665 => conv_std_logic_vector(16776, 16),
18666 => conv_std_logic_vector(16848, 16),
18667 => conv_std_logic_vector(16920, 16),
18668 => conv_std_logic_vector(16992, 16),
18669 => conv_std_logic_vector(17064, 16),
18670 => conv_std_logic_vector(17136, 16),
18671 => conv_std_logic_vector(17208, 16),
18672 => conv_std_logic_vector(17280, 16),
18673 => conv_std_logic_vector(17352, 16),
18674 => conv_std_logic_vector(17424, 16),
18675 => conv_std_logic_vector(17496, 16),
18676 => conv_std_logic_vector(17568, 16),
18677 => conv_std_logic_vector(17640, 16),
18678 => conv_std_logic_vector(17712, 16),
18679 => conv_std_logic_vector(17784, 16),
18680 => conv_std_logic_vector(17856, 16),
18681 => conv_std_logic_vector(17928, 16),
18682 => conv_std_logic_vector(18000, 16),
18683 => conv_std_logic_vector(18072, 16),
18684 => conv_std_logic_vector(18144, 16),
18685 => conv_std_logic_vector(18216, 16),
18686 => conv_std_logic_vector(18288, 16),
18687 => conv_std_logic_vector(18360, 16),
18688 => conv_std_logic_vector(0, 16),
18689 => conv_std_logic_vector(73, 16),
18690 => conv_std_logic_vector(146, 16),
18691 => conv_std_logic_vector(219, 16),
18692 => conv_std_logic_vector(292, 16),
18693 => conv_std_logic_vector(365, 16),
18694 => conv_std_logic_vector(438, 16),
18695 => conv_std_logic_vector(511, 16),
18696 => conv_std_logic_vector(584, 16),
18697 => conv_std_logic_vector(657, 16),
18698 => conv_std_logic_vector(730, 16),
18699 => conv_std_logic_vector(803, 16),
18700 => conv_std_logic_vector(876, 16),
18701 => conv_std_logic_vector(949, 16),
18702 => conv_std_logic_vector(1022, 16),
18703 => conv_std_logic_vector(1095, 16),
18704 => conv_std_logic_vector(1168, 16),
18705 => conv_std_logic_vector(1241, 16),
18706 => conv_std_logic_vector(1314, 16),
18707 => conv_std_logic_vector(1387, 16),
18708 => conv_std_logic_vector(1460, 16),
18709 => conv_std_logic_vector(1533, 16),
18710 => conv_std_logic_vector(1606, 16),
18711 => conv_std_logic_vector(1679, 16),
18712 => conv_std_logic_vector(1752, 16),
18713 => conv_std_logic_vector(1825, 16),
18714 => conv_std_logic_vector(1898, 16),
18715 => conv_std_logic_vector(1971, 16),
18716 => conv_std_logic_vector(2044, 16),
18717 => conv_std_logic_vector(2117, 16),
18718 => conv_std_logic_vector(2190, 16),
18719 => conv_std_logic_vector(2263, 16),
18720 => conv_std_logic_vector(2336, 16),
18721 => conv_std_logic_vector(2409, 16),
18722 => conv_std_logic_vector(2482, 16),
18723 => conv_std_logic_vector(2555, 16),
18724 => conv_std_logic_vector(2628, 16),
18725 => conv_std_logic_vector(2701, 16),
18726 => conv_std_logic_vector(2774, 16),
18727 => conv_std_logic_vector(2847, 16),
18728 => conv_std_logic_vector(2920, 16),
18729 => conv_std_logic_vector(2993, 16),
18730 => conv_std_logic_vector(3066, 16),
18731 => conv_std_logic_vector(3139, 16),
18732 => conv_std_logic_vector(3212, 16),
18733 => conv_std_logic_vector(3285, 16),
18734 => conv_std_logic_vector(3358, 16),
18735 => conv_std_logic_vector(3431, 16),
18736 => conv_std_logic_vector(3504, 16),
18737 => conv_std_logic_vector(3577, 16),
18738 => conv_std_logic_vector(3650, 16),
18739 => conv_std_logic_vector(3723, 16),
18740 => conv_std_logic_vector(3796, 16),
18741 => conv_std_logic_vector(3869, 16),
18742 => conv_std_logic_vector(3942, 16),
18743 => conv_std_logic_vector(4015, 16),
18744 => conv_std_logic_vector(4088, 16),
18745 => conv_std_logic_vector(4161, 16),
18746 => conv_std_logic_vector(4234, 16),
18747 => conv_std_logic_vector(4307, 16),
18748 => conv_std_logic_vector(4380, 16),
18749 => conv_std_logic_vector(4453, 16),
18750 => conv_std_logic_vector(4526, 16),
18751 => conv_std_logic_vector(4599, 16),
18752 => conv_std_logic_vector(4672, 16),
18753 => conv_std_logic_vector(4745, 16),
18754 => conv_std_logic_vector(4818, 16),
18755 => conv_std_logic_vector(4891, 16),
18756 => conv_std_logic_vector(4964, 16),
18757 => conv_std_logic_vector(5037, 16),
18758 => conv_std_logic_vector(5110, 16),
18759 => conv_std_logic_vector(5183, 16),
18760 => conv_std_logic_vector(5256, 16),
18761 => conv_std_logic_vector(5329, 16),
18762 => conv_std_logic_vector(5402, 16),
18763 => conv_std_logic_vector(5475, 16),
18764 => conv_std_logic_vector(5548, 16),
18765 => conv_std_logic_vector(5621, 16),
18766 => conv_std_logic_vector(5694, 16),
18767 => conv_std_logic_vector(5767, 16),
18768 => conv_std_logic_vector(5840, 16),
18769 => conv_std_logic_vector(5913, 16),
18770 => conv_std_logic_vector(5986, 16),
18771 => conv_std_logic_vector(6059, 16),
18772 => conv_std_logic_vector(6132, 16),
18773 => conv_std_logic_vector(6205, 16),
18774 => conv_std_logic_vector(6278, 16),
18775 => conv_std_logic_vector(6351, 16),
18776 => conv_std_logic_vector(6424, 16),
18777 => conv_std_logic_vector(6497, 16),
18778 => conv_std_logic_vector(6570, 16),
18779 => conv_std_logic_vector(6643, 16),
18780 => conv_std_logic_vector(6716, 16),
18781 => conv_std_logic_vector(6789, 16),
18782 => conv_std_logic_vector(6862, 16),
18783 => conv_std_logic_vector(6935, 16),
18784 => conv_std_logic_vector(7008, 16),
18785 => conv_std_logic_vector(7081, 16),
18786 => conv_std_logic_vector(7154, 16),
18787 => conv_std_logic_vector(7227, 16),
18788 => conv_std_logic_vector(7300, 16),
18789 => conv_std_logic_vector(7373, 16),
18790 => conv_std_logic_vector(7446, 16),
18791 => conv_std_logic_vector(7519, 16),
18792 => conv_std_logic_vector(7592, 16),
18793 => conv_std_logic_vector(7665, 16),
18794 => conv_std_logic_vector(7738, 16),
18795 => conv_std_logic_vector(7811, 16),
18796 => conv_std_logic_vector(7884, 16),
18797 => conv_std_logic_vector(7957, 16),
18798 => conv_std_logic_vector(8030, 16),
18799 => conv_std_logic_vector(8103, 16),
18800 => conv_std_logic_vector(8176, 16),
18801 => conv_std_logic_vector(8249, 16),
18802 => conv_std_logic_vector(8322, 16),
18803 => conv_std_logic_vector(8395, 16),
18804 => conv_std_logic_vector(8468, 16),
18805 => conv_std_logic_vector(8541, 16),
18806 => conv_std_logic_vector(8614, 16),
18807 => conv_std_logic_vector(8687, 16),
18808 => conv_std_logic_vector(8760, 16),
18809 => conv_std_logic_vector(8833, 16),
18810 => conv_std_logic_vector(8906, 16),
18811 => conv_std_logic_vector(8979, 16),
18812 => conv_std_logic_vector(9052, 16),
18813 => conv_std_logic_vector(9125, 16),
18814 => conv_std_logic_vector(9198, 16),
18815 => conv_std_logic_vector(9271, 16),
18816 => conv_std_logic_vector(9344, 16),
18817 => conv_std_logic_vector(9417, 16),
18818 => conv_std_logic_vector(9490, 16),
18819 => conv_std_logic_vector(9563, 16),
18820 => conv_std_logic_vector(9636, 16),
18821 => conv_std_logic_vector(9709, 16),
18822 => conv_std_logic_vector(9782, 16),
18823 => conv_std_logic_vector(9855, 16),
18824 => conv_std_logic_vector(9928, 16),
18825 => conv_std_logic_vector(10001, 16),
18826 => conv_std_logic_vector(10074, 16),
18827 => conv_std_logic_vector(10147, 16),
18828 => conv_std_logic_vector(10220, 16),
18829 => conv_std_logic_vector(10293, 16),
18830 => conv_std_logic_vector(10366, 16),
18831 => conv_std_logic_vector(10439, 16),
18832 => conv_std_logic_vector(10512, 16),
18833 => conv_std_logic_vector(10585, 16),
18834 => conv_std_logic_vector(10658, 16),
18835 => conv_std_logic_vector(10731, 16),
18836 => conv_std_logic_vector(10804, 16),
18837 => conv_std_logic_vector(10877, 16),
18838 => conv_std_logic_vector(10950, 16),
18839 => conv_std_logic_vector(11023, 16),
18840 => conv_std_logic_vector(11096, 16),
18841 => conv_std_logic_vector(11169, 16),
18842 => conv_std_logic_vector(11242, 16),
18843 => conv_std_logic_vector(11315, 16),
18844 => conv_std_logic_vector(11388, 16),
18845 => conv_std_logic_vector(11461, 16),
18846 => conv_std_logic_vector(11534, 16),
18847 => conv_std_logic_vector(11607, 16),
18848 => conv_std_logic_vector(11680, 16),
18849 => conv_std_logic_vector(11753, 16),
18850 => conv_std_logic_vector(11826, 16),
18851 => conv_std_logic_vector(11899, 16),
18852 => conv_std_logic_vector(11972, 16),
18853 => conv_std_logic_vector(12045, 16),
18854 => conv_std_logic_vector(12118, 16),
18855 => conv_std_logic_vector(12191, 16),
18856 => conv_std_logic_vector(12264, 16),
18857 => conv_std_logic_vector(12337, 16),
18858 => conv_std_logic_vector(12410, 16),
18859 => conv_std_logic_vector(12483, 16),
18860 => conv_std_logic_vector(12556, 16),
18861 => conv_std_logic_vector(12629, 16),
18862 => conv_std_logic_vector(12702, 16),
18863 => conv_std_logic_vector(12775, 16),
18864 => conv_std_logic_vector(12848, 16),
18865 => conv_std_logic_vector(12921, 16),
18866 => conv_std_logic_vector(12994, 16),
18867 => conv_std_logic_vector(13067, 16),
18868 => conv_std_logic_vector(13140, 16),
18869 => conv_std_logic_vector(13213, 16),
18870 => conv_std_logic_vector(13286, 16),
18871 => conv_std_logic_vector(13359, 16),
18872 => conv_std_logic_vector(13432, 16),
18873 => conv_std_logic_vector(13505, 16),
18874 => conv_std_logic_vector(13578, 16),
18875 => conv_std_logic_vector(13651, 16),
18876 => conv_std_logic_vector(13724, 16),
18877 => conv_std_logic_vector(13797, 16),
18878 => conv_std_logic_vector(13870, 16),
18879 => conv_std_logic_vector(13943, 16),
18880 => conv_std_logic_vector(14016, 16),
18881 => conv_std_logic_vector(14089, 16),
18882 => conv_std_logic_vector(14162, 16),
18883 => conv_std_logic_vector(14235, 16),
18884 => conv_std_logic_vector(14308, 16),
18885 => conv_std_logic_vector(14381, 16),
18886 => conv_std_logic_vector(14454, 16),
18887 => conv_std_logic_vector(14527, 16),
18888 => conv_std_logic_vector(14600, 16),
18889 => conv_std_logic_vector(14673, 16),
18890 => conv_std_logic_vector(14746, 16),
18891 => conv_std_logic_vector(14819, 16),
18892 => conv_std_logic_vector(14892, 16),
18893 => conv_std_logic_vector(14965, 16),
18894 => conv_std_logic_vector(15038, 16),
18895 => conv_std_logic_vector(15111, 16),
18896 => conv_std_logic_vector(15184, 16),
18897 => conv_std_logic_vector(15257, 16),
18898 => conv_std_logic_vector(15330, 16),
18899 => conv_std_logic_vector(15403, 16),
18900 => conv_std_logic_vector(15476, 16),
18901 => conv_std_logic_vector(15549, 16),
18902 => conv_std_logic_vector(15622, 16),
18903 => conv_std_logic_vector(15695, 16),
18904 => conv_std_logic_vector(15768, 16),
18905 => conv_std_logic_vector(15841, 16),
18906 => conv_std_logic_vector(15914, 16),
18907 => conv_std_logic_vector(15987, 16),
18908 => conv_std_logic_vector(16060, 16),
18909 => conv_std_logic_vector(16133, 16),
18910 => conv_std_logic_vector(16206, 16),
18911 => conv_std_logic_vector(16279, 16),
18912 => conv_std_logic_vector(16352, 16),
18913 => conv_std_logic_vector(16425, 16),
18914 => conv_std_logic_vector(16498, 16),
18915 => conv_std_logic_vector(16571, 16),
18916 => conv_std_logic_vector(16644, 16),
18917 => conv_std_logic_vector(16717, 16),
18918 => conv_std_logic_vector(16790, 16),
18919 => conv_std_logic_vector(16863, 16),
18920 => conv_std_logic_vector(16936, 16),
18921 => conv_std_logic_vector(17009, 16),
18922 => conv_std_logic_vector(17082, 16),
18923 => conv_std_logic_vector(17155, 16),
18924 => conv_std_logic_vector(17228, 16),
18925 => conv_std_logic_vector(17301, 16),
18926 => conv_std_logic_vector(17374, 16),
18927 => conv_std_logic_vector(17447, 16),
18928 => conv_std_logic_vector(17520, 16),
18929 => conv_std_logic_vector(17593, 16),
18930 => conv_std_logic_vector(17666, 16),
18931 => conv_std_logic_vector(17739, 16),
18932 => conv_std_logic_vector(17812, 16),
18933 => conv_std_logic_vector(17885, 16),
18934 => conv_std_logic_vector(17958, 16),
18935 => conv_std_logic_vector(18031, 16),
18936 => conv_std_logic_vector(18104, 16),
18937 => conv_std_logic_vector(18177, 16),
18938 => conv_std_logic_vector(18250, 16),
18939 => conv_std_logic_vector(18323, 16),
18940 => conv_std_logic_vector(18396, 16),
18941 => conv_std_logic_vector(18469, 16),
18942 => conv_std_logic_vector(18542, 16),
18943 => conv_std_logic_vector(18615, 16),
18944 => conv_std_logic_vector(0, 16),
18945 => conv_std_logic_vector(74, 16),
18946 => conv_std_logic_vector(148, 16),
18947 => conv_std_logic_vector(222, 16),
18948 => conv_std_logic_vector(296, 16),
18949 => conv_std_logic_vector(370, 16),
18950 => conv_std_logic_vector(444, 16),
18951 => conv_std_logic_vector(518, 16),
18952 => conv_std_logic_vector(592, 16),
18953 => conv_std_logic_vector(666, 16),
18954 => conv_std_logic_vector(740, 16),
18955 => conv_std_logic_vector(814, 16),
18956 => conv_std_logic_vector(888, 16),
18957 => conv_std_logic_vector(962, 16),
18958 => conv_std_logic_vector(1036, 16),
18959 => conv_std_logic_vector(1110, 16),
18960 => conv_std_logic_vector(1184, 16),
18961 => conv_std_logic_vector(1258, 16),
18962 => conv_std_logic_vector(1332, 16),
18963 => conv_std_logic_vector(1406, 16),
18964 => conv_std_logic_vector(1480, 16),
18965 => conv_std_logic_vector(1554, 16),
18966 => conv_std_logic_vector(1628, 16),
18967 => conv_std_logic_vector(1702, 16),
18968 => conv_std_logic_vector(1776, 16),
18969 => conv_std_logic_vector(1850, 16),
18970 => conv_std_logic_vector(1924, 16),
18971 => conv_std_logic_vector(1998, 16),
18972 => conv_std_logic_vector(2072, 16),
18973 => conv_std_logic_vector(2146, 16),
18974 => conv_std_logic_vector(2220, 16),
18975 => conv_std_logic_vector(2294, 16),
18976 => conv_std_logic_vector(2368, 16),
18977 => conv_std_logic_vector(2442, 16),
18978 => conv_std_logic_vector(2516, 16),
18979 => conv_std_logic_vector(2590, 16),
18980 => conv_std_logic_vector(2664, 16),
18981 => conv_std_logic_vector(2738, 16),
18982 => conv_std_logic_vector(2812, 16),
18983 => conv_std_logic_vector(2886, 16),
18984 => conv_std_logic_vector(2960, 16),
18985 => conv_std_logic_vector(3034, 16),
18986 => conv_std_logic_vector(3108, 16),
18987 => conv_std_logic_vector(3182, 16),
18988 => conv_std_logic_vector(3256, 16),
18989 => conv_std_logic_vector(3330, 16),
18990 => conv_std_logic_vector(3404, 16),
18991 => conv_std_logic_vector(3478, 16),
18992 => conv_std_logic_vector(3552, 16),
18993 => conv_std_logic_vector(3626, 16),
18994 => conv_std_logic_vector(3700, 16),
18995 => conv_std_logic_vector(3774, 16),
18996 => conv_std_logic_vector(3848, 16),
18997 => conv_std_logic_vector(3922, 16),
18998 => conv_std_logic_vector(3996, 16),
18999 => conv_std_logic_vector(4070, 16),
19000 => conv_std_logic_vector(4144, 16),
19001 => conv_std_logic_vector(4218, 16),
19002 => conv_std_logic_vector(4292, 16),
19003 => conv_std_logic_vector(4366, 16),
19004 => conv_std_logic_vector(4440, 16),
19005 => conv_std_logic_vector(4514, 16),
19006 => conv_std_logic_vector(4588, 16),
19007 => conv_std_logic_vector(4662, 16),
19008 => conv_std_logic_vector(4736, 16),
19009 => conv_std_logic_vector(4810, 16),
19010 => conv_std_logic_vector(4884, 16),
19011 => conv_std_logic_vector(4958, 16),
19012 => conv_std_logic_vector(5032, 16),
19013 => conv_std_logic_vector(5106, 16),
19014 => conv_std_logic_vector(5180, 16),
19015 => conv_std_logic_vector(5254, 16),
19016 => conv_std_logic_vector(5328, 16),
19017 => conv_std_logic_vector(5402, 16),
19018 => conv_std_logic_vector(5476, 16),
19019 => conv_std_logic_vector(5550, 16),
19020 => conv_std_logic_vector(5624, 16),
19021 => conv_std_logic_vector(5698, 16),
19022 => conv_std_logic_vector(5772, 16),
19023 => conv_std_logic_vector(5846, 16),
19024 => conv_std_logic_vector(5920, 16),
19025 => conv_std_logic_vector(5994, 16),
19026 => conv_std_logic_vector(6068, 16),
19027 => conv_std_logic_vector(6142, 16),
19028 => conv_std_logic_vector(6216, 16),
19029 => conv_std_logic_vector(6290, 16),
19030 => conv_std_logic_vector(6364, 16),
19031 => conv_std_logic_vector(6438, 16),
19032 => conv_std_logic_vector(6512, 16),
19033 => conv_std_logic_vector(6586, 16),
19034 => conv_std_logic_vector(6660, 16),
19035 => conv_std_logic_vector(6734, 16),
19036 => conv_std_logic_vector(6808, 16),
19037 => conv_std_logic_vector(6882, 16),
19038 => conv_std_logic_vector(6956, 16),
19039 => conv_std_logic_vector(7030, 16),
19040 => conv_std_logic_vector(7104, 16),
19041 => conv_std_logic_vector(7178, 16),
19042 => conv_std_logic_vector(7252, 16),
19043 => conv_std_logic_vector(7326, 16),
19044 => conv_std_logic_vector(7400, 16),
19045 => conv_std_logic_vector(7474, 16),
19046 => conv_std_logic_vector(7548, 16),
19047 => conv_std_logic_vector(7622, 16),
19048 => conv_std_logic_vector(7696, 16),
19049 => conv_std_logic_vector(7770, 16),
19050 => conv_std_logic_vector(7844, 16),
19051 => conv_std_logic_vector(7918, 16),
19052 => conv_std_logic_vector(7992, 16),
19053 => conv_std_logic_vector(8066, 16),
19054 => conv_std_logic_vector(8140, 16),
19055 => conv_std_logic_vector(8214, 16),
19056 => conv_std_logic_vector(8288, 16),
19057 => conv_std_logic_vector(8362, 16),
19058 => conv_std_logic_vector(8436, 16),
19059 => conv_std_logic_vector(8510, 16),
19060 => conv_std_logic_vector(8584, 16),
19061 => conv_std_logic_vector(8658, 16),
19062 => conv_std_logic_vector(8732, 16),
19063 => conv_std_logic_vector(8806, 16),
19064 => conv_std_logic_vector(8880, 16),
19065 => conv_std_logic_vector(8954, 16),
19066 => conv_std_logic_vector(9028, 16),
19067 => conv_std_logic_vector(9102, 16),
19068 => conv_std_logic_vector(9176, 16),
19069 => conv_std_logic_vector(9250, 16),
19070 => conv_std_logic_vector(9324, 16),
19071 => conv_std_logic_vector(9398, 16),
19072 => conv_std_logic_vector(9472, 16),
19073 => conv_std_logic_vector(9546, 16),
19074 => conv_std_logic_vector(9620, 16),
19075 => conv_std_logic_vector(9694, 16),
19076 => conv_std_logic_vector(9768, 16),
19077 => conv_std_logic_vector(9842, 16),
19078 => conv_std_logic_vector(9916, 16),
19079 => conv_std_logic_vector(9990, 16),
19080 => conv_std_logic_vector(10064, 16),
19081 => conv_std_logic_vector(10138, 16),
19082 => conv_std_logic_vector(10212, 16),
19083 => conv_std_logic_vector(10286, 16),
19084 => conv_std_logic_vector(10360, 16),
19085 => conv_std_logic_vector(10434, 16),
19086 => conv_std_logic_vector(10508, 16),
19087 => conv_std_logic_vector(10582, 16),
19088 => conv_std_logic_vector(10656, 16),
19089 => conv_std_logic_vector(10730, 16),
19090 => conv_std_logic_vector(10804, 16),
19091 => conv_std_logic_vector(10878, 16),
19092 => conv_std_logic_vector(10952, 16),
19093 => conv_std_logic_vector(11026, 16),
19094 => conv_std_logic_vector(11100, 16),
19095 => conv_std_logic_vector(11174, 16),
19096 => conv_std_logic_vector(11248, 16),
19097 => conv_std_logic_vector(11322, 16),
19098 => conv_std_logic_vector(11396, 16),
19099 => conv_std_logic_vector(11470, 16),
19100 => conv_std_logic_vector(11544, 16),
19101 => conv_std_logic_vector(11618, 16),
19102 => conv_std_logic_vector(11692, 16),
19103 => conv_std_logic_vector(11766, 16),
19104 => conv_std_logic_vector(11840, 16),
19105 => conv_std_logic_vector(11914, 16),
19106 => conv_std_logic_vector(11988, 16),
19107 => conv_std_logic_vector(12062, 16),
19108 => conv_std_logic_vector(12136, 16),
19109 => conv_std_logic_vector(12210, 16),
19110 => conv_std_logic_vector(12284, 16),
19111 => conv_std_logic_vector(12358, 16),
19112 => conv_std_logic_vector(12432, 16),
19113 => conv_std_logic_vector(12506, 16),
19114 => conv_std_logic_vector(12580, 16),
19115 => conv_std_logic_vector(12654, 16),
19116 => conv_std_logic_vector(12728, 16),
19117 => conv_std_logic_vector(12802, 16),
19118 => conv_std_logic_vector(12876, 16),
19119 => conv_std_logic_vector(12950, 16),
19120 => conv_std_logic_vector(13024, 16),
19121 => conv_std_logic_vector(13098, 16),
19122 => conv_std_logic_vector(13172, 16),
19123 => conv_std_logic_vector(13246, 16),
19124 => conv_std_logic_vector(13320, 16),
19125 => conv_std_logic_vector(13394, 16),
19126 => conv_std_logic_vector(13468, 16),
19127 => conv_std_logic_vector(13542, 16),
19128 => conv_std_logic_vector(13616, 16),
19129 => conv_std_logic_vector(13690, 16),
19130 => conv_std_logic_vector(13764, 16),
19131 => conv_std_logic_vector(13838, 16),
19132 => conv_std_logic_vector(13912, 16),
19133 => conv_std_logic_vector(13986, 16),
19134 => conv_std_logic_vector(14060, 16),
19135 => conv_std_logic_vector(14134, 16),
19136 => conv_std_logic_vector(14208, 16),
19137 => conv_std_logic_vector(14282, 16),
19138 => conv_std_logic_vector(14356, 16),
19139 => conv_std_logic_vector(14430, 16),
19140 => conv_std_logic_vector(14504, 16),
19141 => conv_std_logic_vector(14578, 16),
19142 => conv_std_logic_vector(14652, 16),
19143 => conv_std_logic_vector(14726, 16),
19144 => conv_std_logic_vector(14800, 16),
19145 => conv_std_logic_vector(14874, 16),
19146 => conv_std_logic_vector(14948, 16),
19147 => conv_std_logic_vector(15022, 16),
19148 => conv_std_logic_vector(15096, 16),
19149 => conv_std_logic_vector(15170, 16),
19150 => conv_std_logic_vector(15244, 16),
19151 => conv_std_logic_vector(15318, 16),
19152 => conv_std_logic_vector(15392, 16),
19153 => conv_std_logic_vector(15466, 16),
19154 => conv_std_logic_vector(15540, 16),
19155 => conv_std_logic_vector(15614, 16),
19156 => conv_std_logic_vector(15688, 16),
19157 => conv_std_logic_vector(15762, 16),
19158 => conv_std_logic_vector(15836, 16),
19159 => conv_std_logic_vector(15910, 16),
19160 => conv_std_logic_vector(15984, 16),
19161 => conv_std_logic_vector(16058, 16),
19162 => conv_std_logic_vector(16132, 16),
19163 => conv_std_logic_vector(16206, 16),
19164 => conv_std_logic_vector(16280, 16),
19165 => conv_std_logic_vector(16354, 16),
19166 => conv_std_logic_vector(16428, 16),
19167 => conv_std_logic_vector(16502, 16),
19168 => conv_std_logic_vector(16576, 16),
19169 => conv_std_logic_vector(16650, 16),
19170 => conv_std_logic_vector(16724, 16),
19171 => conv_std_logic_vector(16798, 16),
19172 => conv_std_logic_vector(16872, 16),
19173 => conv_std_logic_vector(16946, 16),
19174 => conv_std_logic_vector(17020, 16),
19175 => conv_std_logic_vector(17094, 16),
19176 => conv_std_logic_vector(17168, 16),
19177 => conv_std_logic_vector(17242, 16),
19178 => conv_std_logic_vector(17316, 16),
19179 => conv_std_logic_vector(17390, 16),
19180 => conv_std_logic_vector(17464, 16),
19181 => conv_std_logic_vector(17538, 16),
19182 => conv_std_logic_vector(17612, 16),
19183 => conv_std_logic_vector(17686, 16),
19184 => conv_std_logic_vector(17760, 16),
19185 => conv_std_logic_vector(17834, 16),
19186 => conv_std_logic_vector(17908, 16),
19187 => conv_std_logic_vector(17982, 16),
19188 => conv_std_logic_vector(18056, 16),
19189 => conv_std_logic_vector(18130, 16),
19190 => conv_std_logic_vector(18204, 16),
19191 => conv_std_logic_vector(18278, 16),
19192 => conv_std_logic_vector(18352, 16),
19193 => conv_std_logic_vector(18426, 16),
19194 => conv_std_logic_vector(18500, 16),
19195 => conv_std_logic_vector(18574, 16),
19196 => conv_std_logic_vector(18648, 16),
19197 => conv_std_logic_vector(18722, 16),
19198 => conv_std_logic_vector(18796, 16),
19199 => conv_std_logic_vector(18870, 16),
19200 => conv_std_logic_vector(0, 16),
19201 => conv_std_logic_vector(75, 16),
19202 => conv_std_logic_vector(150, 16),
19203 => conv_std_logic_vector(225, 16),
19204 => conv_std_logic_vector(300, 16),
19205 => conv_std_logic_vector(375, 16),
19206 => conv_std_logic_vector(450, 16),
19207 => conv_std_logic_vector(525, 16),
19208 => conv_std_logic_vector(600, 16),
19209 => conv_std_logic_vector(675, 16),
19210 => conv_std_logic_vector(750, 16),
19211 => conv_std_logic_vector(825, 16),
19212 => conv_std_logic_vector(900, 16),
19213 => conv_std_logic_vector(975, 16),
19214 => conv_std_logic_vector(1050, 16),
19215 => conv_std_logic_vector(1125, 16),
19216 => conv_std_logic_vector(1200, 16),
19217 => conv_std_logic_vector(1275, 16),
19218 => conv_std_logic_vector(1350, 16),
19219 => conv_std_logic_vector(1425, 16),
19220 => conv_std_logic_vector(1500, 16),
19221 => conv_std_logic_vector(1575, 16),
19222 => conv_std_logic_vector(1650, 16),
19223 => conv_std_logic_vector(1725, 16),
19224 => conv_std_logic_vector(1800, 16),
19225 => conv_std_logic_vector(1875, 16),
19226 => conv_std_logic_vector(1950, 16),
19227 => conv_std_logic_vector(2025, 16),
19228 => conv_std_logic_vector(2100, 16),
19229 => conv_std_logic_vector(2175, 16),
19230 => conv_std_logic_vector(2250, 16),
19231 => conv_std_logic_vector(2325, 16),
19232 => conv_std_logic_vector(2400, 16),
19233 => conv_std_logic_vector(2475, 16),
19234 => conv_std_logic_vector(2550, 16),
19235 => conv_std_logic_vector(2625, 16),
19236 => conv_std_logic_vector(2700, 16),
19237 => conv_std_logic_vector(2775, 16),
19238 => conv_std_logic_vector(2850, 16),
19239 => conv_std_logic_vector(2925, 16),
19240 => conv_std_logic_vector(3000, 16),
19241 => conv_std_logic_vector(3075, 16),
19242 => conv_std_logic_vector(3150, 16),
19243 => conv_std_logic_vector(3225, 16),
19244 => conv_std_logic_vector(3300, 16),
19245 => conv_std_logic_vector(3375, 16),
19246 => conv_std_logic_vector(3450, 16),
19247 => conv_std_logic_vector(3525, 16),
19248 => conv_std_logic_vector(3600, 16),
19249 => conv_std_logic_vector(3675, 16),
19250 => conv_std_logic_vector(3750, 16),
19251 => conv_std_logic_vector(3825, 16),
19252 => conv_std_logic_vector(3900, 16),
19253 => conv_std_logic_vector(3975, 16),
19254 => conv_std_logic_vector(4050, 16),
19255 => conv_std_logic_vector(4125, 16),
19256 => conv_std_logic_vector(4200, 16),
19257 => conv_std_logic_vector(4275, 16),
19258 => conv_std_logic_vector(4350, 16),
19259 => conv_std_logic_vector(4425, 16),
19260 => conv_std_logic_vector(4500, 16),
19261 => conv_std_logic_vector(4575, 16),
19262 => conv_std_logic_vector(4650, 16),
19263 => conv_std_logic_vector(4725, 16),
19264 => conv_std_logic_vector(4800, 16),
19265 => conv_std_logic_vector(4875, 16),
19266 => conv_std_logic_vector(4950, 16),
19267 => conv_std_logic_vector(5025, 16),
19268 => conv_std_logic_vector(5100, 16),
19269 => conv_std_logic_vector(5175, 16),
19270 => conv_std_logic_vector(5250, 16),
19271 => conv_std_logic_vector(5325, 16),
19272 => conv_std_logic_vector(5400, 16),
19273 => conv_std_logic_vector(5475, 16),
19274 => conv_std_logic_vector(5550, 16),
19275 => conv_std_logic_vector(5625, 16),
19276 => conv_std_logic_vector(5700, 16),
19277 => conv_std_logic_vector(5775, 16),
19278 => conv_std_logic_vector(5850, 16),
19279 => conv_std_logic_vector(5925, 16),
19280 => conv_std_logic_vector(6000, 16),
19281 => conv_std_logic_vector(6075, 16),
19282 => conv_std_logic_vector(6150, 16),
19283 => conv_std_logic_vector(6225, 16),
19284 => conv_std_logic_vector(6300, 16),
19285 => conv_std_logic_vector(6375, 16),
19286 => conv_std_logic_vector(6450, 16),
19287 => conv_std_logic_vector(6525, 16),
19288 => conv_std_logic_vector(6600, 16),
19289 => conv_std_logic_vector(6675, 16),
19290 => conv_std_logic_vector(6750, 16),
19291 => conv_std_logic_vector(6825, 16),
19292 => conv_std_logic_vector(6900, 16),
19293 => conv_std_logic_vector(6975, 16),
19294 => conv_std_logic_vector(7050, 16),
19295 => conv_std_logic_vector(7125, 16),
19296 => conv_std_logic_vector(7200, 16),
19297 => conv_std_logic_vector(7275, 16),
19298 => conv_std_logic_vector(7350, 16),
19299 => conv_std_logic_vector(7425, 16),
19300 => conv_std_logic_vector(7500, 16),
19301 => conv_std_logic_vector(7575, 16),
19302 => conv_std_logic_vector(7650, 16),
19303 => conv_std_logic_vector(7725, 16),
19304 => conv_std_logic_vector(7800, 16),
19305 => conv_std_logic_vector(7875, 16),
19306 => conv_std_logic_vector(7950, 16),
19307 => conv_std_logic_vector(8025, 16),
19308 => conv_std_logic_vector(8100, 16),
19309 => conv_std_logic_vector(8175, 16),
19310 => conv_std_logic_vector(8250, 16),
19311 => conv_std_logic_vector(8325, 16),
19312 => conv_std_logic_vector(8400, 16),
19313 => conv_std_logic_vector(8475, 16),
19314 => conv_std_logic_vector(8550, 16),
19315 => conv_std_logic_vector(8625, 16),
19316 => conv_std_logic_vector(8700, 16),
19317 => conv_std_logic_vector(8775, 16),
19318 => conv_std_logic_vector(8850, 16),
19319 => conv_std_logic_vector(8925, 16),
19320 => conv_std_logic_vector(9000, 16),
19321 => conv_std_logic_vector(9075, 16),
19322 => conv_std_logic_vector(9150, 16),
19323 => conv_std_logic_vector(9225, 16),
19324 => conv_std_logic_vector(9300, 16),
19325 => conv_std_logic_vector(9375, 16),
19326 => conv_std_logic_vector(9450, 16),
19327 => conv_std_logic_vector(9525, 16),
19328 => conv_std_logic_vector(9600, 16),
19329 => conv_std_logic_vector(9675, 16),
19330 => conv_std_logic_vector(9750, 16),
19331 => conv_std_logic_vector(9825, 16),
19332 => conv_std_logic_vector(9900, 16),
19333 => conv_std_logic_vector(9975, 16),
19334 => conv_std_logic_vector(10050, 16),
19335 => conv_std_logic_vector(10125, 16),
19336 => conv_std_logic_vector(10200, 16),
19337 => conv_std_logic_vector(10275, 16),
19338 => conv_std_logic_vector(10350, 16),
19339 => conv_std_logic_vector(10425, 16),
19340 => conv_std_logic_vector(10500, 16),
19341 => conv_std_logic_vector(10575, 16),
19342 => conv_std_logic_vector(10650, 16),
19343 => conv_std_logic_vector(10725, 16),
19344 => conv_std_logic_vector(10800, 16),
19345 => conv_std_logic_vector(10875, 16),
19346 => conv_std_logic_vector(10950, 16),
19347 => conv_std_logic_vector(11025, 16),
19348 => conv_std_logic_vector(11100, 16),
19349 => conv_std_logic_vector(11175, 16),
19350 => conv_std_logic_vector(11250, 16),
19351 => conv_std_logic_vector(11325, 16),
19352 => conv_std_logic_vector(11400, 16),
19353 => conv_std_logic_vector(11475, 16),
19354 => conv_std_logic_vector(11550, 16),
19355 => conv_std_logic_vector(11625, 16),
19356 => conv_std_logic_vector(11700, 16),
19357 => conv_std_logic_vector(11775, 16),
19358 => conv_std_logic_vector(11850, 16),
19359 => conv_std_logic_vector(11925, 16),
19360 => conv_std_logic_vector(12000, 16),
19361 => conv_std_logic_vector(12075, 16),
19362 => conv_std_logic_vector(12150, 16),
19363 => conv_std_logic_vector(12225, 16),
19364 => conv_std_logic_vector(12300, 16),
19365 => conv_std_logic_vector(12375, 16),
19366 => conv_std_logic_vector(12450, 16),
19367 => conv_std_logic_vector(12525, 16),
19368 => conv_std_logic_vector(12600, 16),
19369 => conv_std_logic_vector(12675, 16),
19370 => conv_std_logic_vector(12750, 16),
19371 => conv_std_logic_vector(12825, 16),
19372 => conv_std_logic_vector(12900, 16),
19373 => conv_std_logic_vector(12975, 16),
19374 => conv_std_logic_vector(13050, 16),
19375 => conv_std_logic_vector(13125, 16),
19376 => conv_std_logic_vector(13200, 16),
19377 => conv_std_logic_vector(13275, 16),
19378 => conv_std_logic_vector(13350, 16),
19379 => conv_std_logic_vector(13425, 16),
19380 => conv_std_logic_vector(13500, 16),
19381 => conv_std_logic_vector(13575, 16),
19382 => conv_std_logic_vector(13650, 16),
19383 => conv_std_logic_vector(13725, 16),
19384 => conv_std_logic_vector(13800, 16),
19385 => conv_std_logic_vector(13875, 16),
19386 => conv_std_logic_vector(13950, 16),
19387 => conv_std_logic_vector(14025, 16),
19388 => conv_std_logic_vector(14100, 16),
19389 => conv_std_logic_vector(14175, 16),
19390 => conv_std_logic_vector(14250, 16),
19391 => conv_std_logic_vector(14325, 16),
19392 => conv_std_logic_vector(14400, 16),
19393 => conv_std_logic_vector(14475, 16),
19394 => conv_std_logic_vector(14550, 16),
19395 => conv_std_logic_vector(14625, 16),
19396 => conv_std_logic_vector(14700, 16),
19397 => conv_std_logic_vector(14775, 16),
19398 => conv_std_logic_vector(14850, 16),
19399 => conv_std_logic_vector(14925, 16),
19400 => conv_std_logic_vector(15000, 16),
19401 => conv_std_logic_vector(15075, 16),
19402 => conv_std_logic_vector(15150, 16),
19403 => conv_std_logic_vector(15225, 16),
19404 => conv_std_logic_vector(15300, 16),
19405 => conv_std_logic_vector(15375, 16),
19406 => conv_std_logic_vector(15450, 16),
19407 => conv_std_logic_vector(15525, 16),
19408 => conv_std_logic_vector(15600, 16),
19409 => conv_std_logic_vector(15675, 16),
19410 => conv_std_logic_vector(15750, 16),
19411 => conv_std_logic_vector(15825, 16),
19412 => conv_std_logic_vector(15900, 16),
19413 => conv_std_logic_vector(15975, 16),
19414 => conv_std_logic_vector(16050, 16),
19415 => conv_std_logic_vector(16125, 16),
19416 => conv_std_logic_vector(16200, 16),
19417 => conv_std_logic_vector(16275, 16),
19418 => conv_std_logic_vector(16350, 16),
19419 => conv_std_logic_vector(16425, 16),
19420 => conv_std_logic_vector(16500, 16),
19421 => conv_std_logic_vector(16575, 16),
19422 => conv_std_logic_vector(16650, 16),
19423 => conv_std_logic_vector(16725, 16),
19424 => conv_std_logic_vector(16800, 16),
19425 => conv_std_logic_vector(16875, 16),
19426 => conv_std_logic_vector(16950, 16),
19427 => conv_std_logic_vector(17025, 16),
19428 => conv_std_logic_vector(17100, 16),
19429 => conv_std_logic_vector(17175, 16),
19430 => conv_std_logic_vector(17250, 16),
19431 => conv_std_logic_vector(17325, 16),
19432 => conv_std_logic_vector(17400, 16),
19433 => conv_std_logic_vector(17475, 16),
19434 => conv_std_logic_vector(17550, 16),
19435 => conv_std_logic_vector(17625, 16),
19436 => conv_std_logic_vector(17700, 16),
19437 => conv_std_logic_vector(17775, 16),
19438 => conv_std_logic_vector(17850, 16),
19439 => conv_std_logic_vector(17925, 16),
19440 => conv_std_logic_vector(18000, 16),
19441 => conv_std_logic_vector(18075, 16),
19442 => conv_std_logic_vector(18150, 16),
19443 => conv_std_logic_vector(18225, 16),
19444 => conv_std_logic_vector(18300, 16),
19445 => conv_std_logic_vector(18375, 16),
19446 => conv_std_logic_vector(18450, 16),
19447 => conv_std_logic_vector(18525, 16),
19448 => conv_std_logic_vector(18600, 16),
19449 => conv_std_logic_vector(18675, 16),
19450 => conv_std_logic_vector(18750, 16),
19451 => conv_std_logic_vector(18825, 16),
19452 => conv_std_logic_vector(18900, 16),
19453 => conv_std_logic_vector(18975, 16),
19454 => conv_std_logic_vector(19050, 16),
19455 => conv_std_logic_vector(19125, 16),
19456 => conv_std_logic_vector(0, 16),
19457 => conv_std_logic_vector(76, 16),
19458 => conv_std_logic_vector(152, 16),
19459 => conv_std_logic_vector(228, 16),
19460 => conv_std_logic_vector(304, 16),
19461 => conv_std_logic_vector(380, 16),
19462 => conv_std_logic_vector(456, 16),
19463 => conv_std_logic_vector(532, 16),
19464 => conv_std_logic_vector(608, 16),
19465 => conv_std_logic_vector(684, 16),
19466 => conv_std_logic_vector(760, 16),
19467 => conv_std_logic_vector(836, 16),
19468 => conv_std_logic_vector(912, 16),
19469 => conv_std_logic_vector(988, 16),
19470 => conv_std_logic_vector(1064, 16),
19471 => conv_std_logic_vector(1140, 16),
19472 => conv_std_logic_vector(1216, 16),
19473 => conv_std_logic_vector(1292, 16),
19474 => conv_std_logic_vector(1368, 16),
19475 => conv_std_logic_vector(1444, 16),
19476 => conv_std_logic_vector(1520, 16),
19477 => conv_std_logic_vector(1596, 16),
19478 => conv_std_logic_vector(1672, 16),
19479 => conv_std_logic_vector(1748, 16),
19480 => conv_std_logic_vector(1824, 16),
19481 => conv_std_logic_vector(1900, 16),
19482 => conv_std_logic_vector(1976, 16),
19483 => conv_std_logic_vector(2052, 16),
19484 => conv_std_logic_vector(2128, 16),
19485 => conv_std_logic_vector(2204, 16),
19486 => conv_std_logic_vector(2280, 16),
19487 => conv_std_logic_vector(2356, 16),
19488 => conv_std_logic_vector(2432, 16),
19489 => conv_std_logic_vector(2508, 16),
19490 => conv_std_logic_vector(2584, 16),
19491 => conv_std_logic_vector(2660, 16),
19492 => conv_std_logic_vector(2736, 16),
19493 => conv_std_logic_vector(2812, 16),
19494 => conv_std_logic_vector(2888, 16),
19495 => conv_std_logic_vector(2964, 16),
19496 => conv_std_logic_vector(3040, 16),
19497 => conv_std_logic_vector(3116, 16),
19498 => conv_std_logic_vector(3192, 16),
19499 => conv_std_logic_vector(3268, 16),
19500 => conv_std_logic_vector(3344, 16),
19501 => conv_std_logic_vector(3420, 16),
19502 => conv_std_logic_vector(3496, 16),
19503 => conv_std_logic_vector(3572, 16),
19504 => conv_std_logic_vector(3648, 16),
19505 => conv_std_logic_vector(3724, 16),
19506 => conv_std_logic_vector(3800, 16),
19507 => conv_std_logic_vector(3876, 16),
19508 => conv_std_logic_vector(3952, 16),
19509 => conv_std_logic_vector(4028, 16),
19510 => conv_std_logic_vector(4104, 16),
19511 => conv_std_logic_vector(4180, 16),
19512 => conv_std_logic_vector(4256, 16),
19513 => conv_std_logic_vector(4332, 16),
19514 => conv_std_logic_vector(4408, 16),
19515 => conv_std_logic_vector(4484, 16),
19516 => conv_std_logic_vector(4560, 16),
19517 => conv_std_logic_vector(4636, 16),
19518 => conv_std_logic_vector(4712, 16),
19519 => conv_std_logic_vector(4788, 16),
19520 => conv_std_logic_vector(4864, 16),
19521 => conv_std_logic_vector(4940, 16),
19522 => conv_std_logic_vector(5016, 16),
19523 => conv_std_logic_vector(5092, 16),
19524 => conv_std_logic_vector(5168, 16),
19525 => conv_std_logic_vector(5244, 16),
19526 => conv_std_logic_vector(5320, 16),
19527 => conv_std_logic_vector(5396, 16),
19528 => conv_std_logic_vector(5472, 16),
19529 => conv_std_logic_vector(5548, 16),
19530 => conv_std_logic_vector(5624, 16),
19531 => conv_std_logic_vector(5700, 16),
19532 => conv_std_logic_vector(5776, 16),
19533 => conv_std_logic_vector(5852, 16),
19534 => conv_std_logic_vector(5928, 16),
19535 => conv_std_logic_vector(6004, 16),
19536 => conv_std_logic_vector(6080, 16),
19537 => conv_std_logic_vector(6156, 16),
19538 => conv_std_logic_vector(6232, 16),
19539 => conv_std_logic_vector(6308, 16),
19540 => conv_std_logic_vector(6384, 16),
19541 => conv_std_logic_vector(6460, 16),
19542 => conv_std_logic_vector(6536, 16),
19543 => conv_std_logic_vector(6612, 16),
19544 => conv_std_logic_vector(6688, 16),
19545 => conv_std_logic_vector(6764, 16),
19546 => conv_std_logic_vector(6840, 16),
19547 => conv_std_logic_vector(6916, 16),
19548 => conv_std_logic_vector(6992, 16),
19549 => conv_std_logic_vector(7068, 16),
19550 => conv_std_logic_vector(7144, 16),
19551 => conv_std_logic_vector(7220, 16),
19552 => conv_std_logic_vector(7296, 16),
19553 => conv_std_logic_vector(7372, 16),
19554 => conv_std_logic_vector(7448, 16),
19555 => conv_std_logic_vector(7524, 16),
19556 => conv_std_logic_vector(7600, 16),
19557 => conv_std_logic_vector(7676, 16),
19558 => conv_std_logic_vector(7752, 16),
19559 => conv_std_logic_vector(7828, 16),
19560 => conv_std_logic_vector(7904, 16),
19561 => conv_std_logic_vector(7980, 16),
19562 => conv_std_logic_vector(8056, 16),
19563 => conv_std_logic_vector(8132, 16),
19564 => conv_std_logic_vector(8208, 16),
19565 => conv_std_logic_vector(8284, 16),
19566 => conv_std_logic_vector(8360, 16),
19567 => conv_std_logic_vector(8436, 16),
19568 => conv_std_logic_vector(8512, 16),
19569 => conv_std_logic_vector(8588, 16),
19570 => conv_std_logic_vector(8664, 16),
19571 => conv_std_logic_vector(8740, 16),
19572 => conv_std_logic_vector(8816, 16),
19573 => conv_std_logic_vector(8892, 16),
19574 => conv_std_logic_vector(8968, 16),
19575 => conv_std_logic_vector(9044, 16),
19576 => conv_std_logic_vector(9120, 16),
19577 => conv_std_logic_vector(9196, 16),
19578 => conv_std_logic_vector(9272, 16),
19579 => conv_std_logic_vector(9348, 16),
19580 => conv_std_logic_vector(9424, 16),
19581 => conv_std_logic_vector(9500, 16),
19582 => conv_std_logic_vector(9576, 16),
19583 => conv_std_logic_vector(9652, 16),
19584 => conv_std_logic_vector(9728, 16),
19585 => conv_std_logic_vector(9804, 16),
19586 => conv_std_logic_vector(9880, 16),
19587 => conv_std_logic_vector(9956, 16),
19588 => conv_std_logic_vector(10032, 16),
19589 => conv_std_logic_vector(10108, 16),
19590 => conv_std_logic_vector(10184, 16),
19591 => conv_std_logic_vector(10260, 16),
19592 => conv_std_logic_vector(10336, 16),
19593 => conv_std_logic_vector(10412, 16),
19594 => conv_std_logic_vector(10488, 16),
19595 => conv_std_logic_vector(10564, 16),
19596 => conv_std_logic_vector(10640, 16),
19597 => conv_std_logic_vector(10716, 16),
19598 => conv_std_logic_vector(10792, 16),
19599 => conv_std_logic_vector(10868, 16),
19600 => conv_std_logic_vector(10944, 16),
19601 => conv_std_logic_vector(11020, 16),
19602 => conv_std_logic_vector(11096, 16),
19603 => conv_std_logic_vector(11172, 16),
19604 => conv_std_logic_vector(11248, 16),
19605 => conv_std_logic_vector(11324, 16),
19606 => conv_std_logic_vector(11400, 16),
19607 => conv_std_logic_vector(11476, 16),
19608 => conv_std_logic_vector(11552, 16),
19609 => conv_std_logic_vector(11628, 16),
19610 => conv_std_logic_vector(11704, 16),
19611 => conv_std_logic_vector(11780, 16),
19612 => conv_std_logic_vector(11856, 16),
19613 => conv_std_logic_vector(11932, 16),
19614 => conv_std_logic_vector(12008, 16),
19615 => conv_std_logic_vector(12084, 16),
19616 => conv_std_logic_vector(12160, 16),
19617 => conv_std_logic_vector(12236, 16),
19618 => conv_std_logic_vector(12312, 16),
19619 => conv_std_logic_vector(12388, 16),
19620 => conv_std_logic_vector(12464, 16),
19621 => conv_std_logic_vector(12540, 16),
19622 => conv_std_logic_vector(12616, 16),
19623 => conv_std_logic_vector(12692, 16),
19624 => conv_std_logic_vector(12768, 16),
19625 => conv_std_logic_vector(12844, 16),
19626 => conv_std_logic_vector(12920, 16),
19627 => conv_std_logic_vector(12996, 16),
19628 => conv_std_logic_vector(13072, 16),
19629 => conv_std_logic_vector(13148, 16),
19630 => conv_std_logic_vector(13224, 16),
19631 => conv_std_logic_vector(13300, 16),
19632 => conv_std_logic_vector(13376, 16),
19633 => conv_std_logic_vector(13452, 16),
19634 => conv_std_logic_vector(13528, 16),
19635 => conv_std_logic_vector(13604, 16),
19636 => conv_std_logic_vector(13680, 16),
19637 => conv_std_logic_vector(13756, 16),
19638 => conv_std_logic_vector(13832, 16),
19639 => conv_std_logic_vector(13908, 16),
19640 => conv_std_logic_vector(13984, 16),
19641 => conv_std_logic_vector(14060, 16),
19642 => conv_std_logic_vector(14136, 16),
19643 => conv_std_logic_vector(14212, 16),
19644 => conv_std_logic_vector(14288, 16),
19645 => conv_std_logic_vector(14364, 16),
19646 => conv_std_logic_vector(14440, 16),
19647 => conv_std_logic_vector(14516, 16),
19648 => conv_std_logic_vector(14592, 16),
19649 => conv_std_logic_vector(14668, 16),
19650 => conv_std_logic_vector(14744, 16),
19651 => conv_std_logic_vector(14820, 16),
19652 => conv_std_logic_vector(14896, 16),
19653 => conv_std_logic_vector(14972, 16),
19654 => conv_std_logic_vector(15048, 16),
19655 => conv_std_logic_vector(15124, 16),
19656 => conv_std_logic_vector(15200, 16),
19657 => conv_std_logic_vector(15276, 16),
19658 => conv_std_logic_vector(15352, 16),
19659 => conv_std_logic_vector(15428, 16),
19660 => conv_std_logic_vector(15504, 16),
19661 => conv_std_logic_vector(15580, 16),
19662 => conv_std_logic_vector(15656, 16),
19663 => conv_std_logic_vector(15732, 16),
19664 => conv_std_logic_vector(15808, 16),
19665 => conv_std_logic_vector(15884, 16),
19666 => conv_std_logic_vector(15960, 16),
19667 => conv_std_logic_vector(16036, 16),
19668 => conv_std_logic_vector(16112, 16),
19669 => conv_std_logic_vector(16188, 16),
19670 => conv_std_logic_vector(16264, 16),
19671 => conv_std_logic_vector(16340, 16),
19672 => conv_std_logic_vector(16416, 16),
19673 => conv_std_logic_vector(16492, 16),
19674 => conv_std_logic_vector(16568, 16),
19675 => conv_std_logic_vector(16644, 16),
19676 => conv_std_logic_vector(16720, 16),
19677 => conv_std_logic_vector(16796, 16),
19678 => conv_std_logic_vector(16872, 16),
19679 => conv_std_logic_vector(16948, 16),
19680 => conv_std_logic_vector(17024, 16),
19681 => conv_std_logic_vector(17100, 16),
19682 => conv_std_logic_vector(17176, 16),
19683 => conv_std_logic_vector(17252, 16),
19684 => conv_std_logic_vector(17328, 16),
19685 => conv_std_logic_vector(17404, 16),
19686 => conv_std_logic_vector(17480, 16),
19687 => conv_std_logic_vector(17556, 16),
19688 => conv_std_logic_vector(17632, 16),
19689 => conv_std_logic_vector(17708, 16),
19690 => conv_std_logic_vector(17784, 16),
19691 => conv_std_logic_vector(17860, 16),
19692 => conv_std_logic_vector(17936, 16),
19693 => conv_std_logic_vector(18012, 16),
19694 => conv_std_logic_vector(18088, 16),
19695 => conv_std_logic_vector(18164, 16),
19696 => conv_std_logic_vector(18240, 16),
19697 => conv_std_logic_vector(18316, 16),
19698 => conv_std_logic_vector(18392, 16),
19699 => conv_std_logic_vector(18468, 16),
19700 => conv_std_logic_vector(18544, 16),
19701 => conv_std_logic_vector(18620, 16),
19702 => conv_std_logic_vector(18696, 16),
19703 => conv_std_logic_vector(18772, 16),
19704 => conv_std_logic_vector(18848, 16),
19705 => conv_std_logic_vector(18924, 16),
19706 => conv_std_logic_vector(19000, 16),
19707 => conv_std_logic_vector(19076, 16),
19708 => conv_std_logic_vector(19152, 16),
19709 => conv_std_logic_vector(19228, 16),
19710 => conv_std_logic_vector(19304, 16),
19711 => conv_std_logic_vector(19380, 16),
19712 => conv_std_logic_vector(0, 16),
19713 => conv_std_logic_vector(77, 16),
19714 => conv_std_logic_vector(154, 16),
19715 => conv_std_logic_vector(231, 16),
19716 => conv_std_logic_vector(308, 16),
19717 => conv_std_logic_vector(385, 16),
19718 => conv_std_logic_vector(462, 16),
19719 => conv_std_logic_vector(539, 16),
19720 => conv_std_logic_vector(616, 16),
19721 => conv_std_logic_vector(693, 16),
19722 => conv_std_logic_vector(770, 16),
19723 => conv_std_logic_vector(847, 16),
19724 => conv_std_logic_vector(924, 16),
19725 => conv_std_logic_vector(1001, 16),
19726 => conv_std_logic_vector(1078, 16),
19727 => conv_std_logic_vector(1155, 16),
19728 => conv_std_logic_vector(1232, 16),
19729 => conv_std_logic_vector(1309, 16),
19730 => conv_std_logic_vector(1386, 16),
19731 => conv_std_logic_vector(1463, 16),
19732 => conv_std_logic_vector(1540, 16),
19733 => conv_std_logic_vector(1617, 16),
19734 => conv_std_logic_vector(1694, 16),
19735 => conv_std_logic_vector(1771, 16),
19736 => conv_std_logic_vector(1848, 16),
19737 => conv_std_logic_vector(1925, 16),
19738 => conv_std_logic_vector(2002, 16),
19739 => conv_std_logic_vector(2079, 16),
19740 => conv_std_logic_vector(2156, 16),
19741 => conv_std_logic_vector(2233, 16),
19742 => conv_std_logic_vector(2310, 16),
19743 => conv_std_logic_vector(2387, 16),
19744 => conv_std_logic_vector(2464, 16),
19745 => conv_std_logic_vector(2541, 16),
19746 => conv_std_logic_vector(2618, 16),
19747 => conv_std_logic_vector(2695, 16),
19748 => conv_std_logic_vector(2772, 16),
19749 => conv_std_logic_vector(2849, 16),
19750 => conv_std_logic_vector(2926, 16),
19751 => conv_std_logic_vector(3003, 16),
19752 => conv_std_logic_vector(3080, 16),
19753 => conv_std_logic_vector(3157, 16),
19754 => conv_std_logic_vector(3234, 16),
19755 => conv_std_logic_vector(3311, 16),
19756 => conv_std_logic_vector(3388, 16),
19757 => conv_std_logic_vector(3465, 16),
19758 => conv_std_logic_vector(3542, 16),
19759 => conv_std_logic_vector(3619, 16),
19760 => conv_std_logic_vector(3696, 16),
19761 => conv_std_logic_vector(3773, 16),
19762 => conv_std_logic_vector(3850, 16),
19763 => conv_std_logic_vector(3927, 16),
19764 => conv_std_logic_vector(4004, 16),
19765 => conv_std_logic_vector(4081, 16),
19766 => conv_std_logic_vector(4158, 16),
19767 => conv_std_logic_vector(4235, 16),
19768 => conv_std_logic_vector(4312, 16),
19769 => conv_std_logic_vector(4389, 16),
19770 => conv_std_logic_vector(4466, 16),
19771 => conv_std_logic_vector(4543, 16),
19772 => conv_std_logic_vector(4620, 16),
19773 => conv_std_logic_vector(4697, 16),
19774 => conv_std_logic_vector(4774, 16),
19775 => conv_std_logic_vector(4851, 16),
19776 => conv_std_logic_vector(4928, 16),
19777 => conv_std_logic_vector(5005, 16),
19778 => conv_std_logic_vector(5082, 16),
19779 => conv_std_logic_vector(5159, 16),
19780 => conv_std_logic_vector(5236, 16),
19781 => conv_std_logic_vector(5313, 16),
19782 => conv_std_logic_vector(5390, 16),
19783 => conv_std_logic_vector(5467, 16),
19784 => conv_std_logic_vector(5544, 16),
19785 => conv_std_logic_vector(5621, 16),
19786 => conv_std_logic_vector(5698, 16),
19787 => conv_std_logic_vector(5775, 16),
19788 => conv_std_logic_vector(5852, 16),
19789 => conv_std_logic_vector(5929, 16),
19790 => conv_std_logic_vector(6006, 16),
19791 => conv_std_logic_vector(6083, 16),
19792 => conv_std_logic_vector(6160, 16),
19793 => conv_std_logic_vector(6237, 16),
19794 => conv_std_logic_vector(6314, 16),
19795 => conv_std_logic_vector(6391, 16),
19796 => conv_std_logic_vector(6468, 16),
19797 => conv_std_logic_vector(6545, 16),
19798 => conv_std_logic_vector(6622, 16),
19799 => conv_std_logic_vector(6699, 16),
19800 => conv_std_logic_vector(6776, 16),
19801 => conv_std_logic_vector(6853, 16),
19802 => conv_std_logic_vector(6930, 16),
19803 => conv_std_logic_vector(7007, 16),
19804 => conv_std_logic_vector(7084, 16),
19805 => conv_std_logic_vector(7161, 16),
19806 => conv_std_logic_vector(7238, 16),
19807 => conv_std_logic_vector(7315, 16),
19808 => conv_std_logic_vector(7392, 16),
19809 => conv_std_logic_vector(7469, 16),
19810 => conv_std_logic_vector(7546, 16),
19811 => conv_std_logic_vector(7623, 16),
19812 => conv_std_logic_vector(7700, 16),
19813 => conv_std_logic_vector(7777, 16),
19814 => conv_std_logic_vector(7854, 16),
19815 => conv_std_logic_vector(7931, 16),
19816 => conv_std_logic_vector(8008, 16),
19817 => conv_std_logic_vector(8085, 16),
19818 => conv_std_logic_vector(8162, 16),
19819 => conv_std_logic_vector(8239, 16),
19820 => conv_std_logic_vector(8316, 16),
19821 => conv_std_logic_vector(8393, 16),
19822 => conv_std_logic_vector(8470, 16),
19823 => conv_std_logic_vector(8547, 16),
19824 => conv_std_logic_vector(8624, 16),
19825 => conv_std_logic_vector(8701, 16),
19826 => conv_std_logic_vector(8778, 16),
19827 => conv_std_logic_vector(8855, 16),
19828 => conv_std_logic_vector(8932, 16),
19829 => conv_std_logic_vector(9009, 16),
19830 => conv_std_logic_vector(9086, 16),
19831 => conv_std_logic_vector(9163, 16),
19832 => conv_std_logic_vector(9240, 16),
19833 => conv_std_logic_vector(9317, 16),
19834 => conv_std_logic_vector(9394, 16),
19835 => conv_std_logic_vector(9471, 16),
19836 => conv_std_logic_vector(9548, 16),
19837 => conv_std_logic_vector(9625, 16),
19838 => conv_std_logic_vector(9702, 16),
19839 => conv_std_logic_vector(9779, 16),
19840 => conv_std_logic_vector(9856, 16),
19841 => conv_std_logic_vector(9933, 16),
19842 => conv_std_logic_vector(10010, 16),
19843 => conv_std_logic_vector(10087, 16),
19844 => conv_std_logic_vector(10164, 16),
19845 => conv_std_logic_vector(10241, 16),
19846 => conv_std_logic_vector(10318, 16),
19847 => conv_std_logic_vector(10395, 16),
19848 => conv_std_logic_vector(10472, 16),
19849 => conv_std_logic_vector(10549, 16),
19850 => conv_std_logic_vector(10626, 16),
19851 => conv_std_logic_vector(10703, 16),
19852 => conv_std_logic_vector(10780, 16),
19853 => conv_std_logic_vector(10857, 16),
19854 => conv_std_logic_vector(10934, 16),
19855 => conv_std_logic_vector(11011, 16),
19856 => conv_std_logic_vector(11088, 16),
19857 => conv_std_logic_vector(11165, 16),
19858 => conv_std_logic_vector(11242, 16),
19859 => conv_std_logic_vector(11319, 16),
19860 => conv_std_logic_vector(11396, 16),
19861 => conv_std_logic_vector(11473, 16),
19862 => conv_std_logic_vector(11550, 16),
19863 => conv_std_logic_vector(11627, 16),
19864 => conv_std_logic_vector(11704, 16),
19865 => conv_std_logic_vector(11781, 16),
19866 => conv_std_logic_vector(11858, 16),
19867 => conv_std_logic_vector(11935, 16),
19868 => conv_std_logic_vector(12012, 16),
19869 => conv_std_logic_vector(12089, 16),
19870 => conv_std_logic_vector(12166, 16),
19871 => conv_std_logic_vector(12243, 16),
19872 => conv_std_logic_vector(12320, 16),
19873 => conv_std_logic_vector(12397, 16),
19874 => conv_std_logic_vector(12474, 16),
19875 => conv_std_logic_vector(12551, 16),
19876 => conv_std_logic_vector(12628, 16),
19877 => conv_std_logic_vector(12705, 16),
19878 => conv_std_logic_vector(12782, 16),
19879 => conv_std_logic_vector(12859, 16),
19880 => conv_std_logic_vector(12936, 16),
19881 => conv_std_logic_vector(13013, 16),
19882 => conv_std_logic_vector(13090, 16),
19883 => conv_std_logic_vector(13167, 16),
19884 => conv_std_logic_vector(13244, 16),
19885 => conv_std_logic_vector(13321, 16),
19886 => conv_std_logic_vector(13398, 16),
19887 => conv_std_logic_vector(13475, 16),
19888 => conv_std_logic_vector(13552, 16),
19889 => conv_std_logic_vector(13629, 16),
19890 => conv_std_logic_vector(13706, 16),
19891 => conv_std_logic_vector(13783, 16),
19892 => conv_std_logic_vector(13860, 16),
19893 => conv_std_logic_vector(13937, 16),
19894 => conv_std_logic_vector(14014, 16),
19895 => conv_std_logic_vector(14091, 16),
19896 => conv_std_logic_vector(14168, 16),
19897 => conv_std_logic_vector(14245, 16),
19898 => conv_std_logic_vector(14322, 16),
19899 => conv_std_logic_vector(14399, 16),
19900 => conv_std_logic_vector(14476, 16),
19901 => conv_std_logic_vector(14553, 16),
19902 => conv_std_logic_vector(14630, 16),
19903 => conv_std_logic_vector(14707, 16),
19904 => conv_std_logic_vector(14784, 16),
19905 => conv_std_logic_vector(14861, 16),
19906 => conv_std_logic_vector(14938, 16),
19907 => conv_std_logic_vector(15015, 16),
19908 => conv_std_logic_vector(15092, 16),
19909 => conv_std_logic_vector(15169, 16),
19910 => conv_std_logic_vector(15246, 16),
19911 => conv_std_logic_vector(15323, 16),
19912 => conv_std_logic_vector(15400, 16),
19913 => conv_std_logic_vector(15477, 16),
19914 => conv_std_logic_vector(15554, 16),
19915 => conv_std_logic_vector(15631, 16),
19916 => conv_std_logic_vector(15708, 16),
19917 => conv_std_logic_vector(15785, 16),
19918 => conv_std_logic_vector(15862, 16),
19919 => conv_std_logic_vector(15939, 16),
19920 => conv_std_logic_vector(16016, 16),
19921 => conv_std_logic_vector(16093, 16),
19922 => conv_std_logic_vector(16170, 16),
19923 => conv_std_logic_vector(16247, 16),
19924 => conv_std_logic_vector(16324, 16),
19925 => conv_std_logic_vector(16401, 16),
19926 => conv_std_logic_vector(16478, 16),
19927 => conv_std_logic_vector(16555, 16),
19928 => conv_std_logic_vector(16632, 16),
19929 => conv_std_logic_vector(16709, 16),
19930 => conv_std_logic_vector(16786, 16),
19931 => conv_std_logic_vector(16863, 16),
19932 => conv_std_logic_vector(16940, 16),
19933 => conv_std_logic_vector(17017, 16),
19934 => conv_std_logic_vector(17094, 16),
19935 => conv_std_logic_vector(17171, 16),
19936 => conv_std_logic_vector(17248, 16),
19937 => conv_std_logic_vector(17325, 16),
19938 => conv_std_logic_vector(17402, 16),
19939 => conv_std_logic_vector(17479, 16),
19940 => conv_std_logic_vector(17556, 16),
19941 => conv_std_logic_vector(17633, 16),
19942 => conv_std_logic_vector(17710, 16),
19943 => conv_std_logic_vector(17787, 16),
19944 => conv_std_logic_vector(17864, 16),
19945 => conv_std_logic_vector(17941, 16),
19946 => conv_std_logic_vector(18018, 16),
19947 => conv_std_logic_vector(18095, 16),
19948 => conv_std_logic_vector(18172, 16),
19949 => conv_std_logic_vector(18249, 16),
19950 => conv_std_logic_vector(18326, 16),
19951 => conv_std_logic_vector(18403, 16),
19952 => conv_std_logic_vector(18480, 16),
19953 => conv_std_logic_vector(18557, 16),
19954 => conv_std_logic_vector(18634, 16),
19955 => conv_std_logic_vector(18711, 16),
19956 => conv_std_logic_vector(18788, 16),
19957 => conv_std_logic_vector(18865, 16),
19958 => conv_std_logic_vector(18942, 16),
19959 => conv_std_logic_vector(19019, 16),
19960 => conv_std_logic_vector(19096, 16),
19961 => conv_std_logic_vector(19173, 16),
19962 => conv_std_logic_vector(19250, 16),
19963 => conv_std_logic_vector(19327, 16),
19964 => conv_std_logic_vector(19404, 16),
19965 => conv_std_logic_vector(19481, 16),
19966 => conv_std_logic_vector(19558, 16),
19967 => conv_std_logic_vector(19635, 16),
19968 => conv_std_logic_vector(0, 16),
19969 => conv_std_logic_vector(78, 16),
19970 => conv_std_logic_vector(156, 16),
19971 => conv_std_logic_vector(234, 16),
19972 => conv_std_logic_vector(312, 16),
19973 => conv_std_logic_vector(390, 16),
19974 => conv_std_logic_vector(468, 16),
19975 => conv_std_logic_vector(546, 16),
19976 => conv_std_logic_vector(624, 16),
19977 => conv_std_logic_vector(702, 16),
19978 => conv_std_logic_vector(780, 16),
19979 => conv_std_logic_vector(858, 16),
19980 => conv_std_logic_vector(936, 16),
19981 => conv_std_logic_vector(1014, 16),
19982 => conv_std_logic_vector(1092, 16),
19983 => conv_std_logic_vector(1170, 16),
19984 => conv_std_logic_vector(1248, 16),
19985 => conv_std_logic_vector(1326, 16),
19986 => conv_std_logic_vector(1404, 16),
19987 => conv_std_logic_vector(1482, 16),
19988 => conv_std_logic_vector(1560, 16),
19989 => conv_std_logic_vector(1638, 16),
19990 => conv_std_logic_vector(1716, 16),
19991 => conv_std_logic_vector(1794, 16),
19992 => conv_std_logic_vector(1872, 16),
19993 => conv_std_logic_vector(1950, 16),
19994 => conv_std_logic_vector(2028, 16),
19995 => conv_std_logic_vector(2106, 16),
19996 => conv_std_logic_vector(2184, 16),
19997 => conv_std_logic_vector(2262, 16),
19998 => conv_std_logic_vector(2340, 16),
19999 => conv_std_logic_vector(2418, 16),
20000 => conv_std_logic_vector(2496, 16),
20001 => conv_std_logic_vector(2574, 16),
20002 => conv_std_logic_vector(2652, 16),
20003 => conv_std_logic_vector(2730, 16),
20004 => conv_std_logic_vector(2808, 16),
20005 => conv_std_logic_vector(2886, 16),
20006 => conv_std_logic_vector(2964, 16),
20007 => conv_std_logic_vector(3042, 16),
20008 => conv_std_logic_vector(3120, 16),
20009 => conv_std_logic_vector(3198, 16),
20010 => conv_std_logic_vector(3276, 16),
20011 => conv_std_logic_vector(3354, 16),
20012 => conv_std_logic_vector(3432, 16),
20013 => conv_std_logic_vector(3510, 16),
20014 => conv_std_logic_vector(3588, 16),
20015 => conv_std_logic_vector(3666, 16),
20016 => conv_std_logic_vector(3744, 16),
20017 => conv_std_logic_vector(3822, 16),
20018 => conv_std_logic_vector(3900, 16),
20019 => conv_std_logic_vector(3978, 16),
20020 => conv_std_logic_vector(4056, 16),
20021 => conv_std_logic_vector(4134, 16),
20022 => conv_std_logic_vector(4212, 16),
20023 => conv_std_logic_vector(4290, 16),
20024 => conv_std_logic_vector(4368, 16),
20025 => conv_std_logic_vector(4446, 16),
20026 => conv_std_logic_vector(4524, 16),
20027 => conv_std_logic_vector(4602, 16),
20028 => conv_std_logic_vector(4680, 16),
20029 => conv_std_logic_vector(4758, 16),
20030 => conv_std_logic_vector(4836, 16),
20031 => conv_std_logic_vector(4914, 16),
20032 => conv_std_logic_vector(4992, 16),
20033 => conv_std_logic_vector(5070, 16),
20034 => conv_std_logic_vector(5148, 16),
20035 => conv_std_logic_vector(5226, 16),
20036 => conv_std_logic_vector(5304, 16),
20037 => conv_std_logic_vector(5382, 16),
20038 => conv_std_logic_vector(5460, 16),
20039 => conv_std_logic_vector(5538, 16),
20040 => conv_std_logic_vector(5616, 16),
20041 => conv_std_logic_vector(5694, 16),
20042 => conv_std_logic_vector(5772, 16),
20043 => conv_std_logic_vector(5850, 16),
20044 => conv_std_logic_vector(5928, 16),
20045 => conv_std_logic_vector(6006, 16),
20046 => conv_std_logic_vector(6084, 16),
20047 => conv_std_logic_vector(6162, 16),
20048 => conv_std_logic_vector(6240, 16),
20049 => conv_std_logic_vector(6318, 16),
20050 => conv_std_logic_vector(6396, 16),
20051 => conv_std_logic_vector(6474, 16),
20052 => conv_std_logic_vector(6552, 16),
20053 => conv_std_logic_vector(6630, 16),
20054 => conv_std_logic_vector(6708, 16),
20055 => conv_std_logic_vector(6786, 16),
20056 => conv_std_logic_vector(6864, 16),
20057 => conv_std_logic_vector(6942, 16),
20058 => conv_std_logic_vector(7020, 16),
20059 => conv_std_logic_vector(7098, 16),
20060 => conv_std_logic_vector(7176, 16),
20061 => conv_std_logic_vector(7254, 16),
20062 => conv_std_logic_vector(7332, 16),
20063 => conv_std_logic_vector(7410, 16),
20064 => conv_std_logic_vector(7488, 16),
20065 => conv_std_logic_vector(7566, 16),
20066 => conv_std_logic_vector(7644, 16),
20067 => conv_std_logic_vector(7722, 16),
20068 => conv_std_logic_vector(7800, 16),
20069 => conv_std_logic_vector(7878, 16),
20070 => conv_std_logic_vector(7956, 16),
20071 => conv_std_logic_vector(8034, 16),
20072 => conv_std_logic_vector(8112, 16),
20073 => conv_std_logic_vector(8190, 16),
20074 => conv_std_logic_vector(8268, 16),
20075 => conv_std_logic_vector(8346, 16),
20076 => conv_std_logic_vector(8424, 16),
20077 => conv_std_logic_vector(8502, 16),
20078 => conv_std_logic_vector(8580, 16),
20079 => conv_std_logic_vector(8658, 16),
20080 => conv_std_logic_vector(8736, 16),
20081 => conv_std_logic_vector(8814, 16),
20082 => conv_std_logic_vector(8892, 16),
20083 => conv_std_logic_vector(8970, 16),
20084 => conv_std_logic_vector(9048, 16),
20085 => conv_std_logic_vector(9126, 16),
20086 => conv_std_logic_vector(9204, 16),
20087 => conv_std_logic_vector(9282, 16),
20088 => conv_std_logic_vector(9360, 16),
20089 => conv_std_logic_vector(9438, 16),
20090 => conv_std_logic_vector(9516, 16),
20091 => conv_std_logic_vector(9594, 16),
20092 => conv_std_logic_vector(9672, 16),
20093 => conv_std_logic_vector(9750, 16),
20094 => conv_std_logic_vector(9828, 16),
20095 => conv_std_logic_vector(9906, 16),
20096 => conv_std_logic_vector(9984, 16),
20097 => conv_std_logic_vector(10062, 16),
20098 => conv_std_logic_vector(10140, 16),
20099 => conv_std_logic_vector(10218, 16),
20100 => conv_std_logic_vector(10296, 16),
20101 => conv_std_logic_vector(10374, 16),
20102 => conv_std_logic_vector(10452, 16),
20103 => conv_std_logic_vector(10530, 16),
20104 => conv_std_logic_vector(10608, 16),
20105 => conv_std_logic_vector(10686, 16),
20106 => conv_std_logic_vector(10764, 16),
20107 => conv_std_logic_vector(10842, 16),
20108 => conv_std_logic_vector(10920, 16),
20109 => conv_std_logic_vector(10998, 16),
20110 => conv_std_logic_vector(11076, 16),
20111 => conv_std_logic_vector(11154, 16),
20112 => conv_std_logic_vector(11232, 16),
20113 => conv_std_logic_vector(11310, 16),
20114 => conv_std_logic_vector(11388, 16),
20115 => conv_std_logic_vector(11466, 16),
20116 => conv_std_logic_vector(11544, 16),
20117 => conv_std_logic_vector(11622, 16),
20118 => conv_std_logic_vector(11700, 16),
20119 => conv_std_logic_vector(11778, 16),
20120 => conv_std_logic_vector(11856, 16),
20121 => conv_std_logic_vector(11934, 16),
20122 => conv_std_logic_vector(12012, 16),
20123 => conv_std_logic_vector(12090, 16),
20124 => conv_std_logic_vector(12168, 16),
20125 => conv_std_logic_vector(12246, 16),
20126 => conv_std_logic_vector(12324, 16),
20127 => conv_std_logic_vector(12402, 16),
20128 => conv_std_logic_vector(12480, 16),
20129 => conv_std_logic_vector(12558, 16),
20130 => conv_std_logic_vector(12636, 16),
20131 => conv_std_logic_vector(12714, 16),
20132 => conv_std_logic_vector(12792, 16),
20133 => conv_std_logic_vector(12870, 16),
20134 => conv_std_logic_vector(12948, 16),
20135 => conv_std_logic_vector(13026, 16),
20136 => conv_std_logic_vector(13104, 16),
20137 => conv_std_logic_vector(13182, 16),
20138 => conv_std_logic_vector(13260, 16),
20139 => conv_std_logic_vector(13338, 16),
20140 => conv_std_logic_vector(13416, 16),
20141 => conv_std_logic_vector(13494, 16),
20142 => conv_std_logic_vector(13572, 16),
20143 => conv_std_logic_vector(13650, 16),
20144 => conv_std_logic_vector(13728, 16),
20145 => conv_std_logic_vector(13806, 16),
20146 => conv_std_logic_vector(13884, 16),
20147 => conv_std_logic_vector(13962, 16),
20148 => conv_std_logic_vector(14040, 16),
20149 => conv_std_logic_vector(14118, 16),
20150 => conv_std_logic_vector(14196, 16),
20151 => conv_std_logic_vector(14274, 16),
20152 => conv_std_logic_vector(14352, 16),
20153 => conv_std_logic_vector(14430, 16),
20154 => conv_std_logic_vector(14508, 16),
20155 => conv_std_logic_vector(14586, 16),
20156 => conv_std_logic_vector(14664, 16),
20157 => conv_std_logic_vector(14742, 16),
20158 => conv_std_logic_vector(14820, 16),
20159 => conv_std_logic_vector(14898, 16),
20160 => conv_std_logic_vector(14976, 16),
20161 => conv_std_logic_vector(15054, 16),
20162 => conv_std_logic_vector(15132, 16),
20163 => conv_std_logic_vector(15210, 16),
20164 => conv_std_logic_vector(15288, 16),
20165 => conv_std_logic_vector(15366, 16),
20166 => conv_std_logic_vector(15444, 16),
20167 => conv_std_logic_vector(15522, 16),
20168 => conv_std_logic_vector(15600, 16),
20169 => conv_std_logic_vector(15678, 16),
20170 => conv_std_logic_vector(15756, 16),
20171 => conv_std_logic_vector(15834, 16),
20172 => conv_std_logic_vector(15912, 16),
20173 => conv_std_logic_vector(15990, 16),
20174 => conv_std_logic_vector(16068, 16),
20175 => conv_std_logic_vector(16146, 16),
20176 => conv_std_logic_vector(16224, 16),
20177 => conv_std_logic_vector(16302, 16),
20178 => conv_std_logic_vector(16380, 16),
20179 => conv_std_logic_vector(16458, 16),
20180 => conv_std_logic_vector(16536, 16),
20181 => conv_std_logic_vector(16614, 16),
20182 => conv_std_logic_vector(16692, 16),
20183 => conv_std_logic_vector(16770, 16),
20184 => conv_std_logic_vector(16848, 16),
20185 => conv_std_logic_vector(16926, 16),
20186 => conv_std_logic_vector(17004, 16),
20187 => conv_std_logic_vector(17082, 16),
20188 => conv_std_logic_vector(17160, 16),
20189 => conv_std_logic_vector(17238, 16),
20190 => conv_std_logic_vector(17316, 16),
20191 => conv_std_logic_vector(17394, 16),
20192 => conv_std_logic_vector(17472, 16),
20193 => conv_std_logic_vector(17550, 16),
20194 => conv_std_logic_vector(17628, 16),
20195 => conv_std_logic_vector(17706, 16),
20196 => conv_std_logic_vector(17784, 16),
20197 => conv_std_logic_vector(17862, 16),
20198 => conv_std_logic_vector(17940, 16),
20199 => conv_std_logic_vector(18018, 16),
20200 => conv_std_logic_vector(18096, 16),
20201 => conv_std_logic_vector(18174, 16),
20202 => conv_std_logic_vector(18252, 16),
20203 => conv_std_logic_vector(18330, 16),
20204 => conv_std_logic_vector(18408, 16),
20205 => conv_std_logic_vector(18486, 16),
20206 => conv_std_logic_vector(18564, 16),
20207 => conv_std_logic_vector(18642, 16),
20208 => conv_std_logic_vector(18720, 16),
20209 => conv_std_logic_vector(18798, 16),
20210 => conv_std_logic_vector(18876, 16),
20211 => conv_std_logic_vector(18954, 16),
20212 => conv_std_logic_vector(19032, 16),
20213 => conv_std_logic_vector(19110, 16),
20214 => conv_std_logic_vector(19188, 16),
20215 => conv_std_logic_vector(19266, 16),
20216 => conv_std_logic_vector(19344, 16),
20217 => conv_std_logic_vector(19422, 16),
20218 => conv_std_logic_vector(19500, 16),
20219 => conv_std_logic_vector(19578, 16),
20220 => conv_std_logic_vector(19656, 16),
20221 => conv_std_logic_vector(19734, 16),
20222 => conv_std_logic_vector(19812, 16),
20223 => conv_std_logic_vector(19890, 16),
20224 => conv_std_logic_vector(0, 16),
20225 => conv_std_logic_vector(79, 16),
20226 => conv_std_logic_vector(158, 16),
20227 => conv_std_logic_vector(237, 16),
20228 => conv_std_logic_vector(316, 16),
20229 => conv_std_logic_vector(395, 16),
20230 => conv_std_logic_vector(474, 16),
20231 => conv_std_logic_vector(553, 16),
20232 => conv_std_logic_vector(632, 16),
20233 => conv_std_logic_vector(711, 16),
20234 => conv_std_logic_vector(790, 16),
20235 => conv_std_logic_vector(869, 16),
20236 => conv_std_logic_vector(948, 16),
20237 => conv_std_logic_vector(1027, 16),
20238 => conv_std_logic_vector(1106, 16),
20239 => conv_std_logic_vector(1185, 16),
20240 => conv_std_logic_vector(1264, 16),
20241 => conv_std_logic_vector(1343, 16),
20242 => conv_std_logic_vector(1422, 16),
20243 => conv_std_logic_vector(1501, 16),
20244 => conv_std_logic_vector(1580, 16),
20245 => conv_std_logic_vector(1659, 16),
20246 => conv_std_logic_vector(1738, 16),
20247 => conv_std_logic_vector(1817, 16),
20248 => conv_std_logic_vector(1896, 16),
20249 => conv_std_logic_vector(1975, 16),
20250 => conv_std_logic_vector(2054, 16),
20251 => conv_std_logic_vector(2133, 16),
20252 => conv_std_logic_vector(2212, 16),
20253 => conv_std_logic_vector(2291, 16),
20254 => conv_std_logic_vector(2370, 16),
20255 => conv_std_logic_vector(2449, 16),
20256 => conv_std_logic_vector(2528, 16),
20257 => conv_std_logic_vector(2607, 16),
20258 => conv_std_logic_vector(2686, 16),
20259 => conv_std_logic_vector(2765, 16),
20260 => conv_std_logic_vector(2844, 16),
20261 => conv_std_logic_vector(2923, 16),
20262 => conv_std_logic_vector(3002, 16),
20263 => conv_std_logic_vector(3081, 16),
20264 => conv_std_logic_vector(3160, 16),
20265 => conv_std_logic_vector(3239, 16),
20266 => conv_std_logic_vector(3318, 16),
20267 => conv_std_logic_vector(3397, 16),
20268 => conv_std_logic_vector(3476, 16),
20269 => conv_std_logic_vector(3555, 16),
20270 => conv_std_logic_vector(3634, 16),
20271 => conv_std_logic_vector(3713, 16),
20272 => conv_std_logic_vector(3792, 16),
20273 => conv_std_logic_vector(3871, 16),
20274 => conv_std_logic_vector(3950, 16),
20275 => conv_std_logic_vector(4029, 16),
20276 => conv_std_logic_vector(4108, 16),
20277 => conv_std_logic_vector(4187, 16),
20278 => conv_std_logic_vector(4266, 16),
20279 => conv_std_logic_vector(4345, 16),
20280 => conv_std_logic_vector(4424, 16),
20281 => conv_std_logic_vector(4503, 16),
20282 => conv_std_logic_vector(4582, 16),
20283 => conv_std_logic_vector(4661, 16),
20284 => conv_std_logic_vector(4740, 16),
20285 => conv_std_logic_vector(4819, 16),
20286 => conv_std_logic_vector(4898, 16),
20287 => conv_std_logic_vector(4977, 16),
20288 => conv_std_logic_vector(5056, 16),
20289 => conv_std_logic_vector(5135, 16),
20290 => conv_std_logic_vector(5214, 16),
20291 => conv_std_logic_vector(5293, 16),
20292 => conv_std_logic_vector(5372, 16),
20293 => conv_std_logic_vector(5451, 16),
20294 => conv_std_logic_vector(5530, 16),
20295 => conv_std_logic_vector(5609, 16),
20296 => conv_std_logic_vector(5688, 16),
20297 => conv_std_logic_vector(5767, 16),
20298 => conv_std_logic_vector(5846, 16),
20299 => conv_std_logic_vector(5925, 16),
20300 => conv_std_logic_vector(6004, 16),
20301 => conv_std_logic_vector(6083, 16),
20302 => conv_std_logic_vector(6162, 16),
20303 => conv_std_logic_vector(6241, 16),
20304 => conv_std_logic_vector(6320, 16),
20305 => conv_std_logic_vector(6399, 16),
20306 => conv_std_logic_vector(6478, 16),
20307 => conv_std_logic_vector(6557, 16),
20308 => conv_std_logic_vector(6636, 16),
20309 => conv_std_logic_vector(6715, 16),
20310 => conv_std_logic_vector(6794, 16),
20311 => conv_std_logic_vector(6873, 16),
20312 => conv_std_logic_vector(6952, 16),
20313 => conv_std_logic_vector(7031, 16),
20314 => conv_std_logic_vector(7110, 16),
20315 => conv_std_logic_vector(7189, 16),
20316 => conv_std_logic_vector(7268, 16),
20317 => conv_std_logic_vector(7347, 16),
20318 => conv_std_logic_vector(7426, 16),
20319 => conv_std_logic_vector(7505, 16),
20320 => conv_std_logic_vector(7584, 16),
20321 => conv_std_logic_vector(7663, 16),
20322 => conv_std_logic_vector(7742, 16),
20323 => conv_std_logic_vector(7821, 16),
20324 => conv_std_logic_vector(7900, 16),
20325 => conv_std_logic_vector(7979, 16),
20326 => conv_std_logic_vector(8058, 16),
20327 => conv_std_logic_vector(8137, 16),
20328 => conv_std_logic_vector(8216, 16),
20329 => conv_std_logic_vector(8295, 16),
20330 => conv_std_logic_vector(8374, 16),
20331 => conv_std_logic_vector(8453, 16),
20332 => conv_std_logic_vector(8532, 16),
20333 => conv_std_logic_vector(8611, 16),
20334 => conv_std_logic_vector(8690, 16),
20335 => conv_std_logic_vector(8769, 16),
20336 => conv_std_logic_vector(8848, 16),
20337 => conv_std_logic_vector(8927, 16),
20338 => conv_std_logic_vector(9006, 16),
20339 => conv_std_logic_vector(9085, 16),
20340 => conv_std_logic_vector(9164, 16),
20341 => conv_std_logic_vector(9243, 16),
20342 => conv_std_logic_vector(9322, 16),
20343 => conv_std_logic_vector(9401, 16),
20344 => conv_std_logic_vector(9480, 16),
20345 => conv_std_logic_vector(9559, 16),
20346 => conv_std_logic_vector(9638, 16),
20347 => conv_std_logic_vector(9717, 16),
20348 => conv_std_logic_vector(9796, 16),
20349 => conv_std_logic_vector(9875, 16),
20350 => conv_std_logic_vector(9954, 16),
20351 => conv_std_logic_vector(10033, 16),
20352 => conv_std_logic_vector(10112, 16),
20353 => conv_std_logic_vector(10191, 16),
20354 => conv_std_logic_vector(10270, 16),
20355 => conv_std_logic_vector(10349, 16),
20356 => conv_std_logic_vector(10428, 16),
20357 => conv_std_logic_vector(10507, 16),
20358 => conv_std_logic_vector(10586, 16),
20359 => conv_std_logic_vector(10665, 16),
20360 => conv_std_logic_vector(10744, 16),
20361 => conv_std_logic_vector(10823, 16),
20362 => conv_std_logic_vector(10902, 16),
20363 => conv_std_logic_vector(10981, 16),
20364 => conv_std_logic_vector(11060, 16),
20365 => conv_std_logic_vector(11139, 16),
20366 => conv_std_logic_vector(11218, 16),
20367 => conv_std_logic_vector(11297, 16),
20368 => conv_std_logic_vector(11376, 16),
20369 => conv_std_logic_vector(11455, 16),
20370 => conv_std_logic_vector(11534, 16),
20371 => conv_std_logic_vector(11613, 16),
20372 => conv_std_logic_vector(11692, 16),
20373 => conv_std_logic_vector(11771, 16),
20374 => conv_std_logic_vector(11850, 16),
20375 => conv_std_logic_vector(11929, 16),
20376 => conv_std_logic_vector(12008, 16),
20377 => conv_std_logic_vector(12087, 16),
20378 => conv_std_logic_vector(12166, 16),
20379 => conv_std_logic_vector(12245, 16),
20380 => conv_std_logic_vector(12324, 16),
20381 => conv_std_logic_vector(12403, 16),
20382 => conv_std_logic_vector(12482, 16),
20383 => conv_std_logic_vector(12561, 16),
20384 => conv_std_logic_vector(12640, 16),
20385 => conv_std_logic_vector(12719, 16),
20386 => conv_std_logic_vector(12798, 16),
20387 => conv_std_logic_vector(12877, 16),
20388 => conv_std_logic_vector(12956, 16),
20389 => conv_std_logic_vector(13035, 16),
20390 => conv_std_logic_vector(13114, 16),
20391 => conv_std_logic_vector(13193, 16),
20392 => conv_std_logic_vector(13272, 16),
20393 => conv_std_logic_vector(13351, 16),
20394 => conv_std_logic_vector(13430, 16),
20395 => conv_std_logic_vector(13509, 16),
20396 => conv_std_logic_vector(13588, 16),
20397 => conv_std_logic_vector(13667, 16),
20398 => conv_std_logic_vector(13746, 16),
20399 => conv_std_logic_vector(13825, 16),
20400 => conv_std_logic_vector(13904, 16),
20401 => conv_std_logic_vector(13983, 16),
20402 => conv_std_logic_vector(14062, 16),
20403 => conv_std_logic_vector(14141, 16),
20404 => conv_std_logic_vector(14220, 16),
20405 => conv_std_logic_vector(14299, 16),
20406 => conv_std_logic_vector(14378, 16),
20407 => conv_std_logic_vector(14457, 16),
20408 => conv_std_logic_vector(14536, 16),
20409 => conv_std_logic_vector(14615, 16),
20410 => conv_std_logic_vector(14694, 16),
20411 => conv_std_logic_vector(14773, 16),
20412 => conv_std_logic_vector(14852, 16),
20413 => conv_std_logic_vector(14931, 16),
20414 => conv_std_logic_vector(15010, 16),
20415 => conv_std_logic_vector(15089, 16),
20416 => conv_std_logic_vector(15168, 16),
20417 => conv_std_logic_vector(15247, 16),
20418 => conv_std_logic_vector(15326, 16),
20419 => conv_std_logic_vector(15405, 16),
20420 => conv_std_logic_vector(15484, 16),
20421 => conv_std_logic_vector(15563, 16),
20422 => conv_std_logic_vector(15642, 16),
20423 => conv_std_logic_vector(15721, 16),
20424 => conv_std_logic_vector(15800, 16),
20425 => conv_std_logic_vector(15879, 16),
20426 => conv_std_logic_vector(15958, 16),
20427 => conv_std_logic_vector(16037, 16),
20428 => conv_std_logic_vector(16116, 16),
20429 => conv_std_logic_vector(16195, 16),
20430 => conv_std_logic_vector(16274, 16),
20431 => conv_std_logic_vector(16353, 16),
20432 => conv_std_logic_vector(16432, 16),
20433 => conv_std_logic_vector(16511, 16),
20434 => conv_std_logic_vector(16590, 16),
20435 => conv_std_logic_vector(16669, 16),
20436 => conv_std_logic_vector(16748, 16),
20437 => conv_std_logic_vector(16827, 16),
20438 => conv_std_logic_vector(16906, 16),
20439 => conv_std_logic_vector(16985, 16),
20440 => conv_std_logic_vector(17064, 16),
20441 => conv_std_logic_vector(17143, 16),
20442 => conv_std_logic_vector(17222, 16),
20443 => conv_std_logic_vector(17301, 16),
20444 => conv_std_logic_vector(17380, 16),
20445 => conv_std_logic_vector(17459, 16),
20446 => conv_std_logic_vector(17538, 16),
20447 => conv_std_logic_vector(17617, 16),
20448 => conv_std_logic_vector(17696, 16),
20449 => conv_std_logic_vector(17775, 16),
20450 => conv_std_logic_vector(17854, 16),
20451 => conv_std_logic_vector(17933, 16),
20452 => conv_std_logic_vector(18012, 16),
20453 => conv_std_logic_vector(18091, 16),
20454 => conv_std_logic_vector(18170, 16),
20455 => conv_std_logic_vector(18249, 16),
20456 => conv_std_logic_vector(18328, 16),
20457 => conv_std_logic_vector(18407, 16),
20458 => conv_std_logic_vector(18486, 16),
20459 => conv_std_logic_vector(18565, 16),
20460 => conv_std_logic_vector(18644, 16),
20461 => conv_std_logic_vector(18723, 16),
20462 => conv_std_logic_vector(18802, 16),
20463 => conv_std_logic_vector(18881, 16),
20464 => conv_std_logic_vector(18960, 16),
20465 => conv_std_logic_vector(19039, 16),
20466 => conv_std_logic_vector(19118, 16),
20467 => conv_std_logic_vector(19197, 16),
20468 => conv_std_logic_vector(19276, 16),
20469 => conv_std_logic_vector(19355, 16),
20470 => conv_std_logic_vector(19434, 16),
20471 => conv_std_logic_vector(19513, 16),
20472 => conv_std_logic_vector(19592, 16),
20473 => conv_std_logic_vector(19671, 16),
20474 => conv_std_logic_vector(19750, 16),
20475 => conv_std_logic_vector(19829, 16),
20476 => conv_std_logic_vector(19908, 16),
20477 => conv_std_logic_vector(19987, 16),
20478 => conv_std_logic_vector(20066, 16),
20479 => conv_std_logic_vector(20145, 16),
20480 => conv_std_logic_vector(0, 16),
20481 => conv_std_logic_vector(80, 16),
20482 => conv_std_logic_vector(160, 16),
20483 => conv_std_logic_vector(240, 16),
20484 => conv_std_logic_vector(320, 16),
20485 => conv_std_logic_vector(400, 16),
20486 => conv_std_logic_vector(480, 16),
20487 => conv_std_logic_vector(560, 16),
20488 => conv_std_logic_vector(640, 16),
20489 => conv_std_logic_vector(720, 16),
20490 => conv_std_logic_vector(800, 16),
20491 => conv_std_logic_vector(880, 16),
20492 => conv_std_logic_vector(960, 16),
20493 => conv_std_logic_vector(1040, 16),
20494 => conv_std_logic_vector(1120, 16),
20495 => conv_std_logic_vector(1200, 16),
20496 => conv_std_logic_vector(1280, 16),
20497 => conv_std_logic_vector(1360, 16),
20498 => conv_std_logic_vector(1440, 16),
20499 => conv_std_logic_vector(1520, 16),
20500 => conv_std_logic_vector(1600, 16),
20501 => conv_std_logic_vector(1680, 16),
20502 => conv_std_logic_vector(1760, 16),
20503 => conv_std_logic_vector(1840, 16),
20504 => conv_std_logic_vector(1920, 16),
20505 => conv_std_logic_vector(2000, 16),
20506 => conv_std_logic_vector(2080, 16),
20507 => conv_std_logic_vector(2160, 16),
20508 => conv_std_logic_vector(2240, 16),
20509 => conv_std_logic_vector(2320, 16),
20510 => conv_std_logic_vector(2400, 16),
20511 => conv_std_logic_vector(2480, 16),
20512 => conv_std_logic_vector(2560, 16),
20513 => conv_std_logic_vector(2640, 16),
20514 => conv_std_logic_vector(2720, 16),
20515 => conv_std_logic_vector(2800, 16),
20516 => conv_std_logic_vector(2880, 16),
20517 => conv_std_logic_vector(2960, 16),
20518 => conv_std_logic_vector(3040, 16),
20519 => conv_std_logic_vector(3120, 16),
20520 => conv_std_logic_vector(3200, 16),
20521 => conv_std_logic_vector(3280, 16),
20522 => conv_std_logic_vector(3360, 16),
20523 => conv_std_logic_vector(3440, 16),
20524 => conv_std_logic_vector(3520, 16),
20525 => conv_std_logic_vector(3600, 16),
20526 => conv_std_logic_vector(3680, 16),
20527 => conv_std_logic_vector(3760, 16),
20528 => conv_std_logic_vector(3840, 16),
20529 => conv_std_logic_vector(3920, 16),
20530 => conv_std_logic_vector(4000, 16),
20531 => conv_std_logic_vector(4080, 16),
20532 => conv_std_logic_vector(4160, 16),
20533 => conv_std_logic_vector(4240, 16),
20534 => conv_std_logic_vector(4320, 16),
20535 => conv_std_logic_vector(4400, 16),
20536 => conv_std_logic_vector(4480, 16),
20537 => conv_std_logic_vector(4560, 16),
20538 => conv_std_logic_vector(4640, 16),
20539 => conv_std_logic_vector(4720, 16),
20540 => conv_std_logic_vector(4800, 16),
20541 => conv_std_logic_vector(4880, 16),
20542 => conv_std_logic_vector(4960, 16),
20543 => conv_std_logic_vector(5040, 16),
20544 => conv_std_logic_vector(5120, 16),
20545 => conv_std_logic_vector(5200, 16),
20546 => conv_std_logic_vector(5280, 16),
20547 => conv_std_logic_vector(5360, 16),
20548 => conv_std_logic_vector(5440, 16),
20549 => conv_std_logic_vector(5520, 16),
20550 => conv_std_logic_vector(5600, 16),
20551 => conv_std_logic_vector(5680, 16),
20552 => conv_std_logic_vector(5760, 16),
20553 => conv_std_logic_vector(5840, 16),
20554 => conv_std_logic_vector(5920, 16),
20555 => conv_std_logic_vector(6000, 16),
20556 => conv_std_logic_vector(6080, 16),
20557 => conv_std_logic_vector(6160, 16),
20558 => conv_std_logic_vector(6240, 16),
20559 => conv_std_logic_vector(6320, 16),
20560 => conv_std_logic_vector(6400, 16),
20561 => conv_std_logic_vector(6480, 16),
20562 => conv_std_logic_vector(6560, 16),
20563 => conv_std_logic_vector(6640, 16),
20564 => conv_std_logic_vector(6720, 16),
20565 => conv_std_logic_vector(6800, 16),
20566 => conv_std_logic_vector(6880, 16),
20567 => conv_std_logic_vector(6960, 16),
20568 => conv_std_logic_vector(7040, 16),
20569 => conv_std_logic_vector(7120, 16),
20570 => conv_std_logic_vector(7200, 16),
20571 => conv_std_logic_vector(7280, 16),
20572 => conv_std_logic_vector(7360, 16),
20573 => conv_std_logic_vector(7440, 16),
20574 => conv_std_logic_vector(7520, 16),
20575 => conv_std_logic_vector(7600, 16),
20576 => conv_std_logic_vector(7680, 16),
20577 => conv_std_logic_vector(7760, 16),
20578 => conv_std_logic_vector(7840, 16),
20579 => conv_std_logic_vector(7920, 16),
20580 => conv_std_logic_vector(8000, 16),
20581 => conv_std_logic_vector(8080, 16),
20582 => conv_std_logic_vector(8160, 16),
20583 => conv_std_logic_vector(8240, 16),
20584 => conv_std_logic_vector(8320, 16),
20585 => conv_std_logic_vector(8400, 16),
20586 => conv_std_logic_vector(8480, 16),
20587 => conv_std_logic_vector(8560, 16),
20588 => conv_std_logic_vector(8640, 16),
20589 => conv_std_logic_vector(8720, 16),
20590 => conv_std_logic_vector(8800, 16),
20591 => conv_std_logic_vector(8880, 16),
20592 => conv_std_logic_vector(8960, 16),
20593 => conv_std_logic_vector(9040, 16),
20594 => conv_std_logic_vector(9120, 16),
20595 => conv_std_logic_vector(9200, 16),
20596 => conv_std_logic_vector(9280, 16),
20597 => conv_std_logic_vector(9360, 16),
20598 => conv_std_logic_vector(9440, 16),
20599 => conv_std_logic_vector(9520, 16),
20600 => conv_std_logic_vector(9600, 16),
20601 => conv_std_logic_vector(9680, 16),
20602 => conv_std_logic_vector(9760, 16),
20603 => conv_std_logic_vector(9840, 16),
20604 => conv_std_logic_vector(9920, 16),
20605 => conv_std_logic_vector(10000, 16),
20606 => conv_std_logic_vector(10080, 16),
20607 => conv_std_logic_vector(10160, 16),
20608 => conv_std_logic_vector(10240, 16),
20609 => conv_std_logic_vector(10320, 16),
20610 => conv_std_logic_vector(10400, 16),
20611 => conv_std_logic_vector(10480, 16),
20612 => conv_std_logic_vector(10560, 16),
20613 => conv_std_logic_vector(10640, 16),
20614 => conv_std_logic_vector(10720, 16),
20615 => conv_std_logic_vector(10800, 16),
20616 => conv_std_logic_vector(10880, 16),
20617 => conv_std_logic_vector(10960, 16),
20618 => conv_std_logic_vector(11040, 16),
20619 => conv_std_logic_vector(11120, 16),
20620 => conv_std_logic_vector(11200, 16),
20621 => conv_std_logic_vector(11280, 16),
20622 => conv_std_logic_vector(11360, 16),
20623 => conv_std_logic_vector(11440, 16),
20624 => conv_std_logic_vector(11520, 16),
20625 => conv_std_logic_vector(11600, 16),
20626 => conv_std_logic_vector(11680, 16),
20627 => conv_std_logic_vector(11760, 16),
20628 => conv_std_logic_vector(11840, 16),
20629 => conv_std_logic_vector(11920, 16),
20630 => conv_std_logic_vector(12000, 16),
20631 => conv_std_logic_vector(12080, 16),
20632 => conv_std_logic_vector(12160, 16),
20633 => conv_std_logic_vector(12240, 16),
20634 => conv_std_logic_vector(12320, 16),
20635 => conv_std_logic_vector(12400, 16),
20636 => conv_std_logic_vector(12480, 16),
20637 => conv_std_logic_vector(12560, 16),
20638 => conv_std_logic_vector(12640, 16),
20639 => conv_std_logic_vector(12720, 16),
20640 => conv_std_logic_vector(12800, 16),
20641 => conv_std_logic_vector(12880, 16),
20642 => conv_std_logic_vector(12960, 16),
20643 => conv_std_logic_vector(13040, 16),
20644 => conv_std_logic_vector(13120, 16),
20645 => conv_std_logic_vector(13200, 16),
20646 => conv_std_logic_vector(13280, 16),
20647 => conv_std_logic_vector(13360, 16),
20648 => conv_std_logic_vector(13440, 16),
20649 => conv_std_logic_vector(13520, 16),
20650 => conv_std_logic_vector(13600, 16),
20651 => conv_std_logic_vector(13680, 16),
20652 => conv_std_logic_vector(13760, 16),
20653 => conv_std_logic_vector(13840, 16),
20654 => conv_std_logic_vector(13920, 16),
20655 => conv_std_logic_vector(14000, 16),
20656 => conv_std_logic_vector(14080, 16),
20657 => conv_std_logic_vector(14160, 16),
20658 => conv_std_logic_vector(14240, 16),
20659 => conv_std_logic_vector(14320, 16),
20660 => conv_std_logic_vector(14400, 16),
20661 => conv_std_logic_vector(14480, 16),
20662 => conv_std_logic_vector(14560, 16),
20663 => conv_std_logic_vector(14640, 16),
20664 => conv_std_logic_vector(14720, 16),
20665 => conv_std_logic_vector(14800, 16),
20666 => conv_std_logic_vector(14880, 16),
20667 => conv_std_logic_vector(14960, 16),
20668 => conv_std_logic_vector(15040, 16),
20669 => conv_std_logic_vector(15120, 16),
20670 => conv_std_logic_vector(15200, 16),
20671 => conv_std_logic_vector(15280, 16),
20672 => conv_std_logic_vector(15360, 16),
20673 => conv_std_logic_vector(15440, 16),
20674 => conv_std_logic_vector(15520, 16),
20675 => conv_std_logic_vector(15600, 16),
20676 => conv_std_logic_vector(15680, 16),
20677 => conv_std_logic_vector(15760, 16),
20678 => conv_std_logic_vector(15840, 16),
20679 => conv_std_logic_vector(15920, 16),
20680 => conv_std_logic_vector(16000, 16),
20681 => conv_std_logic_vector(16080, 16),
20682 => conv_std_logic_vector(16160, 16),
20683 => conv_std_logic_vector(16240, 16),
20684 => conv_std_logic_vector(16320, 16),
20685 => conv_std_logic_vector(16400, 16),
20686 => conv_std_logic_vector(16480, 16),
20687 => conv_std_logic_vector(16560, 16),
20688 => conv_std_logic_vector(16640, 16),
20689 => conv_std_logic_vector(16720, 16),
20690 => conv_std_logic_vector(16800, 16),
20691 => conv_std_logic_vector(16880, 16),
20692 => conv_std_logic_vector(16960, 16),
20693 => conv_std_logic_vector(17040, 16),
20694 => conv_std_logic_vector(17120, 16),
20695 => conv_std_logic_vector(17200, 16),
20696 => conv_std_logic_vector(17280, 16),
20697 => conv_std_logic_vector(17360, 16),
20698 => conv_std_logic_vector(17440, 16),
20699 => conv_std_logic_vector(17520, 16),
20700 => conv_std_logic_vector(17600, 16),
20701 => conv_std_logic_vector(17680, 16),
20702 => conv_std_logic_vector(17760, 16),
20703 => conv_std_logic_vector(17840, 16),
20704 => conv_std_logic_vector(17920, 16),
20705 => conv_std_logic_vector(18000, 16),
20706 => conv_std_logic_vector(18080, 16),
20707 => conv_std_logic_vector(18160, 16),
20708 => conv_std_logic_vector(18240, 16),
20709 => conv_std_logic_vector(18320, 16),
20710 => conv_std_logic_vector(18400, 16),
20711 => conv_std_logic_vector(18480, 16),
20712 => conv_std_logic_vector(18560, 16),
20713 => conv_std_logic_vector(18640, 16),
20714 => conv_std_logic_vector(18720, 16),
20715 => conv_std_logic_vector(18800, 16),
20716 => conv_std_logic_vector(18880, 16),
20717 => conv_std_logic_vector(18960, 16),
20718 => conv_std_logic_vector(19040, 16),
20719 => conv_std_logic_vector(19120, 16),
20720 => conv_std_logic_vector(19200, 16),
20721 => conv_std_logic_vector(19280, 16),
20722 => conv_std_logic_vector(19360, 16),
20723 => conv_std_logic_vector(19440, 16),
20724 => conv_std_logic_vector(19520, 16),
20725 => conv_std_logic_vector(19600, 16),
20726 => conv_std_logic_vector(19680, 16),
20727 => conv_std_logic_vector(19760, 16),
20728 => conv_std_logic_vector(19840, 16),
20729 => conv_std_logic_vector(19920, 16),
20730 => conv_std_logic_vector(20000, 16),
20731 => conv_std_logic_vector(20080, 16),
20732 => conv_std_logic_vector(20160, 16),
20733 => conv_std_logic_vector(20240, 16),
20734 => conv_std_logic_vector(20320, 16),
20735 => conv_std_logic_vector(20400, 16),
20736 => conv_std_logic_vector(0, 16),
20737 => conv_std_logic_vector(81, 16),
20738 => conv_std_logic_vector(162, 16),
20739 => conv_std_logic_vector(243, 16),
20740 => conv_std_logic_vector(324, 16),
20741 => conv_std_logic_vector(405, 16),
20742 => conv_std_logic_vector(486, 16),
20743 => conv_std_logic_vector(567, 16),
20744 => conv_std_logic_vector(648, 16),
20745 => conv_std_logic_vector(729, 16),
20746 => conv_std_logic_vector(810, 16),
20747 => conv_std_logic_vector(891, 16),
20748 => conv_std_logic_vector(972, 16),
20749 => conv_std_logic_vector(1053, 16),
20750 => conv_std_logic_vector(1134, 16),
20751 => conv_std_logic_vector(1215, 16),
20752 => conv_std_logic_vector(1296, 16),
20753 => conv_std_logic_vector(1377, 16),
20754 => conv_std_logic_vector(1458, 16),
20755 => conv_std_logic_vector(1539, 16),
20756 => conv_std_logic_vector(1620, 16),
20757 => conv_std_logic_vector(1701, 16),
20758 => conv_std_logic_vector(1782, 16),
20759 => conv_std_logic_vector(1863, 16),
20760 => conv_std_logic_vector(1944, 16),
20761 => conv_std_logic_vector(2025, 16),
20762 => conv_std_logic_vector(2106, 16),
20763 => conv_std_logic_vector(2187, 16),
20764 => conv_std_logic_vector(2268, 16),
20765 => conv_std_logic_vector(2349, 16),
20766 => conv_std_logic_vector(2430, 16),
20767 => conv_std_logic_vector(2511, 16),
20768 => conv_std_logic_vector(2592, 16),
20769 => conv_std_logic_vector(2673, 16),
20770 => conv_std_logic_vector(2754, 16),
20771 => conv_std_logic_vector(2835, 16),
20772 => conv_std_logic_vector(2916, 16),
20773 => conv_std_logic_vector(2997, 16),
20774 => conv_std_logic_vector(3078, 16),
20775 => conv_std_logic_vector(3159, 16),
20776 => conv_std_logic_vector(3240, 16),
20777 => conv_std_logic_vector(3321, 16),
20778 => conv_std_logic_vector(3402, 16),
20779 => conv_std_logic_vector(3483, 16),
20780 => conv_std_logic_vector(3564, 16),
20781 => conv_std_logic_vector(3645, 16),
20782 => conv_std_logic_vector(3726, 16),
20783 => conv_std_logic_vector(3807, 16),
20784 => conv_std_logic_vector(3888, 16),
20785 => conv_std_logic_vector(3969, 16),
20786 => conv_std_logic_vector(4050, 16),
20787 => conv_std_logic_vector(4131, 16),
20788 => conv_std_logic_vector(4212, 16),
20789 => conv_std_logic_vector(4293, 16),
20790 => conv_std_logic_vector(4374, 16),
20791 => conv_std_logic_vector(4455, 16),
20792 => conv_std_logic_vector(4536, 16),
20793 => conv_std_logic_vector(4617, 16),
20794 => conv_std_logic_vector(4698, 16),
20795 => conv_std_logic_vector(4779, 16),
20796 => conv_std_logic_vector(4860, 16),
20797 => conv_std_logic_vector(4941, 16),
20798 => conv_std_logic_vector(5022, 16),
20799 => conv_std_logic_vector(5103, 16),
20800 => conv_std_logic_vector(5184, 16),
20801 => conv_std_logic_vector(5265, 16),
20802 => conv_std_logic_vector(5346, 16),
20803 => conv_std_logic_vector(5427, 16),
20804 => conv_std_logic_vector(5508, 16),
20805 => conv_std_logic_vector(5589, 16),
20806 => conv_std_logic_vector(5670, 16),
20807 => conv_std_logic_vector(5751, 16),
20808 => conv_std_logic_vector(5832, 16),
20809 => conv_std_logic_vector(5913, 16),
20810 => conv_std_logic_vector(5994, 16),
20811 => conv_std_logic_vector(6075, 16),
20812 => conv_std_logic_vector(6156, 16),
20813 => conv_std_logic_vector(6237, 16),
20814 => conv_std_logic_vector(6318, 16),
20815 => conv_std_logic_vector(6399, 16),
20816 => conv_std_logic_vector(6480, 16),
20817 => conv_std_logic_vector(6561, 16),
20818 => conv_std_logic_vector(6642, 16),
20819 => conv_std_logic_vector(6723, 16),
20820 => conv_std_logic_vector(6804, 16),
20821 => conv_std_logic_vector(6885, 16),
20822 => conv_std_logic_vector(6966, 16),
20823 => conv_std_logic_vector(7047, 16),
20824 => conv_std_logic_vector(7128, 16),
20825 => conv_std_logic_vector(7209, 16),
20826 => conv_std_logic_vector(7290, 16),
20827 => conv_std_logic_vector(7371, 16),
20828 => conv_std_logic_vector(7452, 16),
20829 => conv_std_logic_vector(7533, 16),
20830 => conv_std_logic_vector(7614, 16),
20831 => conv_std_logic_vector(7695, 16),
20832 => conv_std_logic_vector(7776, 16),
20833 => conv_std_logic_vector(7857, 16),
20834 => conv_std_logic_vector(7938, 16),
20835 => conv_std_logic_vector(8019, 16),
20836 => conv_std_logic_vector(8100, 16),
20837 => conv_std_logic_vector(8181, 16),
20838 => conv_std_logic_vector(8262, 16),
20839 => conv_std_logic_vector(8343, 16),
20840 => conv_std_logic_vector(8424, 16),
20841 => conv_std_logic_vector(8505, 16),
20842 => conv_std_logic_vector(8586, 16),
20843 => conv_std_logic_vector(8667, 16),
20844 => conv_std_logic_vector(8748, 16),
20845 => conv_std_logic_vector(8829, 16),
20846 => conv_std_logic_vector(8910, 16),
20847 => conv_std_logic_vector(8991, 16),
20848 => conv_std_logic_vector(9072, 16),
20849 => conv_std_logic_vector(9153, 16),
20850 => conv_std_logic_vector(9234, 16),
20851 => conv_std_logic_vector(9315, 16),
20852 => conv_std_logic_vector(9396, 16),
20853 => conv_std_logic_vector(9477, 16),
20854 => conv_std_logic_vector(9558, 16),
20855 => conv_std_logic_vector(9639, 16),
20856 => conv_std_logic_vector(9720, 16),
20857 => conv_std_logic_vector(9801, 16),
20858 => conv_std_logic_vector(9882, 16),
20859 => conv_std_logic_vector(9963, 16),
20860 => conv_std_logic_vector(10044, 16),
20861 => conv_std_logic_vector(10125, 16),
20862 => conv_std_logic_vector(10206, 16),
20863 => conv_std_logic_vector(10287, 16),
20864 => conv_std_logic_vector(10368, 16),
20865 => conv_std_logic_vector(10449, 16),
20866 => conv_std_logic_vector(10530, 16),
20867 => conv_std_logic_vector(10611, 16),
20868 => conv_std_logic_vector(10692, 16),
20869 => conv_std_logic_vector(10773, 16),
20870 => conv_std_logic_vector(10854, 16),
20871 => conv_std_logic_vector(10935, 16),
20872 => conv_std_logic_vector(11016, 16),
20873 => conv_std_logic_vector(11097, 16),
20874 => conv_std_logic_vector(11178, 16),
20875 => conv_std_logic_vector(11259, 16),
20876 => conv_std_logic_vector(11340, 16),
20877 => conv_std_logic_vector(11421, 16),
20878 => conv_std_logic_vector(11502, 16),
20879 => conv_std_logic_vector(11583, 16),
20880 => conv_std_logic_vector(11664, 16),
20881 => conv_std_logic_vector(11745, 16),
20882 => conv_std_logic_vector(11826, 16),
20883 => conv_std_logic_vector(11907, 16),
20884 => conv_std_logic_vector(11988, 16),
20885 => conv_std_logic_vector(12069, 16),
20886 => conv_std_logic_vector(12150, 16),
20887 => conv_std_logic_vector(12231, 16),
20888 => conv_std_logic_vector(12312, 16),
20889 => conv_std_logic_vector(12393, 16),
20890 => conv_std_logic_vector(12474, 16),
20891 => conv_std_logic_vector(12555, 16),
20892 => conv_std_logic_vector(12636, 16),
20893 => conv_std_logic_vector(12717, 16),
20894 => conv_std_logic_vector(12798, 16),
20895 => conv_std_logic_vector(12879, 16),
20896 => conv_std_logic_vector(12960, 16),
20897 => conv_std_logic_vector(13041, 16),
20898 => conv_std_logic_vector(13122, 16),
20899 => conv_std_logic_vector(13203, 16),
20900 => conv_std_logic_vector(13284, 16),
20901 => conv_std_logic_vector(13365, 16),
20902 => conv_std_logic_vector(13446, 16),
20903 => conv_std_logic_vector(13527, 16),
20904 => conv_std_logic_vector(13608, 16),
20905 => conv_std_logic_vector(13689, 16),
20906 => conv_std_logic_vector(13770, 16),
20907 => conv_std_logic_vector(13851, 16),
20908 => conv_std_logic_vector(13932, 16),
20909 => conv_std_logic_vector(14013, 16),
20910 => conv_std_logic_vector(14094, 16),
20911 => conv_std_logic_vector(14175, 16),
20912 => conv_std_logic_vector(14256, 16),
20913 => conv_std_logic_vector(14337, 16),
20914 => conv_std_logic_vector(14418, 16),
20915 => conv_std_logic_vector(14499, 16),
20916 => conv_std_logic_vector(14580, 16),
20917 => conv_std_logic_vector(14661, 16),
20918 => conv_std_logic_vector(14742, 16),
20919 => conv_std_logic_vector(14823, 16),
20920 => conv_std_logic_vector(14904, 16),
20921 => conv_std_logic_vector(14985, 16),
20922 => conv_std_logic_vector(15066, 16),
20923 => conv_std_logic_vector(15147, 16),
20924 => conv_std_logic_vector(15228, 16),
20925 => conv_std_logic_vector(15309, 16),
20926 => conv_std_logic_vector(15390, 16),
20927 => conv_std_logic_vector(15471, 16),
20928 => conv_std_logic_vector(15552, 16),
20929 => conv_std_logic_vector(15633, 16),
20930 => conv_std_logic_vector(15714, 16),
20931 => conv_std_logic_vector(15795, 16),
20932 => conv_std_logic_vector(15876, 16),
20933 => conv_std_logic_vector(15957, 16),
20934 => conv_std_logic_vector(16038, 16),
20935 => conv_std_logic_vector(16119, 16),
20936 => conv_std_logic_vector(16200, 16),
20937 => conv_std_logic_vector(16281, 16),
20938 => conv_std_logic_vector(16362, 16),
20939 => conv_std_logic_vector(16443, 16),
20940 => conv_std_logic_vector(16524, 16),
20941 => conv_std_logic_vector(16605, 16),
20942 => conv_std_logic_vector(16686, 16),
20943 => conv_std_logic_vector(16767, 16),
20944 => conv_std_logic_vector(16848, 16),
20945 => conv_std_logic_vector(16929, 16),
20946 => conv_std_logic_vector(17010, 16),
20947 => conv_std_logic_vector(17091, 16),
20948 => conv_std_logic_vector(17172, 16),
20949 => conv_std_logic_vector(17253, 16),
20950 => conv_std_logic_vector(17334, 16),
20951 => conv_std_logic_vector(17415, 16),
20952 => conv_std_logic_vector(17496, 16),
20953 => conv_std_logic_vector(17577, 16),
20954 => conv_std_logic_vector(17658, 16),
20955 => conv_std_logic_vector(17739, 16),
20956 => conv_std_logic_vector(17820, 16),
20957 => conv_std_logic_vector(17901, 16),
20958 => conv_std_logic_vector(17982, 16),
20959 => conv_std_logic_vector(18063, 16),
20960 => conv_std_logic_vector(18144, 16),
20961 => conv_std_logic_vector(18225, 16),
20962 => conv_std_logic_vector(18306, 16),
20963 => conv_std_logic_vector(18387, 16),
20964 => conv_std_logic_vector(18468, 16),
20965 => conv_std_logic_vector(18549, 16),
20966 => conv_std_logic_vector(18630, 16),
20967 => conv_std_logic_vector(18711, 16),
20968 => conv_std_logic_vector(18792, 16),
20969 => conv_std_logic_vector(18873, 16),
20970 => conv_std_logic_vector(18954, 16),
20971 => conv_std_logic_vector(19035, 16),
20972 => conv_std_logic_vector(19116, 16),
20973 => conv_std_logic_vector(19197, 16),
20974 => conv_std_logic_vector(19278, 16),
20975 => conv_std_logic_vector(19359, 16),
20976 => conv_std_logic_vector(19440, 16),
20977 => conv_std_logic_vector(19521, 16),
20978 => conv_std_logic_vector(19602, 16),
20979 => conv_std_logic_vector(19683, 16),
20980 => conv_std_logic_vector(19764, 16),
20981 => conv_std_logic_vector(19845, 16),
20982 => conv_std_logic_vector(19926, 16),
20983 => conv_std_logic_vector(20007, 16),
20984 => conv_std_logic_vector(20088, 16),
20985 => conv_std_logic_vector(20169, 16),
20986 => conv_std_logic_vector(20250, 16),
20987 => conv_std_logic_vector(20331, 16),
20988 => conv_std_logic_vector(20412, 16),
20989 => conv_std_logic_vector(20493, 16),
20990 => conv_std_logic_vector(20574, 16),
20991 => conv_std_logic_vector(20655, 16),
20992 => conv_std_logic_vector(0, 16),
20993 => conv_std_logic_vector(82, 16),
20994 => conv_std_logic_vector(164, 16),
20995 => conv_std_logic_vector(246, 16),
20996 => conv_std_logic_vector(328, 16),
20997 => conv_std_logic_vector(410, 16),
20998 => conv_std_logic_vector(492, 16),
20999 => conv_std_logic_vector(574, 16),
21000 => conv_std_logic_vector(656, 16),
21001 => conv_std_logic_vector(738, 16),
21002 => conv_std_logic_vector(820, 16),
21003 => conv_std_logic_vector(902, 16),
21004 => conv_std_logic_vector(984, 16),
21005 => conv_std_logic_vector(1066, 16),
21006 => conv_std_logic_vector(1148, 16),
21007 => conv_std_logic_vector(1230, 16),
21008 => conv_std_logic_vector(1312, 16),
21009 => conv_std_logic_vector(1394, 16),
21010 => conv_std_logic_vector(1476, 16),
21011 => conv_std_logic_vector(1558, 16),
21012 => conv_std_logic_vector(1640, 16),
21013 => conv_std_logic_vector(1722, 16),
21014 => conv_std_logic_vector(1804, 16),
21015 => conv_std_logic_vector(1886, 16),
21016 => conv_std_logic_vector(1968, 16),
21017 => conv_std_logic_vector(2050, 16),
21018 => conv_std_logic_vector(2132, 16),
21019 => conv_std_logic_vector(2214, 16),
21020 => conv_std_logic_vector(2296, 16),
21021 => conv_std_logic_vector(2378, 16),
21022 => conv_std_logic_vector(2460, 16),
21023 => conv_std_logic_vector(2542, 16),
21024 => conv_std_logic_vector(2624, 16),
21025 => conv_std_logic_vector(2706, 16),
21026 => conv_std_logic_vector(2788, 16),
21027 => conv_std_logic_vector(2870, 16),
21028 => conv_std_logic_vector(2952, 16),
21029 => conv_std_logic_vector(3034, 16),
21030 => conv_std_logic_vector(3116, 16),
21031 => conv_std_logic_vector(3198, 16),
21032 => conv_std_logic_vector(3280, 16),
21033 => conv_std_logic_vector(3362, 16),
21034 => conv_std_logic_vector(3444, 16),
21035 => conv_std_logic_vector(3526, 16),
21036 => conv_std_logic_vector(3608, 16),
21037 => conv_std_logic_vector(3690, 16),
21038 => conv_std_logic_vector(3772, 16),
21039 => conv_std_logic_vector(3854, 16),
21040 => conv_std_logic_vector(3936, 16),
21041 => conv_std_logic_vector(4018, 16),
21042 => conv_std_logic_vector(4100, 16),
21043 => conv_std_logic_vector(4182, 16),
21044 => conv_std_logic_vector(4264, 16),
21045 => conv_std_logic_vector(4346, 16),
21046 => conv_std_logic_vector(4428, 16),
21047 => conv_std_logic_vector(4510, 16),
21048 => conv_std_logic_vector(4592, 16),
21049 => conv_std_logic_vector(4674, 16),
21050 => conv_std_logic_vector(4756, 16),
21051 => conv_std_logic_vector(4838, 16),
21052 => conv_std_logic_vector(4920, 16),
21053 => conv_std_logic_vector(5002, 16),
21054 => conv_std_logic_vector(5084, 16),
21055 => conv_std_logic_vector(5166, 16),
21056 => conv_std_logic_vector(5248, 16),
21057 => conv_std_logic_vector(5330, 16),
21058 => conv_std_logic_vector(5412, 16),
21059 => conv_std_logic_vector(5494, 16),
21060 => conv_std_logic_vector(5576, 16),
21061 => conv_std_logic_vector(5658, 16),
21062 => conv_std_logic_vector(5740, 16),
21063 => conv_std_logic_vector(5822, 16),
21064 => conv_std_logic_vector(5904, 16),
21065 => conv_std_logic_vector(5986, 16),
21066 => conv_std_logic_vector(6068, 16),
21067 => conv_std_logic_vector(6150, 16),
21068 => conv_std_logic_vector(6232, 16),
21069 => conv_std_logic_vector(6314, 16),
21070 => conv_std_logic_vector(6396, 16),
21071 => conv_std_logic_vector(6478, 16),
21072 => conv_std_logic_vector(6560, 16),
21073 => conv_std_logic_vector(6642, 16),
21074 => conv_std_logic_vector(6724, 16),
21075 => conv_std_logic_vector(6806, 16),
21076 => conv_std_logic_vector(6888, 16),
21077 => conv_std_logic_vector(6970, 16),
21078 => conv_std_logic_vector(7052, 16),
21079 => conv_std_logic_vector(7134, 16),
21080 => conv_std_logic_vector(7216, 16),
21081 => conv_std_logic_vector(7298, 16),
21082 => conv_std_logic_vector(7380, 16),
21083 => conv_std_logic_vector(7462, 16),
21084 => conv_std_logic_vector(7544, 16),
21085 => conv_std_logic_vector(7626, 16),
21086 => conv_std_logic_vector(7708, 16),
21087 => conv_std_logic_vector(7790, 16),
21088 => conv_std_logic_vector(7872, 16),
21089 => conv_std_logic_vector(7954, 16),
21090 => conv_std_logic_vector(8036, 16),
21091 => conv_std_logic_vector(8118, 16),
21092 => conv_std_logic_vector(8200, 16),
21093 => conv_std_logic_vector(8282, 16),
21094 => conv_std_logic_vector(8364, 16),
21095 => conv_std_logic_vector(8446, 16),
21096 => conv_std_logic_vector(8528, 16),
21097 => conv_std_logic_vector(8610, 16),
21098 => conv_std_logic_vector(8692, 16),
21099 => conv_std_logic_vector(8774, 16),
21100 => conv_std_logic_vector(8856, 16),
21101 => conv_std_logic_vector(8938, 16),
21102 => conv_std_logic_vector(9020, 16),
21103 => conv_std_logic_vector(9102, 16),
21104 => conv_std_logic_vector(9184, 16),
21105 => conv_std_logic_vector(9266, 16),
21106 => conv_std_logic_vector(9348, 16),
21107 => conv_std_logic_vector(9430, 16),
21108 => conv_std_logic_vector(9512, 16),
21109 => conv_std_logic_vector(9594, 16),
21110 => conv_std_logic_vector(9676, 16),
21111 => conv_std_logic_vector(9758, 16),
21112 => conv_std_logic_vector(9840, 16),
21113 => conv_std_logic_vector(9922, 16),
21114 => conv_std_logic_vector(10004, 16),
21115 => conv_std_logic_vector(10086, 16),
21116 => conv_std_logic_vector(10168, 16),
21117 => conv_std_logic_vector(10250, 16),
21118 => conv_std_logic_vector(10332, 16),
21119 => conv_std_logic_vector(10414, 16),
21120 => conv_std_logic_vector(10496, 16),
21121 => conv_std_logic_vector(10578, 16),
21122 => conv_std_logic_vector(10660, 16),
21123 => conv_std_logic_vector(10742, 16),
21124 => conv_std_logic_vector(10824, 16),
21125 => conv_std_logic_vector(10906, 16),
21126 => conv_std_logic_vector(10988, 16),
21127 => conv_std_logic_vector(11070, 16),
21128 => conv_std_logic_vector(11152, 16),
21129 => conv_std_logic_vector(11234, 16),
21130 => conv_std_logic_vector(11316, 16),
21131 => conv_std_logic_vector(11398, 16),
21132 => conv_std_logic_vector(11480, 16),
21133 => conv_std_logic_vector(11562, 16),
21134 => conv_std_logic_vector(11644, 16),
21135 => conv_std_logic_vector(11726, 16),
21136 => conv_std_logic_vector(11808, 16),
21137 => conv_std_logic_vector(11890, 16),
21138 => conv_std_logic_vector(11972, 16),
21139 => conv_std_logic_vector(12054, 16),
21140 => conv_std_logic_vector(12136, 16),
21141 => conv_std_logic_vector(12218, 16),
21142 => conv_std_logic_vector(12300, 16),
21143 => conv_std_logic_vector(12382, 16),
21144 => conv_std_logic_vector(12464, 16),
21145 => conv_std_logic_vector(12546, 16),
21146 => conv_std_logic_vector(12628, 16),
21147 => conv_std_logic_vector(12710, 16),
21148 => conv_std_logic_vector(12792, 16),
21149 => conv_std_logic_vector(12874, 16),
21150 => conv_std_logic_vector(12956, 16),
21151 => conv_std_logic_vector(13038, 16),
21152 => conv_std_logic_vector(13120, 16),
21153 => conv_std_logic_vector(13202, 16),
21154 => conv_std_logic_vector(13284, 16),
21155 => conv_std_logic_vector(13366, 16),
21156 => conv_std_logic_vector(13448, 16),
21157 => conv_std_logic_vector(13530, 16),
21158 => conv_std_logic_vector(13612, 16),
21159 => conv_std_logic_vector(13694, 16),
21160 => conv_std_logic_vector(13776, 16),
21161 => conv_std_logic_vector(13858, 16),
21162 => conv_std_logic_vector(13940, 16),
21163 => conv_std_logic_vector(14022, 16),
21164 => conv_std_logic_vector(14104, 16),
21165 => conv_std_logic_vector(14186, 16),
21166 => conv_std_logic_vector(14268, 16),
21167 => conv_std_logic_vector(14350, 16),
21168 => conv_std_logic_vector(14432, 16),
21169 => conv_std_logic_vector(14514, 16),
21170 => conv_std_logic_vector(14596, 16),
21171 => conv_std_logic_vector(14678, 16),
21172 => conv_std_logic_vector(14760, 16),
21173 => conv_std_logic_vector(14842, 16),
21174 => conv_std_logic_vector(14924, 16),
21175 => conv_std_logic_vector(15006, 16),
21176 => conv_std_logic_vector(15088, 16),
21177 => conv_std_logic_vector(15170, 16),
21178 => conv_std_logic_vector(15252, 16),
21179 => conv_std_logic_vector(15334, 16),
21180 => conv_std_logic_vector(15416, 16),
21181 => conv_std_logic_vector(15498, 16),
21182 => conv_std_logic_vector(15580, 16),
21183 => conv_std_logic_vector(15662, 16),
21184 => conv_std_logic_vector(15744, 16),
21185 => conv_std_logic_vector(15826, 16),
21186 => conv_std_logic_vector(15908, 16),
21187 => conv_std_logic_vector(15990, 16),
21188 => conv_std_logic_vector(16072, 16),
21189 => conv_std_logic_vector(16154, 16),
21190 => conv_std_logic_vector(16236, 16),
21191 => conv_std_logic_vector(16318, 16),
21192 => conv_std_logic_vector(16400, 16),
21193 => conv_std_logic_vector(16482, 16),
21194 => conv_std_logic_vector(16564, 16),
21195 => conv_std_logic_vector(16646, 16),
21196 => conv_std_logic_vector(16728, 16),
21197 => conv_std_logic_vector(16810, 16),
21198 => conv_std_logic_vector(16892, 16),
21199 => conv_std_logic_vector(16974, 16),
21200 => conv_std_logic_vector(17056, 16),
21201 => conv_std_logic_vector(17138, 16),
21202 => conv_std_logic_vector(17220, 16),
21203 => conv_std_logic_vector(17302, 16),
21204 => conv_std_logic_vector(17384, 16),
21205 => conv_std_logic_vector(17466, 16),
21206 => conv_std_logic_vector(17548, 16),
21207 => conv_std_logic_vector(17630, 16),
21208 => conv_std_logic_vector(17712, 16),
21209 => conv_std_logic_vector(17794, 16),
21210 => conv_std_logic_vector(17876, 16),
21211 => conv_std_logic_vector(17958, 16),
21212 => conv_std_logic_vector(18040, 16),
21213 => conv_std_logic_vector(18122, 16),
21214 => conv_std_logic_vector(18204, 16),
21215 => conv_std_logic_vector(18286, 16),
21216 => conv_std_logic_vector(18368, 16),
21217 => conv_std_logic_vector(18450, 16),
21218 => conv_std_logic_vector(18532, 16),
21219 => conv_std_logic_vector(18614, 16),
21220 => conv_std_logic_vector(18696, 16),
21221 => conv_std_logic_vector(18778, 16),
21222 => conv_std_logic_vector(18860, 16),
21223 => conv_std_logic_vector(18942, 16),
21224 => conv_std_logic_vector(19024, 16),
21225 => conv_std_logic_vector(19106, 16),
21226 => conv_std_logic_vector(19188, 16),
21227 => conv_std_logic_vector(19270, 16),
21228 => conv_std_logic_vector(19352, 16),
21229 => conv_std_logic_vector(19434, 16),
21230 => conv_std_logic_vector(19516, 16),
21231 => conv_std_logic_vector(19598, 16),
21232 => conv_std_logic_vector(19680, 16),
21233 => conv_std_logic_vector(19762, 16),
21234 => conv_std_logic_vector(19844, 16),
21235 => conv_std_logic_vector(19926, 16),
21236 => conv_std_logic_vector(20008, 16),
21237 => conv_std_logic_vector(20090, 16),
21238 => conv_std_logic_vector(20172, 16),
21239 => conv_std_logic_vector(20254, 16),
21240 => conv_std_logic_vector(20336, 16),
21241 => conv_std_logic_vector(20418, 16),
21242 => conv_std_logic_vector(20500, 16),
21243 => conv_std_logic_vector(20582, 16),
21244 => conv_std_logic_vector(20664, 16),
21245 => conv_std_logic_vector(20746, 16),
21246 => conv_std_logic_vector(20828, 16),
21247 => conv_std_logic_vector(20910, 16),
21248 => conv_std_logic_vector(0, 16),
21249 => conv_std_logic_vector(83, 16),
21250 => conv_std_logic_vector(166, 16),
21251 => conv_std_logic_vector(249, 16),
21252 => conv_std_logic_vector(332, 16),
21253 => conv_std_logic_vector(415, 16),
21254 => conv_std_logic_vector(498, 16),
21255 => conv_std_logic_vector(581, 16),
21256 => conv_std_logic_vector(664, 16),
21257 => conv_std_logic_vector(747, 16),
21258 => conv_std_logic_vector(830, 16),
21259 => conv_std_logic_vector(913, 16),
21260 => conv_std_logic_vector(996, 16),
21261 => conv_std_logic_vector(1079, 16),
21262 => conv_std_logic_vector(1162, 16),
21263 => conv_std_logic_vector(1245, 16),
21264 => conv_std_logic_vector(1328, 16),
21265 => conv_std_logic_vector(1411, 16),
21266 => conv_std_logic_vector(1494, 16),
21267 => conv_std_logic_vector(1577, 16),
21268 => conv_std_logic_vector(1660, 16),
21269 => conv_std_logic_vector(1743, 16),
21270 => conv_std_logic_vector(1826, 16),
21271 => conv_std_logic_vector(1909, 16),
21272 => conv_std_logic_vector(1992, 16),
21273 => conv_std_logic_vector(2075, 16),
21274 => conv_std_logic_vector(2158, 16),
21275 => conv_std_logic_vector(2241, 16),
21276 => conv_std_logic_vector(2324, 16),
21277 => conv_std_logic_vector(2407, 16),
21278 => conv_std_logic_vector(2490, 16),
21279 => conv_std_logic_vector(2573, 16),
21280 => conv_std_logic_vector(2656, 16),
21281 => conv_std_logic_vector(2739, 16),
21282 => conv_std_logic_vector(2822, 16),
21283 => conv_std_logic_vector(2905, 16),
21284 => conv_std_logic_vector(2988, 16),
21285 => conv_std_logic_vector(3071, 16),
21286 => conv_std_logic_vector(3154, 16),
21287 => conv_std_logic_vector(3237, 16),
21288 => conv_std_logic_vector(3320, 16),
21289 => conv_std_logic_vector(3403, 16),
21290 => conv_std_logic_vector(3486, 16),
21291 => conv_std_logic_vector(3569, 16),
21292 => conv_std_logic_vector(3652, 16),
21293 => conv_std_logic_vector(3735, 16),
21294 => conv_std_logic_vector(3818, 16),
21295 => conv_std_logic_vector(3901, 16),
21296 => conv_std_logic_vector(3984, 16),
21297 => conv_std_logic_vector(4067, 16),
21298 => conv_std_logic_vector(4150, 16),
21299 => conv_std_logic_vector(4233, 16),
21300 => conv_std_logic_vector(4316, 16),
21301 => conv_std_logic_vector(4399, 16),
21302 => conv_std_logic_vector(4482, 16),
21303 => conv_std_logic_vector(4565, 16),
21304 => conv_std_logic_vector(4648, 16),
21305 => conv_std_logic_vector(4731, 16),
21306 => conv_std_logic_vector(4814, 16),
21307 => conv_std_logic_vector(4897, 16),
21308 => conv_std_logic_vector(4980, 16),
21309 => conv_std_logic_vector(5063, 16),
21310 => conv_std_logic_vector(5146, 16),
21311 => conv_std_logic_vector(5229, 16),
21312 => conv_std_logic_vector(5312, 16),
21313 => conv_std_logic_vector(5395, 16),
21314 => conv_std_logic_vector(5478, 16),
21315 => conv_std_logic_vector(5561, 16),
21316 => conv_std_logic_vector(5644, 16),
21317 => conv_std_logic_vector(5727, 16),
21318 => conv_std_logic_vector(5810, 16),
21319 => conv_std_logic_vector(5893, 16),
21320 => conv_std_logic_vector(5976, 16),
21321 => conv_std_logic_vector(6059, 16),
21322 => conv_std_logic_vector(6142, 16),
21323 => conv_std_logic_vector(6225, 16),
21324 => conv_std_logic_vector(6308, 16),
21325 => conv_std_logic_vector(6391, 16),
21326 => conv_std_logic_vector(6474, 16),
21327 => conv_std_logic_vector(6557, 16),
21328 => conv_std_logic_vector(6640, 16),
21329 => conv_std_logic_vector(6723, 16),
21330 => conv_std_logic_vector(6806, 16),
21331 => conv_std_logic_vector(6889, 16),
21332 => conv_std_logic_vector(6972, 16),
21333 => conv_std_logic_vector(7055, 16),
21334 => conv_std_logic_vector(7138, 16),
21335 => conv_std_logic_vector(7221, 16),
21336 => conv_std_logic_vector(7304, 16),
21337 => conv_std_logic_vector(7387, 16),
21338 => conv_std_logic_vector(7470, 16),
21339 => conv_std_logic_vector(7553, 16),
21340 => conv_std_logic_vector(7636, 16),
21341 => conv_std_logic_vector(7719, 16),
21342 => conv_std_logic_vector(7802, 16),
21343 => conv_std_logic_vector(7885, 16),
21344 => conv_std_logic_vector(7968, 16),
21345 => conv_std_logic_vector(8051, 16),
21346 => conv_std_logic_vector(8134, 16),
21347 => conv_std_logic_vector(8217, 16),
21348 => conv_std_logic_vector(8300, 16),
21349 => conv_std_logic_vector(8383, 16),
21350 => conv_std_logic_vector(8466, 16),
21351 => conv_std_logic_vector(8549, 16),
21352 => conv_std_logic_vector(8632, 16),
21353 => conv_std_logic_vector(8715, 16),
21354 => conv_std_logic_vector(8798, 16),
21355 => conv_std_logic_vector(8881, 16),
21356 => conv_std_logic_vector(8964, 16),
21357 => conv_std_logic_vector(9047, 16),
21358 => conv_std_logic_vector(9130, 16),
21359 => conv_std_logic_vector(9213, 16),
21360 => conv_std_logic_vector(9296, 16),
21361 => conv_std_logic_vector(9379, 16),
21362 => conv_std_logic_vector(9462, 16),
21363 => conv_std_logic_vector(9545, 16),
21364 => conv_std_logic_vector(9628, 16),
21365 => conv_std_logic_vector(9711, 16),
21366 => conv_std_logic_vector(9794, 16),
21367 => conv_std_logic_vector(9877, 16),
21368 => conv_std_logic_vector(9960, 16),
21369 => conv_std_logic_vector(10043, 16),
21370 => conv_std_logic_vector(10126, 16),
21371 => conv_std_logic_vector(10209, 16),
21372 => conv_std_logic_vector(10292, 16),
21373 => conv_std_logic_vector(10375, 16),
21374 => conv_std_logic_vector(10458, 16),
21375 => conv_std_logic_vector(10541, 16),
21376 => conv_std_logic_vector(10624, 16),
21377 => conv_std_logic_vector(10707, 16),
21378 => conv_std_logic_vector(10790, 16),
21379 => conv_std_logic_vector(10873, 16),
21380 => conv_std_logic_vector(10956, 16),
21381 => conv_std_logic_vector(11039, 16),
21382 => conv_std_logic_vector(11122, 16),
21383 => conv_std_logic_vector(11205, 16),
21384 => conv_std_logic_vector(11288, 16),
21385 => conv_std_logic_vector(11371, 16),
21386 => conv_std_logic_vector(11454, 16),
21387 => conv_std_logic_vector(11537, 16),
21388 => conv_std_logic_vector(11620, 16),
21389 => conv_std_logic_vector(11703, 16),
21390 => conv_std_logic_vector(11786, 16),
21391 => conv_std_logic_vector(11869, 16),
21392 => conv_std_logic_vector(11952, 16),
21393 => conv_std_logic_vector(12035, 16),
21394 => conv_std_logic_vector(12118, 16),
21395 => conv_std_logic_vector(12201, 16),
21396 => conv_std_logic_vector(12284, 16),
21397 => conv_std_logic_vector(12367, 16),
21398 => conv_std_logic_vector(12450, 16),
21399 => conv_std_logic_vector(12533, 16),
21400 => conv_std_logic_vector(12616, 16),
21401 => conv_std_logic_vector(12699, 16),
21402 => conv_std_logic_vector(12782, 16),
21403 => conv_std_logic_vector(12865, 16),
21404 => conv_std_logic_vector(12948, 16),
21405 => conv_std_logic_vector(13031, 16),
21406 => conv_std_logic_vector(13114, 16),
21407 => conv_std_logic_vector(13197, 16),
21408 => conv_std_logic_vector(13280, 16),
21409 => conv_std_logic_vector(13363, 16),
21410 => conv_std_logic_vector(13446, 16),
21411 => conv_std_logic_vector(13529, 16),
21412 => conv_std_logic_vector(13612, 16),
21413 => conv_std_logic_vector(13695, 16),
21414 => conv_std_logic_vector(13778, 16),
21415 => conv_std_logic_vector(13861, 16),
21416 => conv_std_logic_vector(13944, 16),
21417 => conv_std_logic_vector(14027, 16),
21418 => conv_std_logic_vector(14110, 16),
21419 => conv_std_logic_vector(14193, 16),
21420 => conv_std_logic_vector(14276, 16),
21421 => conv_std_logic_vector(14359, 16),
21422 => conv_std_logic_vector(14442, 16),
21423 => conv_std_logic_vector(14525, 16),
21424 => conv_std_logic_vector(14608, 16),
21425 => conv_std_logic_vector(14691, 16),
21426 => conv_std_logic_vector(14774, 16),
21427 => conv_std_logic_vector(14857, 16),
21428 => conv_std_logic_vector(14940, 16),
21429 => conv_std_logic_vector(15023, 16),
21430 => conv_std_logic_vector(15106, 16),
21431 => conv_std_logic_vector(15189, 16),
21432 => conv_std_logic_vector(15272, 16),
21433 => conv_std_logic_vector(15355, 16),
21434 => conv_std_logic_vector(15438, 16),
21435 => conv_std_logic_vector(15521, 16),
21436 => conv_std_logic_vector(15604, 16),
21437 => conv_std_logic_vector(15687, 16),
21438 => conv_std_logic_vector(15770, 16),
21439 => conv_std_logic_vector(15853, 16),
21440 => conv_std_logic_vector(15936, 16),
21441 => conv_std_logic_vector(16019, 16),
21442 => conv_std_logic_vector(16102, 16),
21443 => conv_std_logic_vector(16185, 16),
21444 => conv_std_logic_vector(16268, 16),
21445 => conv_std_logic_vector(16351, 16),
21446 => conv_std_logic_vector(16434, 16),
21447 => conv_std_logic_vector(16517, 16),
21448 => conv_std_logic_vector(16600, 16),
21449 => conv_std_logic_vector(16683, 16),
21450 => conv_std_logic_vector(16766, 16),
21451 => conv_std_logic_vector(16849, 16),
21452 => conv_std_logic_vector(16932, 16),
21453 => conv_std_logic_vector(17015, 16),
21454 => conv_std_logic_vector(17098, 16),
21455 => conv_std_logic_vector(17181, 16),
21456 => conv_std_logic_vector(17264, 16),
21457 => conv_std_logic_vector(17347, 16),
21458 => conv_std_logic_vector(17430, 16),
21459 => conv_std_logic_vector(17513, 16),
21460 => conv_std_logic_vector(17596, 16),
21461 => conv_std_logic_vector(17679, 16),
21462 => conv_std_logic_vector(17762, 16),
21463 => conv_std_logic_vector(17845, 16),
21464 => conv_std_logic_vector(17928, 16),
21465 => conv_std_logic_vector(18011, 16),
21466 => conv_std_logic_vector(18094, 16),
21467 => conv_std_logic_vector(18177, 16),
21468 => conv_std_logic_vector(18260, 16),
21469 => conv_std_logic_vector(18343, 16),
21470 => conv_std_logic_vector(18426, 16),
21471 => conv_std_logic_vector(18509, 16),
21472 => conv_std_logic_vector(18592, 16),
21473 => conv_std_logic_vector(18675, 16),
21474 => conv_std_logic_vector(18758, 16),
21475 => conv_std_logic_vector(18841, 16),
21476 => conv_std_logic_vector(18924, 16),
21477 => conv_std_logic_vector(19007, 16),
21478 => conv_std_logic_vector(19090, 16),
21479 => conv_std_logic_vector(19173, 16),
21480 => conv_std_logic_vector(19256, 16),
21481 => conv_std_logic_vector(19339, 16),
21482 => conv_std_logic_vector(19422, 16),
21483 => conv_std_logic_vector(19505, 16),
21484 => conv_std_logic_vector(19588, 16),
21485 => conv_std_logic_vector(19671, 16),
21486 => conv_std_logic_vector(19754, 16),
21487 => conv_std_logic_vector(19837, 16),
21488 => conv_std_logic_vector(19920, 16),
21489 => conv_std_logic_vector(20003, 16),
21490 => conv_std_logic_vector(20086, 16),
21491 => conv_std_logic_vector(20169, 16),
21492 => conv_std_logic_vector(20252, 16),
21493 => conv_std_logic_vector(20335, 16),
21494 => conv_std_logic_vector(20418, 16),
21495 => conv_std_logic_vector(20501, 16),
21496 => conv_std_logic_vector(20584, 16),
21497 => conv_std_logic_vector(20667, 16),
21498 => conv_std_logic_vector(20750, 16),
21499 => conv_std_logic_vector(20833, 16),
21500 => conv_std_logic_vector(20916, 16),
21501 => conv_std_logic_vector(20999, 16),
21502 => conv_std_logic_vector(21082, 16),
21503 => conv_std_logic_vector(21165, 16),
21504 => conv_std_logic_vector(0, 16),
21505 => conv_std_logic_vector(84, 16),
21506 => conv_std_logic_vector(168, 16),
21507 => conv_std_logic_vector(252, 16),
21508 => conv_std_logic_vector(336, 16),
21509 => conv_std_logic_vector(420, 16),
21510 => conv_std_logic_vector(504, 16),
21511 => conv_std_logic_vector(588, 16),
21512 => conv_std_logic_vector(672, 16),
21513 => conv_std_logic_vector(756, 16),
21514 => conv_std_logic_vector(840, 16),
21515 => conv_std_logic_vector(924, 16),
21516 => conv_std_logic_vector(1008, 16),
21517 => conv_std_logic_vector(1092, 16),
21518 => conv_std_logic_vector(1176, 16),
21519 => conv_std_logic_vector(1260, 16),
21520 => conv_std_logic_vector(1344, 16),
21521 => conv_std_logic_vector(1428, 16),
21522 => conv_std_logic_vector(1512, 16),
21523 => conv_std_logic_vector(1596, 16),
21524 => conv_std_logic_vector(1680, 16),
21525 => conv_std_logic_vector(1764, 16),
21526 => conv_std_logic_vector(1848, 16),
21527 => conv_std_logic_vector(1932, 16),
21528 => conv_std_logic_vector(2016, 16),
21529 => conv_std_logic_vector(2100, 16),
21530 => conv_std_logic_vector(2184, 16),
21531 => conv_std_logic_vector(2268, 16),
21532 => conv_std_logic_vector(2352, 16),
21533 => conv_std_logic_vector(2436, 16),
21534 => conv_std_logic_vector(2520, 16),
21535 => conv_std_logic_vector(2604, 16),
21536 => conv_std_logic_vector(2688, 16),
21537 => conv_std_logic_vector(2772, 16),
21538 => conv_std_logic_vector(2856, 16),
21539 => conv_std_logic_vector(2940, 16),
21540 => conv_std_logic_vector(3024, 16),
21541 => conv_std_logic_vector(3108, 16),
21542 => conv_std_logic_vector(3192, 16),
21543 => conv_std_logic_vector(3276, 16),
21544 => conv_std_logic_vector(3360, 16),
21545 => conv_std_logic_vector(3444, 16),
21546 => conv_std_logic_vector(3528, 16),
21547 => conv_std_logic_vector(3612, 16),
21548 => conv_std_logic_vector(3696, 16),
21549 => conv_std_logic_vector(3780, 16),
21550 => conv_std_logic_vector(3864, 16),
21551 => conv_std_logic_vector(3948, 16),
21552 => conv_std_logic_vector(4032, 16),
21553 => conv_std_logic_vector(4116, 16),
21554 => conv_std_logic_vector(4200, 16),
21555 => conv_std_logic_vector(4284, 16),
21556 => conv_std_logic_vector(4368, 16),
21557 => conv_std_logic_vector(4452, 16),
21558 => conv_std_logic_vector(4536, 16),
21559 => conv_std_logic_vector(4620, 16),
21560 => conv_std_logic_vector(4704, 16),
21561 => conv_std_logic_vector(4788, 16),
21562 => conv_std_logic_vector(4872, 16),
21563 => conv_std_logic_vector(4956, 16),
21564 => conv_std_logic_vector(5040, 16),
21565 => conv_std_logic_vector(5124, 16),
21566 => conv_std_logic_vector(5208, 16),
21567 => conv_std_logic_vector(5292, 16),
21568 => conv_std_logic_vector(5376, 16),
21569 => conv_std_logic_vector(5460, 16),
21570 => conv_std_logic_vector(5544, 16),
21571 => conv_std_logic_vector(5628, 16),
21572 => conv_std_logic_vector(5712, 16),
21573 => conv_std_logic_vector(5796, 16),
21574 => conv_std_logic_vector(5880, 16),
21575 => conv_std_logic_vector(5964, 16),
21576 => conv_std_logic_vector(6048, 16),
21577 => conv_std_logic_vector(6132, 16),
21578 => conv_std_logic_vector(6216, 16),
21579 => conv_std_logic_vector(6300, 16),
21580 => conv_std_logic_vector(6384, 16),
21581 => conv_std_logic_vector(6468, 16),
21582 => conv_std_logic_vector(6552, 16),
21583 => conv_std_logic_vector(6636, 16),
21584 => conv_std_logic_vector(6720, 16),
21585 => conv_std_logic_vector(6804, 16),
21586 => conv_std_logic_vector(6888, 16),
21587 => conv_std_logic_vector(6972, 16),
21588 => conv_std_logic_vector(7056, 16),
21589 => conv_std_logic_vector(7140, 16),
21590 => conv_std_logic_vector(7224, 16),
21591 => conv_std_logic_vector(7308, 16),
21592 => conv_std_logic_vector(7392, 16),
21593 => conv_std_logic_vector(7476, 16),
21594 => conv_std_logic_vector(7560, 16),
21595 => conv_std_logic_vector(7644, 16),
21596 => conv_std_logic_vector(7728, 16),
21597 => conv_std_logic_vector(7812, 16),
21598 => conv_std_logic_vector(7896, 16),
21599 => conv_std_logic_vector(7980, 16),
21600 => conv_std_logic_vector(8064, 16),
21601 => conv_std_logic_vector(8148, 16),
21602 => conv_std_logic_vector(8232, 16),
21603 => conv_std_logic_vector(8316, 16),
21604 => conv_std_logic_vector(8400, 16),
21605 => conv_std_logic_vector(8484, 16),
21606 => conv_std_logic_vector(8568, 16),
21607 => conv_std_logic_vector(8652, 16),
21608 => conv_std_logic_vector(8736, 16),
21609 => conv_std_logic_vector(8820, 16),
21610 => conv_std_logic_vector(8904, 16),
21611 => conv_std_logic_vector(8988, 16),
21612 => conv_std_logic_vector(9072, 16),
21613 => conv_std_logic_vector(9156, 16),
21614 => conv_std_logic_vector(9240, 16),
21615 => conv_std_logic_vector(9324, 16),
21616 => conv_std_logic_vector(9408, 16),
21617 => conv_std_logic_vector(9492, 16),
21618 => conv_std_logic_vector(9576, 16),
21619 => conv_std_logic_vector(9660, 16),
21620 => conv_std_logic_vector(9744, 16),
21621 => conv_std_logic_vector(9828, 16),
21622 => conv_std_logic_vector(9912, 16),
21623 => conv_std_logic_vector(9996, 16),
21624 => conv_std_logic_vector(10080, 16),
21625 => conv_std_logic_vector(10164, 16),
21626 => conv_std_logic_vector(10248, 16),
21627 => conv_std_logic_vector(10332, 16),
21628 => conv_std_logic_vector(10416, 16),
21629 => conv_std_logic_vector(10500, 16),
21630 => conv_std_logic_vector(10584, 16),
21631 => conv_std_logic_vector(10668, 16),
21632 => conv_std_logic_vector(10752, 16),
21633 => conv_std_logic_vector(10836, 16),
21634 => conv_std_logic_vector(10920, 16),
21635 => conv_std_logic_vector(11004, 16),
21636 => conv_std_logic_vector(11088, 16),
21637 => conv_std_logic_vector(11172, 16),
21638 => conv_std_logic_vector(11256, 16),
21639 => conv_std_logic_vector(11340, 16),
21640 => conv_std_logic_vector(11424, 16),
21641 => conv_std_logic_vector(11508, 16),
21642 => conv_std_logic_vector(11592, 16),
21643 => conv_std_logic_vector(11676, 16),
21644 => conv_std_logic_vector(11760, 16),
21645 => conv_std_logic_vector(11844, 16),
21646 => conv_std_logic_vector(11928, 16),
21647 => conv_std_logic_vector(12012, 16),
21648 => conv_std_logic_vector(12096, 16),
21649 => conv_std_logic_vector(12180, 16),
21650 => conv_std_logic_vector(12264, 16),
21651 => conv_std_logic_vector(12348, 16),
21652 => conv_std_logic_vector(12432, 16),
21653 => conv_std_logic_vector(12516, 16),
21654 => conv_std_logic_vector(12600, 16),
21655 => conv_std_logic_vector(12684, 16),
21656 => conv_std_logic_vector(12768, 16),
21657 => conv_std_logic_vector(12852, 16),
21658 => conv_std_logic_vector(12936, 16),
21659 => conv_std_logic_vector(13020, 16),
21660 => conv_std_logic_vector(13104, 16),
21661 => conv_std_logic_vector(13188, 16),
21662 => conv_std_logic_vector(13272, 16),
21663 => conv_std_logic_vector(13356, 16),
21664 => conv_std_logic_vector(13440, 16),
21665 => conv_std_logic_vector(13524, 16),
21666 => conv_std_logic_vector(13608, 16),
21667 => conv_std_logic_vector(13692, 16),
21668 => conv_std_logic_vector(13776, 16),
21669 => conv_std_logic_vector(13860, 16),
21670 => conv_std_logic_vector(13944, 16),
21671 => conv_std_logic_vector(14028, 16),
21672 => conv_std_logic_vector(14112, 16),
21673 => conv_std_logic_vector(14196, 16),
21674 => conv_std_logic_vector(14280, 16),
21675 => conv_std_logic_vector(14364, 16),
21676 => conv_std_logic_vector(14448, 16),
21677 => conv_std_logic_vector(14532, 16),
21678 => conv_std_logic_vector(14616, 16),
21679 => conv_std_logic_vector(14700, 16),
21680 => conv_std_logic_vector(14784, 16),
21681 => conv_std_logic_vector(14868, 16),
21682 => conv_std_logic_vector(14952, 16),
21683 => conv_std_logic_vector(15036, 16),
21684 => conv_std_logic_vector(15120, 16),
21685 => conv_std_logic_vector(15204, 16),
21686 => conv_std_logic_vector(15288, 16),
21687 => conv_std_logic_vector(15372, 16),
21688 => conv_std_logic_vector(15456, 16),
21689 => conv_std_logic_vector(15540, 16),
21690 => conv_std_logic_vector(15624, 16),
21691 => conv_std_logic_vector(15708, 16),
21692 => conv_std_logic_vector(15792, 16),
21693 => conv_std_logic_vector(15876, 16),
21694 => conv_std_logic_vector(15960, 16),
21695 => conv_std_logic_vector(16044, 16),
21696 => conv_std_logic_vector(16128, 16),
21697 => conv_std_logic_vector(16212, 16),
21698 => conv_std_logic_vector(16296, 16),
21699 => conv_std_logic_vector(16380, 16),
21700 => conv_std_logic_vector(16464, 16),
21701 => conv_std_logic_vector(16548, 16),
21702 => conv_std_logic_vector(16632, 16),
21703 => conv_std_logic_vector(16716, 16),
21704 => conv_std_logic_vector(16800, 16),
21705 => conv_std_logic_vector(16884, 16),
21706 => conv_std_logic_vector(16968, 16),
21707 => conv_std_logic_vector(17052, 16),
21708 => conv_std_logic_vector(17136, 16),
21709 => conv_std_logic_vector(17220, 16),
21710 => conv_std_logic_vector(17304, 16),
21711 => conv_std_logic_vector(17388, 16),
21712 => conv_std_logic_vector(17472, 16),
21713 => conv_std_logic_vector(17556, 16),
21714 => conv_std_logic_vector(17640, 16),
21715 => conv_std_logic_vector(17724, 16),
21716 => conv_std_logic_vector(17808, 16),
21717 => conv_std_logic_vector(17892, 16),
21718 => conv_std_logic_vector(17976, 16),
21719 => conv_std_logic_vector(18060, 16),
21720 => conv_std_logic_vector(18144, 16),
21721 => conv_std_logic_vector(18228, 16),
21722 => conv_std_logic_vector(18312, 16),
21723 => conv_std_logic_vector(18396, 16),
21724 => conv_std_logic_vector(18480, 16),
21725 => conv_std_logic_vector(18564, 16),
21726 => conv_std_logic_vector(18648, 16),
21727 => conv_std_logic_vector(18732, 16),
21728 => conv_std_logic_vector(18816, 16),
21729 => conv_std_logic_vector(18900, 16),
21730 => conv_std_logic_vector(18984, 16),
21731 => conv_std_logic_vector(19068, 16),
21732 => conv_std_logic_vector(19152, 16),
21733 => conv_std_logic_vector(19236, 16),
21734 => conv_std_logic_vector(19320, 16),
21735 => conv_std_logic_vector(19404, 16),
21736 => conv_std_logic_vector(19488, 16),
21737 => conv_std_logic_vector(19572, 16),
21738 => conv_std_logic_vector(19656, 16),
21739 => conv_std_logic_vector(19740, 16),
21740 => conv_std_logic_vector(19824, 16),
21741 => conv_std_logic_vector(19908, 16),
21742 => conv_std_logic_vector(19992, 16),
21743 => conv_std_logic_vector(20076, 16),
21744 => conv_std_logic_vector(20160, 16),
21745 => conv_std_logic_vector(20244, 16),
21746 => conv_std_logic_vector(20328, 16),
21747 => conv_std_logic_vector(20412, 16),
21748 => conv_std_logic_vector(20496, 16),
21749 => conv_std_logic_vector(20580, 16),
21750 => conv_std_logic_vector(20664, 16),
21751 => conv_std_logic_vector(20748, 16),
21752 => conv_std_logic_vector(20832, 16),
21753 => conv_std_logic_vector(20916, 16),
21754 => conv_std_logic_vector(21000, 16),
21755 => conv_std_logic_vector(21084, 16),
21756 => conv_std_logic_vector(21168, 16),
21757 => conv_std_logic_vector(21252, 16),
21758 => conv_std_logic_vector(21336, 16),
21759 => conv_std_logic_vector(21420, 16),
21760 => conv_std_logic_vector(0, 16),
21761 => conv_std_logic_vector(85, 16),
21762 => conv_std_logic_vector(170, 16),
21763 => conv_std_logic_vector(255, 16),
21764 => conv_std_logic_vector(340, 16),
21765 => conv_std_logic_vector(425, 16),
21766 => conv_std_logic_vector(510, 16),
21767 => conv_std_logic_vector(595, 16),
21768 => conv_std_logic_vector(680, 16),
21769 => conv_std_logic_vector(765, 16),
21770 => conv_std_logic_vector(850, 16),
21771 => conv_std_logic_vector(935, 16),
21772 => conv_std_logic_vector(1020, 16),
21773 => conv_std_logic_vector(1105, 16),
21774 => conv_std_logic_vector(1190, 16),
21775 => conv_std_logic_vector(1275, 16),
21776 => conv_std_logic_vector(1360, 16),
21777 => conv_std_logic_vector(1445, 16),
21778 => conv_std_logic_vector(1530, 16),
21779 => conv_std_logic_vector(1615, 16),
21780 => conv_std_logic_vector(1700, 16),
21781 => conv_std_logic_vector(1785, 16),
21782 => conv_std_logic_vector(1870, 16),
21783 => conv_std_logic_vector(1955, 16),
21784 => conv_std_logic_vector(2040, 16),
21785 => conv_std_logic_vector(2125, 16),
21786 => conv_std_logic_vector(2210, 16),
21787 => conv_std_logic_vector(2295, 16),
21788 => conv_std_logic_vector(2380, 16),
21789 => conv_std_logic_vector(2465, 16),
21790 => conv_std_logic_vector(2550, 16),
21791 => conv_std_logic_vector(2635, 16),
21792 => conv_std_logic_vector(2720, 16),
21793 => conv_std_logic_vector(2805, 16),
21794 => conv_std_logic_vector(2890, 16),
21795 => conv_std_logic_vector(2975, 16),
21796 => conv_std_logic_vector(3060, 16),
21797 => conv_std_logic_vector(3145, 16),
21798 => conv_std_logic_vector(3230, 16),
21799 => conv_std_logic_vector(3315, 16),
21800 => conv_std_logic_vector(3400, 16),
21801 => conv_std_logic_vector(3485, 16),
21802 => conv_std_logic_vector(3570, 16),
21803 => conv_std_logic_vector(3655, 16),
21804 => conv_std_logic_vector(3740, 16),
21805 => conv_std_logic_vector(3825, 16),
21806 => conv_std_logic_vector(3910, 16),
21807 => conv_std_logic_vector(3995, 16),
21808 => conv_std_logic_vector(4080, 16),
21809 => conv_std_logic_vector(4165, 16),
21810 => conv_std_logic_vector(4250, 16),
21811 => conv_std_logic_vector(4335, 16),
21812 => conv_std_logic_vector(4420, 16),
21813 => conv_std_logic_vector(4505, 16),
21814 => conv_std_logic_vector(4590, 16),
21815 => conv_std_logic_vector(4675, 16),
21816 => conv_std_logic_vector(4760, 16),
21817 => conv_std_logic_vector(4845, 16),
21818 => conv_std_logic_vector(4930, 16),
21819 => conv_std_logic_vector(5015, 16),
21820 => conv_std_logic_vector(5100, 16),
21821 => conv_std_logic_vector(5185, 16),
21822 => conv_std_logic_vector(5270, 16),
21823 => conv_std_logic_vector(5355, 16),
21824 => conv_std_logic_vector(5440, 16),
21825 => conv_std_logic_vector(5525, 16),
21826 => conv_std_logic_vector(5610, 16),
21827 => conv_std_logic_vector(5695, 16),
21828 => conv_std_logic_vector(5780, 16),
21829 => conv_std_logic_vector(5865, 16),
21830 => conv_std_logic_vector(5950, 16),
21831 => conv_std_logic_vector(6035, 16),
21832 => conv_std_logic_vector(6120, 16),
21833 => conv_std_logic_vector(6205, 16),
21834 => conv_std_logic_vector(6290, 16),
21835 => conv_std_logic_vector(6375, 16),
21836 => conv_std_logic_vector(6460, 16),
21837 => conv_std_logic_vector(6545, 16),
21838 => conv_std_logic_vector(6630, 16),
21839 => conv_std_logic_vector(6715, 16),
21840 => conv_std_logic_vector(6800, 16),
21841 => conv_std_logic_vector(6885, 16),
21842 => conv_std_logic_vector(6970, 16),
21843 => conv_std_logic_vector(7055, 16),
21844 => conv_std_logic_vector(7140, 16),
21845 => conv_std_logic_vector(7225, 16),
21846 => conv_std_logic_vector(7310, 16),
21847 => conv_std_logic_vector(7395, 16),
21848 => conv_std_logic_vector(7480, 16),
21849 => conv_std_logic_vector(7565, 16),
21850 => conv_std_logic_vector(7650, 16),
21851 => conv_std_logic_vector(7735, 16),
21852 => conv_std_logic_vector(7820, 16),
21853 => conv_std_logic_vector(7905, 16),
21854 => conv_std_logic_vector(7990, 16),
21855 => conv_std_logic_vector(8075, 16),
21856 => conv_std_logic_vector(8160, 16),
21857 => conv_std_logic_vector(8245, 16),
21858 => conv_std_logic_vector(8330, 16),
21859 => conv_std_logic_vector(8415, 16),
21860 => conv_std_logic_vector(8500, 16),
21861 => conv_std_logic_vector(8585, 16),
21862 => conv_std_logic_vector(8670, 16),
21863 => conv_std_logic_vector(8755, 16),
21864 => conv_std_logic_vector(8840, 16),
21865 => conv_std_logic_vector(8925, 16),
21866 => conv_std_logic_vector(9010, 16),
21867 => conv_std_logic_vector(9095, 16),
21868 => conv_std_logic_vector(9180, 16),
21869 => conv_std_logic_vector(9265, 16),
21870 => conv_std_logic_vector(9350, 16),
21871 => conv_std_logic_vector(9435, 16),
21872 => conv_std_logic_vector(9520, 16),
21873 => conv_std_logic_vector(9605, 16),
21874 => conv_std_logic_vector(9690, 16),
21875 => conv_std_logic_vector(9775, 16),
21876 => conv_std_logic_vector(9860, 16),
21877 => conv_std_logic_vector(9945, 16),
21878 => conv_std_logic_vector(10030, 16),
21879 => conv_std_logic_vector(10115, 16),
21880 => conv_std_logic_vector(10200, 16),
21881 => conv_std_logic_vector(10285, 16),
21882 => conv_std_logic_vector(10370, 16),
21883 => conv_std_logic_vector(10455, 16),
21884 => conv_std_logic_vector(10540, 16),
21885 => conv_std_logic_vector(10625, 16),
21886 => conv_std_logic_vector(10710, 16),
21887 => conv_std_logic_vector(10795, 16),
21888 => conv_std_logic_vector(10880, 16),
21889 => conv_std_logic_vector(10965, 16),
21890 => conv_std_logic_vector(11050, 16),
21891 => conv_std_logic_vector(11135, 16),
21892 => conv_std_logic_vector(11220, 16),
21893 => conv_std_logic_vector(11305, 16),
21894 => conv_std_logic_vector(11390, 16),
21895 => conv_std_logic_vector(11475, 16),
21896 => conv_std_logic_vector(11560, 16),
21897 => conv_std_logic_vector(11645, 16),
21898 => conv_std_logic_vector(11730, 16),
21899 => conv_std_logic_vector(11815, 16),
21900 => conv_std_logic_vector(11900, 16),
21901 => conv_std_logic_vector(11985, 16),
21902 => conv_std_logic_vector(12070, 16),
21903 => conv_std_logic_vector(12155, 16),
21904 => conv_std_logic_vector(12240, 16),
21905 => conv_std_logic_vector(12325, 16),
21906 => conv_std_logic_vector(12410, 16),
21907 => conv_std_logic_vector(12495, 16),
21908 => conv_std_logic_vector(12580, 16),
21909 => conv_std_logic_vector(12665, 16),
21910 => conv_std_logic_vector(12750, 16),
21911 => conv_std_logic_vector(12835, 16),
21912 => conv_std_logic_vector(12920, 16),
21913 => conv_std_logic_vector(13005, 16),
21914 => conv_std_logic_vector(13090, 16),
21915 => conv_std_logic_vector(13175, 16),
21916 => conv_std_logic_vector(13260, 16),
21917 => conv_std_logic_vector(13345, 16),
21918 => conv_std_logic_vector(13430, 16),
21919 => conv_std_logic_vector(13515, 16),
21920 => conv_std_logic_vector(13600, 16),
21921 => conv_std_logic_vector(13685, 16),
21922 => conv_std_logic_vector(13770, 16),
21923 => conv_std_logic_vector(13855, 16),
21924 => conv_std_logic_vector(13940, 16),
21925 => conv_std_logic_vector(14025, 16),
21926 => conv_std_logic_vector(14110, 16),
21927 => conv_std_logic_vector(14195, 16),
21928 => conv_std_logic_vector(14280, 16),
21929 => conv_std_logic_vector(14365, 16),
21930 => conv_std_logic_vector(14450, 16),
21931 => conv_std_logic_vector(14535, 16),
21932 => conv_std_logic_vector(14620, 16),
21933 => conv_std_logic_vector(14705, 16),
21934 => conv_std_logic_vector(14790, 16),
21935 => conv_std_logic_vector(14875, 16),
21936 => conv_std_logic_vector(14960, 16),
21937 => conv_std_logic_vector(15045, 16),
21938 => conv_std_logic_vector(15130, 16),
21939 => conv_std_logic_vector(15215, 16),
21940 => conv_std_logic_vector(15300, 16),
21941 => conv_std_logic_vector(15385, 16),
21942 => conv_std_logic_vector(15470, 16),
21943 => conv_std_logic_vector(15555, 16),
21944 => conv_std_logic_vector(15640, 16),
21945 => conv_std_logic_vector(15725, 16),
21946 => conv_std_logic_vector(15810, 16),
21947 => conv_std_logic_vector(15895, 16),
21948 => conv_std_logic_vector(15980, 16),
21949 => conv_std_logic_vector(16065, 16),
21950 => conv_std_logic_vector(16150, 16),
21951 => conv_std_logic_vector(16235, 16),
21952 => conv_std_logic_vector(16320, 16),
21953 => conv_std_logic_vector(16405, 16),
21954 => conv_std_logic_vector(16490, 16),
21955 => conv_std_logic_vector(16575, 16),
21956 => conv_std_logic_vector(16660, 16),
21957 => conv_std_logic_vector(16745, 16),
21958 => conv_std_logic_vector(16830, 16),
21959 => conv_std_logic_vector(16915, 16),
21960 => conv_std_logic_vector(17000, 16),
21961 => conv_std_logic_vector(17085, 16),
21962 => conv_std_logic_vector(17170, 16),
21963 => conv_std_logic_vector(17255, 16),
21964 => conv_std_logic_vector(17340, 16),
21965 => conv_std_logic_vector(17425, 16),
21966 => conv_std_logic_vector(17510, 16),
21967 => conv_std_logic_vector(17595, 16),
21968 => conv_std_logic_vector(17680, 16),
21969 => conv_std_logic_vector(17765, 16),
21970 => conv_std_logic_vector(17850, 16),
21971 => conv_std_logic_vector(17935, 16),
21972 => conv_std_logic_vector(18020, 16),
21973 => conv_std_logic_vector(18105, 16),
21974 => conv_std_logic_vector(18190, 16),
21975 => conv_std_logic_vector(18275, 16),
21976 => conv_std_logic_vector(18360, 16),
21977 => conv_std_logic_vector(18445, 16),
21978 => conv_std_logic_vector(18530, 16),
21979 => conv_std_logic_vector(18615, 16),
21980 => conv_std_logic_vector(18700, 16),
21981 => conv_std_logic_vector(18785, 16),
21982 => conv_std_logic_vector(18870, 16),
21983 => conv_std_logic_vector(18955, 16),
21984 => conv_std_logic_vector(19040, 16),
21985 => conv_std_logic_vector(19125, 16),
21986 => conv_std_logic_vector(19210, 16),
21987 => conv_std_logic_vector(19295, 16),
21988 => conv_std_logic_vector(19380, 16),
21989 => conv_std_logic_vector(19465, 16),
21990 => conv_std_logic_vector(19550, 16),
21991 => conv_std_logic_vector(19635, 16),
21992 => conv_std_logic_vector(19720, 16),
21993 => conv_std_logic_vector(19805, 16),
21994 => conv_std_logic_vector(19890, 16),
21995 => conv_std_logic_vector(19975, 16),
21996 => conv_std_logic_vector(20060, 16),
21997 => conv_std_logic_vector(20145, 16),
21998 => conv_std_logic_vector(20230, 16),
21999 => conv_std_logic_vector(20315, 16),
22000 => conv_std_logic_vector(20400, 16),
22001 => conv_std_logic_vector(20485, 16),
22002 => conv_std_logic_vector(20570, 16),
22003 => conv_std_logic_vector(20655, 16),
22004 => conv_std_logic_vector(20740, 16),
22005 => conv_std_logic_vector(20825, 16),
22006 => conv_std_logic_vector(20910, 16),
22007 => conv_std_logic_vector(20995, 16),
22008 => conv_std_logic_vector(21080, 16),
22009 => conv_std_logic_vector(21165, 16),
22010 => conv_std_logic_vector(21250, 16),
22011 => conv_std_logic_vector(21335, 16),
22012 => conv_std_logic_vector(21420, 16),
22013 => conv_std_logic_vector(21505, 16),
22014 => conv_std_logic_vector(21590, 16),
22015 => conv_std_logic_vector(21675, 16),
22016 => conv_std_logic_vector(0, 16),
22017 => conv_std_logic_vector(86, 16),
22018 => conv_std_logic_vector(172, 16),
22019 => conv_std_logic_vector(258, 16),
22020 => conv_std_logic_vector(344, 16),
22021 => conv_std_logic_vector(430, 16),
22022 => conv_std_logic_vector(516, 16),
22023 => conv_std_logic_vector(602, 16),
22024 => conv_std_logic_vector(688, 16),
22025 => conv_std_logic_vector(774, 16),
22026 => conv_std_logic_vector(860, 16),
22027 => conv_std_logic_vector(946, 16),
22028 => conv_std_logic_vector(1032, 16),
22029 => conv_std_logic_vector(1118, 16),
22030 => conv_std_logic_vector(1204, 16),
22031 => conv_std_logic_vector(1290, 16),
22032 => conv_std_logic_vector(1376, 16),
22033 => conv_std_logic_vector(1462, 16),
22034 => conv_std_logic_vector(1548, 16),
22035 => conv_std_logic_vector(1634, 16),
22036 => conv_std_logic_vector(1720, 16),
22037 => conv_std_logic_vector(1806, 16),
22038 => conv_std_logic_vector(1892, 16),
22039 => conv_std_logic_vector(1978, 16),
22040 => conv_std_logic_vector(2064, 16),
22041 => conv_std_logic_vector(2150, 16),
22042 => conv_std_logic_vector(2236, 16),
22043 => conv_std_logic_vector(2322, 16),
22044 => conv_std_logic_vector(2408, 16),
22045 => conv_std_logic_vector(2494, 16),
22046 => conv_std_logic_vector(2580, 16),
22047 => conv_std_logic_vector(2666, 16),
22048 => conv_std_logic_vector(2752, 16),
22049 => conv_std_logic_vector(2838, 16),
22050 => conv_std_logic_vector(2924, 16),
22051 => conv_std_logic_vector(3010, 16),
22052 => conv_std_logic_vector(3096, 16),
22053 => conv_std_logic_vector(3182, 16),
22054 => conv_std_logic_vector(3268, 16),
22055 => conv_std_logic_vector(3354, 16),
22056 => conv_std_logic_vector(3440, 16),
22057 => conv_std_logic_vector(3526, 16),
22058 => conv_std_logic_vector(3612, 16),
22059 => conv_std_logic_vector(3698, 16),
22060 => conv_std_logic_vector(3784, 16),
22061 => conv_std_logic_vector(3870, 16),
22062 => conv_std_logic_vector(3956, 16),
22063 => conv_std_logic_vector(4042, 16),
22064 => conv_std_logic_vector(4128, 16),
22065 => conv_std_logic_vector(4214, 16),
22066 => conv_std_logic_vector(4300, 16),
22067 => conv_std_logic_vector(4386, 16),
22068 => conv_std_logic_vector(4472, 16),
22069 => conv_std_logic_vector(4558, 16),
22070 => conv_std_logic_vector(4644, 16),
22071 => conv_std_logic_vector(4730, 16),
22072 => conv_std_logic_vector(4816, 16),
22073 => conv_std_logic_vector(4902, 16),
22074 => conv_std_logic_vector(4988, 16),
22075 => conv_std_logic_vector(5074, 16),
22076 => conv_std_logic_vector(5160, 16),
22077 => conv_std_logic_vector(5246, 16),
22078 => conv_std_logic_vector(5332, 16),
22079 => conv_std_logic_vector(5418, 16),
22080 => conv_std_logic_vector(5504, 16),
22081 => conv_std_logic_vector(5590, 16),
22082 => conv_std_logic_vector(5676, 16),
22083 => conv_std_logic_vector(5762, 16),
22084 => conv_std_logic_vector(5848, 16),
22085 => conv_std_logic_vector(5934, 16),
22086 => conv_std_logic_vector(6020, 16),
22087 => conv_std_logic_vector(6106, 16),
22088 => conv_std_logic_vector(6192, 16),
22089 => conv_std_logic_vector(6278, 16),
22090 => conv_std_logic_vector(6364, 16),
22091 => conv_std_logic_vector(6450, 16),
22092 => conv_std_logic_vector(6536, 16),
22093 => conv_std_logic_vector(6622, 16),
22094 => conv_std_logic_vector(6708, 16),
22095 => conv_std_logic_vector(6794, 16),
22096 => conv_std_logic_vector(6880, 16),
22097 => conv_std_logic_vector(6966, 16),
22098 => conv_std_logic_vector(7052, 16),
22099 => conv_std_logic_vector(7138, 16),
22100 => conv_std_logic_vector(7224, 16),
22101 => conv_std_logic_vector(7310, 16),
22102 => conv_std_logic_vector(7396, 16),
22103 => conv_std_logic_vector(7482, 16),
22104 => conv_std_logic_vector(7568, 16),
22105 => conv_std_logic_vector(7654, 16),
22106 => conv_std_logic_vector(7740, 16),
22107 => conv_std_logic_vector(7826, 16),
22108 => conv_std_logic_vector(7912, 16),
22109 => conv_std_logic_vector(7998, 16),
22110 => conv_std_logic_vector(8084, 16),
22111 => conv_std_logic_vector(8170, 16),
22112 => conv_std_logic_vector(8256, 16),
22113 => conv_std_logic_vector(8342, 16),
22114 => conv_std_logic_vector(8428, 16),
22115 => conv_std_logic_vector(8514, 16),
22116 => conv_std_logic_vector(8600, 16),
22117 => conv_std_logic_vector(8686, 16),
22118 => conv_std_logic_vector(8772, 16),
22119 => conv_std_logic_vector(8858, 16),
22120 => conv_std_logic_vector(8944, 16),
22121 => conv_std_logic_vector(9030, 16),
22122 => conv_std_logic_vector(9116, 16),
22123 => conv_std_logic_vector(9202, 16),
22124 => conv_std_logic_vector(9288, 16),
22125 => conv_std_logic_vector(9374, 16),
22126 => conv_std_logic_vector(9460, 16),
22127 => conv_std_logic_vector(9546, 16),
22128 => conv_std_logic_vector(9632, 16),
22129 => conv_std_logic_vector(9718, 16),
22130 => conv_std_logic_vector(9804, 16),
22131 => conv_std_logic_vector(9890, 16),
22132 => conv_std_logic_vector(9976, 16),
22133 => conv_std_logic_vector(10062, 16),
22134 => conv_std_logic_vector(10148, 16),
22135 => conv_std_logic_vector(10234, 16),
22136 => conv_std_logic_vector(10320, 16),
22137 => conv_std_logic_vector(10406, 16),
22138 => conv_std_logic_vector(10492, 16),
22139 => conv_std_logic_vector(10578, 16),
22140 => conv_std_logic_vector(10664, 16),
22141 => conv_std_logic_vector(10750, 16),
22142 => conv_std_logic_vector(10836, 16),
22143 => conv_std_logic_vector(10922, 16),
22144 => conv_std_logic_vector(11008, 16),
22145 => conv_std_logic_vector(11094, 16),
22146 => conv_std_logic_vector(11180, 16),
22147 => conv_std_logic_vector(11266, 16),
22148 => conv_std_logic_vector(11352, 16),
22149 => conv_std_logic_vector(11438, 16),
22150 => conv_std_logic_vector(11524, 16),
22151 => conv_std_logic_vector(11610, 16),
22152 => conv_std_logic_vector(11696, 16),
22153 => conv_std_logic_vector(11782, 16),
22154 => conv_std_logic_vector(11868, 16),
22155 => conv_std_logic_vector(11954, 16),
22156 => conv_std_logic_vector(12040, 16),
22157 => conv_std_logic_vector(12126, 16),
22158 => conv_std_logic_vector(12212, 16),
22159 => conv_std_logic_vector(12298, 16),
22160 => conv_std_logic_vector(12384, 16),
22161 => conv_std_logic_vector(12470, 16),
22162 => conv_std_logic_vector(12556, 16),
22163 => conv_std_logic_vector(12642, 16),
22164 => conv_std_logic_vector(12728, 16),
22165 => conv_std_logic_vector(12814, 16),
22166 => conv_std_logic_vector(12900, 16),
22167 => conv_std_logic_vector(12986, 16),
22168 => conv_std_logic_vector(13072, 16),
22169 => conv_std_logic_vector(13158, 16),
22170 => conv_std_logic_vector(13244, 16),
22171 => conv_std_logic_vector(13330, 16),
22172 => conv_std_logic_vector(13416, 16),
22173 => conv_std_logic_vector(13502, 16),
22174 => conv_std_logic_vector(13588, 16),
22175 => conv_std_logic_vector(13674, 16),
22176 => conv_std_logic_vector(13760, 16),
22177 => conv_std_logic_vector(13846, 16),
22178 => conv_std_logic_vector(13932, 16),
22179 => conv_std_logic_vector(14018, 16),
22180 => conv_std_logic_vector(14104, 16),
22181 => conv_std_logic_vector(14190, 16),
22182 => conv_std_logic_vector(14276, 16),
22183 => conv_std_logic_vector(14362, 16),
22184 => conv_std_logic_vector(14448, 16),
22185 => conv_std_logic_vector(14534, 16),
22186 => conv_std_logic_vector(14620, 16),
22187 => conv_std_logic_vector(14706, 16),
22188 => conv_std_logic_vector(14792, 16),
22189 => conv_std_logic_vector(14878, 16),
22190 => conv_std_logic_vector(14964, 16),
22191 => conv_std_logic_vector(15050, 16),
22192 => conv_std_logic_vector(15136, 16),
22193 => conv_std_logic_vector(15222, 16),
22194 => conv_std_logic_vector(15308, 16),
22195 => conv_std_logic_vector(15394, 16),
22196 => conv_std_logic_vector(15480, 16),
22197 => conv_std_logic_vector(15566, 16),
22198 => conv_std_logic_vector(15652, 16),
22199 => conv_std_logic_vector(15738, 16),
22200 => conv_std_logic_vector(15824, 16),
22201 => conv_std_logic_vector(15910, 16),
22202 => conv_std_logic_vector(15996, 16),
22203 => conv_std_logic_vector(16082, 16),
22204 => conv_std_logic_vector(16168, 16),
22205 => conv_std_logic_vector(16254, 16),
22206 => conv_std_logic_vector(16340, 16),
22207 => conv_std_logic_vector(16426, 16),
22208 => conv_std_logic_vector(16512, 16),
22209 => conv_std_logic_vector(16598, 16),
22210 => conv_std_logic_vector(16684, 16),
22211 => conv_std_logic_vector(16770, 16),
22212 => conv_std_logic_vector(16856, 16),
22213 => conv_std_logic_vector(16942, 16),
22214 => conv_std_logic_vector(17028, 16),
22215 => conv_std_logic_vector(17114, 16),
22216 => conv_std_logic_vector(17200, 16),
22217 => conv_std_logic_vector(17286, 16),
22218 => conv_std_logic_vector(17372, 16),
22219 => conv_std_logic_vector(17458, 16),
22220 => conv_std_logic_vector(17544, 16),
22221 => conv_std_logic_vector(17630, 16),
22222 => conv_std_logic_vector(17716, 16),
22223 => conv_std_logic_vector(17802, 16),
22224 => conv_std_logic_vector(17888, 16),
22225 => conv_std_logic_vector(17974, 16),
22226 => conv_std_logic_vector(18060, 16),
22227 => conv_std_logic_vector(18146, 16),
22228 => conv_std_logic_vector(18232, 16),
22229 => conv_std_logic_vector(18318, 16),
22230 => conv_std_logic_vector(18404, 16),
22231 => conv_std_logic_vector(18490, 16),
22232 => conv_std_logic_vector(18576, 16),
22233 => conv_std_logic_vector(18662, 16),
22234 => conv_std_logic_vector(18748, 16),
22235 => conv_std_logic_vector(18834, 16),
22236 => conv_std_logic_vector(18920, 16),
22237 => conv_std_logic_vector(19006, 16),
22238 => conv_std_logic_vector(19092, 16),
22239 => conv_std_logic_vector(19178, 16),
22240 => conv_std_logic_vector(19264, 16),
22241 => conv_std_logic_vector(19350, 16),
22242 => conv_std_logic_vector(19436, 16),
22243 => conv_std_logic_vector(19522, 16),
22244 => conv_std_logic_vector(19608, 16),
22245 => conv_std_logic_vector(19694, 16),
22246 => conv_std_logic_vector(19780, 16),
22247 => conv_std_logic_vector(19866, 16),
22248 => conv_std_logic_vector(19952, 16),
22249 => conv_std_logic_vector(20038, 16),
22250 => conv_std_logic_vector(20124, 16),
22251 => conv_std_logic_vector(20210, 16),
22252 => conv_std_logic_vector(20296, 16),
22253 => conv_std_logic_vector(20382, 16),
22254 => conv_std_logic_vector(20468, 16),
22255 => conv_std_logic_vector(20554, 16),
22256 => conv_std_logic_vector(20640, 16),
22257 => conv_std_logic_vector(20726, 16),
22258 => conv_std_logic_vector(20812, 16),
22259 => conv_std_logic_vector(20898, 16),
22260 => conv_std_logic_vector(20984, 16),
22261 => conv_std_logic_vector(21070, 16),
22262 => conv_std_logic_vector(21156, 16),
22263 => conv_std_logic_vector(21242, 16),
22264 => conv_std_logic_vector(21328, 16),
22265 => conv_std_logic_vector(21414, 16),
22266 => conv_std_logic_vector(21500, 16),
22267 => conv_std_logic_vector(21586, 16),
22268 => conv_std_logic_vector(21672, 16),
22269 => conv_std_logic_vector(21758, 16),
22270 => conv_std_logic_vector(21844, 16),
22271 => conv_std_logic_vector(21930, 16),
22272 => conv_std_logic_vector(0, 16),
22273 => conv_std_logic_vector(87, 16),
22274 => conv_std_logic_vector(174, 16),
22275 => conv_std_logic_vector(261, 16),
22276 => conv_std_logic_vector(348, 16),
22277 => conv_std_logic_vector(435, 16),
22278 => conv_std_logic_vector(522, 16),
22279 => conv_std_logic_vector(609, 16),
22280 => conv_std_logic_vector(696, 16),
22281 => conv_std_logic_vector(783, 16),
22282 => conv_std_logic_vector(870, 16),
22283 => conv_std_logic_vector(957, 16),
22284 => conv_std_logic_vector(1044, 16),
22285 => conv_std_logic_vector(1131, 16),
22286 => conv_std_logic_vector(1218, 16),
22287 => conv_std_logic_vector(1305, 16),
22288 => conv_std_logic_vector(1392, 16),
22289 => conv_std_logic_vector(1479, 16),
22290 => conv_std_logic_vector(1566, 16),
22291 => conv_std_logic_vector(1653, 16),
22292 => conv_std_logic_vector(1740, 16),
22293 => conv_std_logic_vector(1827, 16),
22294 => conv_std_logic_vector(1914, 16),
22295 => conv_std_logic_vector(2001, 16),
22296 => conv_std_logic_vector(2088, 16),
22297 => conv_std_logic_vector(2175, 16),
22298 => conv_std_logic_vector(2262, 16),
22299 => conv_std_logic_vector(2349, 16),
22300 => conv_std_logic_vector(2436, 16),
22301 => conv_std_logic_vector(2523, 16),
22302 => conv_std_logic_vector(2610, 16),
22303 => conv_std_logic_vector(2697, 16),
22304 => conv_std_logic_vector(2784, 16),
22305 => conv_std_logic_vector(2871, 16),
22306 => conv_std_logic_vector(2958, 16),
22307 => conv_std_logic_vector(3045, 16),
22308 => conv_std_logic_vector(3132, 16),
22309 => conv_std_logic_vector(3219, 16),
22310 => conv_std_logic_vector(3306, 16),
22311 => conv_std_logic_vector(3393, 16),
22312 => conv_std_logic_vector(3480, 16),
22313 => conv_std_logic_vector(3567, 16),
22314 => conv_std_logic_vector(3654, 16),
22315 => conv_std_logic_vector(3741, 16),
22316 => conv_std_logic_vector(3828, 16),
22317 => conv_std_logic_vector(3915, 16),
22318 => conv_std_logic_vector(4002, 16),
22319 => conv_std_logic_vector(4089, 16),
22320 => conv_std_logic_vector(4176, 16),
22321 => conv_std_logic_vector(4263, 16),
22322 => conv_std_logic_vector(4350, 16),
22323 => conv_std_logic_vector(4437, 16),
22324 => conv_std_logic_vector(4524, 16),
22325 => conv_std_logic_vector(4611, 16),
22326 => conv_std_logic_vector(4698, 16),
22327 => conv_std_logic_vector(4785, 16),
22328 => conv_std_logic_vector(4872, 16),
22329 => conv_std_logic_vector(4959, 16),
22330 => conv_std_logic_vector(5046, 16),
22331 => conv_std_logic_vector(5133, 16),
22332 => conv_std_logic_vector(5220, 16),
22333 => conv_std_logic_vector(5307, 16),
22334 => conv_std_logic_vector(5394, 16),
22335 => conv_std_logic_vector(5481, 16),
22336 => conv_std_logic_vector(5568, 16),
22337 => conv_std_logic_vector(5655, 16),
22338 => conv_std_logic_vector(5742, 16),
22339 => conv_std_logic_vector(5829, 16),
22340 => conv_std_logic_vector(5916, 16),
22341 => conv_std_logic_vector(6003, 16),
22342 => conv_std_logic_vector(6090, 16),
22343 => conv_std_logic_vector(6177, 16),
22344 => conv_std_logic_vector(6264, 16),
22345 => conv_std_logic_vector(6351, 16),
22346 => conv_std_logic_vector(6438, 16),
22347 => conv_std_logic_vector(6525, 16),
22348 => conv_std_logic_vector(6612, 16),
22349 => conv_std_logic_vector(6699, 16),
22350 => conv_std_logic_vector(6786, 16),
22351 => conv_std_logic_vector(6873, 16),
22352 => conv_std_logic_vector(6960, 16),
22353 => conv_std_logic_vector(7047, 16),
22354 => conv_std_logic_vector(7134, 16),
22355 => conv_std_logic_vector(7221, 16),
22356 => conv_std_logic_vector(7308, 16),
22357 => conv_std_logic_vector(7395, 16),
22358 => conv_std_logic_vector(7482, 16),
22359 => conv_std_logic_vector(7569, 16),
22360 => conv_std_logic_vector(7656, 16),
22361 => conv_std_logic_vector(7743, 16),
22362 => conv_std_logic_vector(7830, 16),
22363 => conv_std_logic_vector(7917, 16),
22364 => conv_std_logic_vector(8004, 16),
22365 => conv_std_logic_vector(8091, 16),
22366 => conv_std_logic_vector(8178, 16),
22367 => conv_std_logic_vector(8265, 16),
22368 => conv_std_logic_vector(8352, 16),
22369 => conv_std_logic_vector(8439, 16),
22370 => conv_std_logic_vector(8526, 16),
22371 => conv_std_logic_vector(8613, 16),
22372 => conv_std_logic_vector(8700, 16),
22373 => conv_std_logic_vector(8787, 16),
22374 => conv_std_logic_vector(8874, 16),
22375 => conv_std_logic_vector(8961, 16),
22376 => conv_std_logic_vector(9048, 16),
22377 => conv_std_logic_vector(9135, 16),
22378 => conv_std_logic_vector(9222, 16),
22379 => conv_std_logic_vector(9309, 16),
22380 => conv_std_logic_vector(9396, 16),
22381 => conv_std_logic_vector(9483, 16),
22382 => conv_std_logic_vector(9570, 16),
22383 => conv_std_logic_vector(9657, 16),
22384 => conv_std_logic_vector(9744, 16),
22385 => conv_std_logic_vector(9831, 16),
22386 => conv_std_logic_vector(9918, 16),
22387 => conv_std_logic_vector(10005, 16),
22388 => conv_std_logic_vector(10092, 16),
22389 => conv_std_logic_vector(10179, 16),
22390 => conv_std_logic_vector(10266, 16),
22391 => conv_std_logic_vector(10353, 16),
22392 => conv_std_logic_vector(10440, 16),
22393 => conv_std_logic_vector(10527, 16),
22394 => conv_std_logic_vector(10614, 16),
22395 => conv_std_logic_vector(10701, 16),
22396 => conv_std_logic_vector(10788, 16),
22397 => conv_std_logic_vector(10875, 16),
22398 => conv_std_logic_vector(10962, 16),
22399 => conv_std_logic_vector(11049, 16),
22400 => conv_std_logic_vector(11136, 16),
22401 => conv_std_logic_vector(11223, 16),
22402 => conv_std_logic_vector(11310, 16),
22403 => conv_std_logic_vector(11397, 16),
22404 => conv_std_logic_vector(11484, 16),
22405 => conv_std_logic_vector(11571, 16),
22406 => conv_std_logic_vector(11658, 16),
22407 => conv_std_logic_vector(11745, 16),
22408 => conv_std_logic_vector(11832, 16),
22409 => conv_std_logic_vector(11919, 16),
22410 => conv_std_logic_vector(12006, 16),
22411 => conv_std_logic_vector(12093, 16),
22412 => conv_std_logic_vector(12180, 16),
22413 => conv_std_logic_vector(12267, 16),
22414 => conv_std_logic_vector(12354, 16),
22415 => conv_std_logic_vector(12441, 16),
22416 => conv_std_logic_vector(12528, 16),
22417 => conv_std_logic_vector(12615, 16),
22418 => conv_std_logic_vector(12702, 16),
22419 => conv_std_logic_vector(12789, 16),
22420 => conv_std_logic_vector(12876, 16),
22421 => conv_std_logic_vector(12963, 16),
22422 => conv_std_logic_vector(13050, 16),
22423 => conv_std_logic_vector(13137, 16),
22424 => conv_std_logic_vector(13224, 16),
22425 => conv_std_logic_vector(13311, 16),
22426 => conv_std_logic_vector(13398, 16),
22427 => conv_std_logic_vector(13485, 16),
22428 => conv_std_logic_vector(13572, 16),
22429 => conv_std_logic_vector(13659, 16),
22430 => conv_std_logic_vector(13746, 16),
22431 => conv_std_logic_vector(13833, 16),
22432 => conv_std_logic_vector(13920, 16),
22433 => conv_std_logic_vector(14007, 16),
22434 => conv_std_logic_vector(14094, 16),
22435 => conv_std_logic_vector(14181, 16),
22436 => conv_std_logic_vector(14268, 16),
22437 => conv_std_logic_vector(14355, 16),
22438 => conv_std_logic_vector(14442, 16),
22439 => conv_std_logic_vector(14529, 16),
22440 => conv_std_logic_vector(14616, 16),
22441 => conv_std_logic_vector(14703, 16),
22442 => conv_std_logic_vector(14790, 16),
22443 => conv_std_logic_vector(14877, 16),
22444 => conv_std_logic_vector(14964, 16),
22445 => conv_std_logic_vector(15051, 16),
22446 => conv_std_logic_vector(15138, 16),
22447 => conv_std_logic_vector(15225, 16),
22448 => conv_std_logic_vector(15312, 16),
22449 => conv_std_logic_vector(15399, 16),
22450 => conv_std_logic_vector(15486, 16),
22451 => conv_std_logic_vector(15573, 16),
22452 => conv_std_logic_vector(15660, 16),
22453 => conv_std_logic_vector(15747, 16),
22454 => conv_std_logic_vector(15834, 16),
22455 => conv_std_logic_vector(15921, 16),
22456 => conv_std_logic_vector(16008, 16),
22457 => conv_std_logic_vector(16095, 16),
22458 => conv_std_logic_vector(16182, 16),
22459 => conv_std_logic_vector(16269, 16),
22460 => conv_std_logic_vector(16356, 16),
22461 => conv_std_logic_vector(16443, 16),
22462 => conv_std_logic_vector(16530, 16),
22463 => conv_std_logic_vector(16617, 16),
22464 => conv_std_logic_vector(16704, 16),
22465 => conv_std_logic_vector(16791, 16),
22466 => conv_std_logic_vector(16878, 16),
22467 => conv_std_logic_vector(16965, 16),
22468 => conv_std_logic_vector(17052, 16),
22469 => conv_std_logic_vector(17139, 16),
22470 => conv_std_logic_vector(17226, 16),
22471 => conv_std_logic_vector(17313, 16),
22472 => conv_std_logic_vector(17400, 16),
22473 => conv_std_logic_vector(17487, 16),
22474 => conv_std_logic_vector(17574, 16),
22475 => conv_std_logic_vector(17661, 16),
22476 => conv_std_logic_vector(17748, 16),
22477 => conv_std_logic_vector(17835, 16),
22478 => conv_std_logic_vector(17922, 16),
22479 => conv_std_logic_vector(18009, 16),
22480 => conv_std_logic_vector(18096, 16),
22481 => conv_std_logic_vector(18183, 16),
22482 => conv_std_logic_vector(18270, 16),
22483 => conv_std_logic_vector(18357, 16),
22484 => conv_std_logic_vector(18444, 16),
22485 => conv_std_logic_vector(18531, 16),
22486 => conv_std_logic_vector(18618, 16),
22487 => conv_std_logic_vector(18705, 16),
22488 => conv_std_logic_vector(18792, 16),
22489 => conv_std_logic_vector(18879, 16),
22490 => conv_std_logic_vector(18966, 16),
22491 => conv_std_logic_vector(19053, 16),
22492 => conv_std_logic_vector(19140, 16),
22493 => conv_std_logic_vector(19227, 16),
22494 => conv_std_logic_vector(19314, 16),
22495 => conv_std_logic_vector(19401, 16),
22496 => conv_std_logic_vector(19488, 16),
22497 => conv_std_logic_vector(19575, 16),
22498 => conv_std_logic_vector(19662, 16),
22499 => conv_std_logic_vector(19749, 16),
22500 => conv_std_logic_vector(19836, 16),
22501 => conv_std_logic_vector(19923, 16),
22502 => conv_std_logic_vector(20010, 16),
22503 => conv_std_logic_vector(20097, 16),
22504 => conv_std_logic_vector(20184, 16),
22505 => conv_std_logic_vector(20271, 16),
22506 => conv_std_logic_vector(20358, 16),
22507 => conv_std_logic_vector(20445, 16),
22508 => conv_std_logic_vector(20532, 16),
22509 => conv_std_logic_vector(20619, 16),
22510 => conv_std_logic_vector(20706, 16),
22511 => conv_std_logic_vector(20793, 16),
22512 => conv_std_logic_vector(20880, 16),
22513 => conv_std_logic_vector(20967, 16),
22514 => conv_std_logic_vector(21054, 16),
22515 => conv_std_logic_vector(21141, 16),
22516 => conv_std_logic_vector(21228, 16),
22517 => conv_std_logic_vector(21315, 16),
22518 => conv_std_logic_vector(21402, 16),
22519 => conv_std_logic_vector(21489, 16),
22520 => conv_std_logic_vector(21576, 16),
22521 => conv_std_logic_vector(21663, 16),
22522 => conv_std_logic_vector(21750, 16),
22523 => conv_std_logic_vector(21837, 16),
22524 => conv_std_logic_vector(21924, 16),
22525 => conv_std_logic_vector(22011, 16),
22526 => conv_std_logic_vector(22098, 16),
22527 => conv_std_logic_vector(22185, 16),
22528 => conv_std_logic_vector(0, 16),
22529 => conv_std_logic_vector(88, 16),
22530 => conv_std_logic_vector(176, 16),
22531 => conv_std_logic_vector(264, 16),
22532 => conv_std_logic_vector(352, 16),
22533 => conv_std_logic_vector(440, 16),
22534 => conv_std_logic_vector(528, 16),
22535 => conv_std_logic_vector(616, 16),
22536 => conv_std_logic_vector(704, 16),
22537 => conv_std_logic_vector(792, 16),
22538 => conv_std_logic_vector(880, 16),
22539 => conv_std_logic_vector(968, 16),
22540 => conv_std_logic_vector(1056, 16),
22541 => conv_std_logic_vector(1144, 16),
22542 => conv_std_logic_vector(1232, 16),
22543 => conv_std_logic_vector(1320, 16),
22544 => conv_std_logic_vector(1408, 16),
22545 => conv_std_logic_vector(1496, 16),
22546 => conv_std_logic_vector(1584, 16),
22547 => conv_std_logic_vector(1672, 16),
22548 => conv_std_logic_vector(1760, 16),
22549 => conv_std_logic_vector(1848, 16),
22550 => conv_std_logic_vector(1936, 16),
22551 => conv_std_logic_vector(2024, 16),
22552 => conv_std_logic_vector(2112, 16),
22553 => conv_std_logic_vector(2200, 16),
22554 => conv_std_logic_vector(2288, 16),
22555 => conv_std_logic_vector(2376, 16),
22556 => conv_std_logic_vector(2464, 16),
22557 => conv_std_logic_vector(2552, 16),
22558 => conv_std_logic_vector(2640, 16),
22559 => conv_std_logic_vector(2728, 16),
22560 => conv_std_logic_vector(2816, 16),
22561 => conv_std_logic_vector(2904, 16),
22562 => conv_std_logic_vector(2992, 16),
22563 => conv_std_logic_vector(3080, 16),
22564 => conv_std_logic_vector(3168, 16),
22565 => conv_std_logic_vector(3256, 16),
22566 => conv_std_logic_vector(3344, 16),
22567 => conv_std_logic_vector(3432, 16),
22568 => conv_std_logic_vector(3520, 16),
22569 => conv_std_logic_vector(3608, 16),
22570 => conv_std_logic_vector(3696, 16),
22571 => conv_std_logic_vector(3784, 16),
22572 => conv_std_logic_vector(3872, 16),
22573 => conv_std_logic_vector(3960, 16),
22574 => conv_std_logic_vector(4048, 16),
22575 => conv_std_logic_vector(4136, 16),
22576 => conv_std_logic_vector(4224, 16),
22577 => conv_std_logic_vector(4312, 16),
22578 => conv_std_logic_vector(4400, 16),
22579 => conv_std_logic_vector(4488, 16),
22580 => conv_std_logic_vector(4576, 16),
22581 => conv_std_logic_vector(4664, 16),
22582 => conv_std_logic_vector(4752, 16),
22583 => conv_std_logic_vector(4840, 16),
22584 => conv_std_logic_vector(4928, 16),
22585 => conv_std_logic_vector(5016, 16),
22586 => conv_std_logic_vector(5104, 16),
22587 => conv_std_logic_vector(5192, 16),
22588 => conv_std_logic_vector(5280, 16),
22589 => conv_std_logic_vector(5368, 16),
22590 => conv_std_logic_vector(5456, 16),
22591 => conv_std_logic_vector(5544, 16),
22592 => conv_std_logic_vector(5632, 16),
22593 => conv_std_logic_vector(5720, 16),
22594 => conv_std_logic_vector(5808, 16),
22595 => conv_std_logic_vector(5896, 16),
22596 => conv_std_logic_vector(5984, 16),
22597 => conv_std_logic_vector(6072, 16),
22598 => conv_std_logic_vector(6160, 16),
22599 => conv_std_logic_vector(6248, 16),
22600 => conv_std_logic_vector(6336, 16),
22601 => conv_std_logic_vector(6424, 16),
22602 => conv_std_logic_vector(6512, 16),
22603 => conv_std_logic_vector(6600, 16),
22604 => conv_std_logic_vector(6688, 16),
22605 => conv_std_logic_vector(6776, 16),
22606 => conv_std_logic_vector(6864, 16),
22607 => conv_std_logic_vector(6952, 16),
22608 => conv_std_logic_vector(7040, 16),
22609 => conv_std_logic_vector(7128, 16),
22610 => conv_std_logic_vector(7216, 16),
22611 => conv_std_logic_vector(7304, 16),
22612 => conv_std_logic_vector(7392, 16),
22613 => conv_std_logic_vector(7480, 16),
22614 => conv_std_logic_vector(7568, 16),
22615 => conv_std_logic_vector(7656, 16),
22616 => conv_std_logic_vector(7744, 16),
22617 => conv_std_logic_vector(7832, 16),
22618 => conv_std_logic_vector(7920, 16),
22619 => conv_std_logic_vector(8008, 16),
22620 => conv_std_logic_vector(8096, 16),
22621 => conv_std_logic_vector(8184, 16),
22622 => conv_std_logic_vector(8272, 16),
22623 => conv_std_logic_vector(8360, 16),
22624 => conv_std_logic_vector(8448, 16),
22625 => conv_std_logic_vector(8536, 16),
22626 => conv_std_logic_vector(8624, 16),
22627 => conv_std_logic_vector(8712, 16),
22628 => conv_std_logic_vector(8800, 16),
22629 => conv_std_logic_vector(8888, 16),
22630 => conv_std_logic_vector(8976, 16),
22631 => conv_std_logic_vector(9064, 16),
22632 => conv_std_logic_vector(9152, 16),
22633 => conv_std_logic_vector(9240, 16),
22634 => conv_std_logic_vector(9328, 16),
22635 => conv_std_logic_vector(9416, 16),
22636 => conv_std_logic_vector(9504, 16),
22637 => conv_std_logic_vector(9592, 16),
22638 => conv_std_logic_vector(9680, 16),
22639 => conv_std_logic_vector(9768, 16),
22640 => conv_std_logic_vector(9856, 16),
22641 => conv_std_logic_vector(9944, 16),
22642 => conv_std_logic_vector(10032, 16),
22643 => conv_std_logic_vector(10120, 16),
22644 => conv_std_logic_vector(10208, 16),
22645 => conv_std_logic_vector(10296, 16),
22646 => conv_std_logic_vector(10384, 16),
22647 => conv_std_logic_vector(10472, 16),
22648 => conv_std_logic_vector(10560, 16),
22649 => conv_std_logic_vector(10648, 16),
22650 => conv_std_logic_vector(10736, 16),
22651 => conv_std_logic_vector(10824, 16),
22652 => conv_std_logic_vector(10912, 16),
22653 => conv_std_logic_vector(11000, 16),
22654 => conv_std_logic_vector(11088, 16),
22655 => conv_std_logic_vector(11176, 16),
22656 => conv_std_logic_vector(11264, 16),
22657 => conv_std_logic_vector(11352, 16),
22658 => conv_std_logic_vector(11440, 16),
22659 => conv_std_logic_vector(11528, 16),
22660 => conv_std_logic_vector(11616, 16),
22661 => conv_std_logic_vector(11704, 16),
22662 => conv_std_logic_vector(11792, 16),
22663 => conv_std_logic_vector(11880, 16),
22664 => conv_std_logic_vector(11968, 16),
22665 => conv_std_logic_vector(12056, 16),
22666 => conv_std_logic_vector(12144, 16),
22667 => conv_std_logic_vector(12232, 16),
22668 => conv_std_logic_vector(12320, 16),
22669 => conv_std_logic_vector(12408, 16),
22670 => conv_std_logic_vector(12496, 16),
22671 => conv_std_logic_vector(12584, 16),
22672 => conv_std_logic_vector(12672, 16),
22673 => conv_std_logic_vector(12760, 16),
22674 => conv_std_logic_vector(12848, 16),
22675 => conv_std_logic_vector(12936, 16),
22676 => conv_std_logic_vector(13024, 16),
22677 => conv_std_logic_vector(13112, 16),
22678 => conv_std_logic_vector(13200, 16),
22679 => conv_std_logic_vector(13288, 16),
22680 => conv_std_logic_vector(13376, 16),
22681 => conv_std_logic_vector(13464, 16),
22682 => conv_std_logic_vector(13552, 16),
22683 => conv_std_logic_vector(13640, 16),
22684 => conv_std_logic_vector(13728, 16),
22685 => conv_std_logic_vector(13816, 16),
22686 => conv_std_logic_vector(13904, 16),
22687 => conv_std_logic_vector(13992, 16),
22688 => conv_std_logic_vector(14080, 16),
22689 => conv_std_logic_vector(14168, 16),
22690 => conv_std_logic_vector(14256, 16),
22691 => conv_std_logic_vector(14344, 16),
22692 => conv_std_logic_vector(14432, 16),
22693 => conv_std_logic_vector(14520, 16),
22694 => conv_std_logic_vector(14608, 16),
22695 => conv_std_logic_vector(14696, 16),
22696 => conv_std_logic_vector(14784, 16),
22697 => conv_std_logic_vector(14872, 16),
22698 => conv_std_logic_vector(14960, 16),
22699 => conv_std_logic_vector(15048, 16),
22700 => conv_std_logic_vector(15136, 16),
22701 => conv_std_logic_vector(15224, 16),
22702 => conv_std_logic_vector(15312, 16),
22703 => conv_std_logic_vector(15400, 16),
22704 => conv_std_logic_vector(15488, 16),
22705 => conv_std_logic_vector(15576, 16),
22706 => conv_std_logic_vector(15664, 16),
22707 => conv_std_logic_vector(15752, 16),
22708 => conv_std_logic_vector(15840, 16),
22709 => conv_std_logic_vector(15928, 16),
22710 => conv_std_logic_vector(16016, 16),
22711 => conv_std_logic_vector(16104, 16),
22712 => conv_std_logic_vector(16192, 16),
22713 => conv_std_logic_vector(16280, 16),
22714 => conv_std_logic_vector(16368, 16),
22715 => conv_std_logic_vector(16456, 16),
22716 => conv_std_logic_vector(16544, 16),
22717 => conv_std_logic_vector(16632, 16),
22718 => conv_std_logic_vector(16720, 16),
22719 => conv_std_logic_vector(16808, 16),
22720 => conv_std_logic_vector(16896, 16),
22721 => conv_std_logic_vector(16984, 16),
22722 => conv_std_logic_vector(17072, 16),
22723 => conv_std_logic_vector(17160, 16),
22724 => conv_std_logic_vector(17248, 16),
22725 => conv_std_logic_vector(17336, 16),
22726 => conv_std_logic_vector(17424, 16),
22727 => conv_std_logic_vector(17512, 16),
22728 => conv_std_logic_vector(17600, 16),
22729 => conv_std_logic_vector(17688, 16),
22730 => conv_std_logic_vector(17776, 16),
22731 => conv_std_logic_vector(17864, 16),
22732 => conv_std_logic_vector(17952, 16),
22733 => conv_std_logic_vector(18040, 16),
22734 => conv_std_logic_vector(18128, 16),
22735 => conv_std_logic_vector(18216, 16),
22736 => conv_std_logic_vector(18304, 16),
22737 => conv_std_logic_vector(18392, 16),
22738 => conv_std_logic_vector(18480, 16),
22739 => conv_std_logic_vector(18568, 16),
22740 => conv_std_logic_vector(18656, 16),
22741 => conv_std_logic_vector(18744, 16),
22742 => conv_std_logic_vector(18832, 16),
22743 => conv_std_logic_vector(18920, 16),
22744 => conv_std_logic_vector(19008, 16),
22745 => conv_std_logic_vector(19096, 16),
22746 => conv_std_logic_vector(19184, 16),
22747 => conv_std_logic_vector(19272, 16),
22748 => conv_std_logic_vector(19360, 16),
22749 => conv_std_logic_vector(19448, 16),
22750 => conv_std_logic_vector(19536, 16),
22751 => conv_std_logic_vector(19624, 16),
22752 => conv_std_logic_vector(19712, 16),
22753 => conv_std_logic_vector(19800, 16),
22754 => conv_std_logic_vector(19888, 16),
22755 => conv_std_logic_vector(19976, 16),
22756 => conv_std_logic_vector(20064, 16),
22757 => conv_std_logic_vector(20152, 16),
22758 => conv_std_logic_vector(20240, 16),
22759 => conv_std_logic_vector(20328, 16),
22760 => conv_std_logic_vector(20416, 16),
22761 => conv_std_logic_vector(20504, 16),
22762 => conv_std_logic_vector(20592, 16),
22763 => conv_std_logic_vector(20680, 16),
22764 => conv_std_logic_vector(20768, 16),
22765 => conv_std_logic_vector(20856, 16),
22766 => conv_std_logic_vector(20944, 16),
22767 => conv_std_logic_vector(21032, 16),
22768 => conv_std_logic_vector(21120, 16),
22769 => conv_std_logic_vector(21208, 16),
22770 => conv_std_logic_vector(21296, 16),
22771 => conv_std_logic_vector(21384, 16),
22772 => conv_std_logic_vector(21472, 16),
22773 => conv_std_logic_vector(21560, 16),
22774 => conv_std_logic_vector(21648, 16),
22775 => conv_std_logic_vector(21736, 16),
22776 => conv_std_logic_vector(21824, 16),
22777 => conv_std_logic_vector(21912, 16),
22778 => conv_std_logic_vector(22000, 16),
22779 => conv_std_logic_vector(22088, 16),
22780 => conv_std_logic_vector(22176, 16),
22781 => conv_std_logic_vector(22264, 16),
22782 => conv_std_logic_vector(22352, 16),
22783 => conv_std_logic_vector(22440, 16),
22784 => conv_std_logic_vector(0, 16),
22785 => conv_std_logic_vector(89, 16),
22786 => conv_std_logic_vector(178, 16),
22787 => conv_std_logic_vector(267, 16),
22788 => conv_std_logic_vector(356, 16),
22789 => conv_std_logic_vector(445, 16),
22790 => conv_std_logic_vector(534, 16),
22791 => conv_std_logic_vector(623, 16),
22792 => conv_std_logic_vector(712, 16),
22793 => conv_std_logic_vector(801, 16),
22794 => conv_std_logic_vector(890, 16),
22795 => conv_std_logic_vector(979, 16),
22796 => conv_std_logic_vector(1068, 16),
22797 => conv_std_logic_vector(1157, 16),
22798 => conv_std_logic_vector(1246, 16),
22799 => conv_std_logic_vector(1335, 16),
22800 => conv_std_logic_vector(1424, 16),
22801 => conv_std_logic_vector(1513, 16),
22802 => conv_std_logic_vector(1602, 16),
22803 => conv_std_logic_vector(1691, 16),
22804 => conv_std_logic_vector(1780, 16),
22805 => conv_std_logic_vector(1869, 16),
22806 => conv_std_logic_vector(1958, 16),
22807 => conv_std_logic_vector(2047, 16),
22808 => conv_std_logic_vector(2136, 16),
22809 => conv_std_logic_vector(2225, 16),
22810 => conv_std_logic_vector(2314, 16),
22811 => conv_std_logic_vector(2403, 16),
22812 => conv_std_logic_vector(2492, 16),
22813 => conv_std_logic_vector(2581, 16),
22814 => conv_std_logic_vector(2670, 16),
22815 => conv_std_logic_vector(2759, 16),
22816 => conv_std_logic_vector(2848, 16),
22817 => conv_std_logic_vector(2937, 16),
22818 => conv_std_logic_vector(3026, 16),
22819 => conv_std_logic_vector(3115, 16),
22820 => conv_std_logic_vector(3204, 16),
22821 => conv_std_logic_vector(3293, 16),
22822 => conv_std_logic_vector(3382, 16),
22823 => conv_std_logic_vector(3471, 16),
22824 => conv_std_logic_vector(3560, 16),
22825 => conv_std_logic_vector(3649, 16),
22826 => conv_std_logic_vector(3738, 16),
22827 => conv_std_logic_vector(3827, 16),
22828 => conv_std_logic_vector(3916, 16),
22829 => conv_std_logic_vector(4005, 16),
22830 => conv_std_logic_vector(4094, 16),
22831 => conv_std_logic_vector(4183, 16),
22832 => conv_std_logic_vector(4272, 16),
22833 => conv_std_logic_vector(4361, 16),
22834 => conv_std_logic_vector(4450, 16),
22835 => conv_std_logic_vector(4539, 16),
22836 => conv_std_logic_vector(4628, 16),
22837 => conv_std_logic_vector(4717, 16),
22838 => conv_std_logic_vector(4806, 16),
22839 => conv_std_logic_vector(4895, 16),
22840 => conv_std_logic_vector(4984, 16),
22841 => conv_std_logic_vector(5073, 16),
22842 => conv_std_logic_vector(5162, 16),
22843 => conv_std_logic_vector(5251, 16),
22844 => conv_std_logic_vector(5340, 16),
22845 => conv_std_logic_vector(5429, 16),
22846 => conv_std_logic_vector(5518, 16),
22847 => conv_std_logic_vector(5607, 16),
22848 => conv_std_logic_vector(5696, 16),
22849 => conv_std_logic_vector(5785, 16),
22850 => conv_std_logic_vector(5874, 16),
22851 => conv_std_logic_vector(5963, 16),
22852 => conv_std_logic_vector(6052, 16),
22853 => conv_std_logic_vector(6141, 16),
22854 => conv_std_logic_vector(6230, 16),
22855 => conv_std_logic_vector(6319, 16),
22856 => conv_std_logic_vector(6408, 16),
22857 => conv_std_logic_vector(6497, 16),
22858 => conv_std_logic_vector(6586, 16),
22859 => conv_std_logic_vector(6675, 16),
22860 => conv_std_logic_vector(6764, 16),
22861 => conv_std_logic_vector(6853, 16),
22862 => conv_std_logic_vector(6942, 16),
22863 => conv_std_logic_vector(7031, 16),
22864 => conv_std_logic_vector(7120, 16),
22865 => conv_std_logic_vector(7209, 16),
22866 => conv_std_logic_vector(7298, 16),
22867 => conv_std_logic_vector(7387, 16),
22868 => conv_std_logic_vector(7476, 16),
22869 => conv_std_logic_vector(7565, 16),
22870 => conv_std_logic_vector(7654, 16),
22871 => conv_std_logic_vector(7743, 16),
22872 => conv_std_logic_vector(7832, 16),
22873 => conv_std_logic_vector(7921, 16),
22874 => conv_std_logic_vector(8010, 16),
22875 => conv_std_logic_vector(8099, 16),
22876 => conv_std_logic_vector(8188, 16),
22877 => conv_std_logic_vector(8277, 16),
22878 => conv_std_logic_vector(8366, 16),
22879 => conv_std_logic_vector(8455, 16),
22880 => conv_std_logic_vector(8544, 16),
22881 => conv_std_logic_vector(8633, 16),
22882 => conv_std_logic_vector(8722, 16),
22883 => conv_std_logic_vector(8811, 16),
22884 => conv_std_logic_vector(8900, 16),
22885 => conv_std_logic_vector(8989, 16),
22886 => conv_std_logic_vector(9078, 16),
22887 => conv_std_logic_vector(9167, 16),
22888 => conv_std_logic_vector(9256, 16),
22889 => conv_std_logic_vector(9345, 16),
22890 => conv_std_logic_vector(9434, 16),
22891 => conv_std_logic_vector(9523, 16),
22892 => conv_std_logic_vector(9612, 16),
22893 => conv_std_logic_vector(9701, 16),
22894 => conv_std_logic_vector(9790, 16),
22895 => conv_std_logic_vector(9879, 16),
22896 => conv_std_logic_vector(9968, 16),
22897 => conv_std_logic_vector(10057, 16),
22898 => conv_std_logic_vector(10146, 16),
22899 => conv_std_logic_vector(10235, 16),
22900 => conv_std_logic_vector(10324, 16),
22901 => conv_std_logic_vector(10413, 16),
22902 => conv_std_logic_vector(10502, 16),
22903 => conv_std_logic_vector(10591, 16),
22904 => conv_std_logic_vector(10680, 16),
22905 => conv_std_logic_vector(10769, 16),
22906 => conv_std_logic_vector(10858, 16),
22907 => conv_std_logic_vector(10947, 16),
22908 => conv_std_logic_vector(11036, 16),
22909 => conv_std_logic_vector(11125, 16),
22910 => conv_std_logic_vector(11214, 16),
22911 => conv_std_logic_vector(11303, 16),
22912 => conv_std_logic_vector(11392, 16),
22913 => conv_std_logic_vector(11481, 16),
22914 => conv_std_logic_vector(11570, 16),
22915 => conv_std_logic_vector(11659, 16),
22916 => conv_std_logic_vector(11748, 16),
22917 => conv_std_logic_vector(11837, 16),
22918 => conv_std_logic_vector(11926, 16),
22919 => conv_std_logic_vector(12015, 16),
22920 => conv_std_logic_vector(12104, 16),
22921 => conv_std_logic_vector(12193, 16),
22922 => conv_std_logic_vector(12282, 16),
22923 => conv_std_logic_vector(12371, 16),
22924 => conv_std_logic_vector(12460, 16),
22925 => conv_std_logic_vector(12549, 16),
22926 => conv_std_logic_vector(12638, 16),
22927 => conv_std_logic_vector(12727, 16),
22928 => conv_std_logic_vector(12816, 16),
22929 => conv_std_logic_vector(12905, 16),
22930 => conv_std_logic_vector(12994, 16),
22931 => conv_std_logic_vector(13083, 16),
22932 => conv_std_logic_vector(13172, 16),
22933 => conv_std_logic_vector(13261, 16),
22934 => conv_std_logic_vector(13350, 16),
22935 => conv_std_logic_vector(13439, 16),
22936 => conv_std_logic_vector(13528, 16),
22937 => conv_std_logic_vector(13617, 16),
22938 => conv_std_logic_vector(13706, 16),
22939 => conv_std_logic_vector(13795, 16),
22940 => conv_std_logic_vector(13884, 16),
22941 => conv_std_logic_vector(13973, 16),
22942 => conv_std_logic_vector(14062, 16),
22943 => conv_std_logic_vector(14151, 16),
22944 => conv_std_logic_vector(14240, 16),
22945 => conv_std_logic_vector(14329, 16),
22946 => conv_std_logic_vector(14418, 16),
22947 => conv_std_logic_vector(14507, 16),
22948 => conv_std_logic_vector(14596, 16),
22949 => conv_std_logic_vector(14685, 16),
22950 => conv_std_logic_vector(14774, 16),
22951 => conv_std_logic_vector(14863, 16),
22952 => conv_std_logic_vector(14952, 16),
22953 => conv_std_logic_vector(15041, 16),
22954 => conv_std_logic_vector(15130, 16),
22955 => conv_std_logic_vector(15219, 16),
22956 => conv_std_logic_vector(15308, 16),
22957 => conv_std_logic_vector(15397, 16),
22958 => conv_std_logic_vector(15486, 16),
22959 => conv_std_logic_vector(15575, 16),
22960 => conv_std_logic_vector(15664, 16),
22961 => conv_std_logic_vector(15753, 16),
22962 => conv_std_logic_vector(15842, 16),
22963 => conv_std_logic_vector(15931, 16),
22964 => conv_std_logic_vector(16020, 16),
22965 => conv_std_logic_vector(16109, 16),
22966 => conv_std_logic_vector(16198, 16),
22967 => conv_std_logic_vector(16287, 16),
22968 => conv_std_logic_vector(16376, 16),
22969 => conv_std_logic_vector(16465, 16),
22970 => conv_std_logic_vector(16554, 16),
22971 => conv_std_logic_vector(16643, 16),
22972 => conv_std_logic_vector(16732, 16),
22973 => conv_std_logic_vector(16821, 16),
22974 => conv_std_logic_vector(16910, 16),
22975 => conv_std_logic_vector(16999, 16),
22976 => conv_std_logic_vector(17088, 16),
22977 => conv_std_logic_vector(17177, 16),
22978 => conv_std_logic_vector(17266, 16),
22979 => conv_std_logic_vector(17355, 16),
22980 => conv_std_logic_vector(17444, 16),
22981 => conv_std_logic_vector(17533, 16),
22982 => conv_std_logic_vector(17622, 16),
22983 => conv_std_logic_vector(17711, 16),
22984 => conv_std_logic_vector(17800, 16),
22985 => conv_std_logic_vector(17889, 16),
22986 => conv_std_logic_vector(17978, 16),
22987 => conv_std_logic_vector(18067, 16),
22988 => conv_std_logic_vector(18156, 16),
22989 => conv_std_logic_vector(18245, 16),
22990 => conv_std_logic_vector(18334, 16),
22991 => conv_std_logic_vector(18423, 16),
22992 => conv_std_logic_vector(18512, 16),
22993 => conv_std_logic_vector(18601, 16),
22994 => conv_std_logic_vector(18690, 16),
22995 => conv_std_logic_vector(18779, 16),
22996 => conv_std_logic_vector(18868, 16),
22997 => conv_std_logic_vector(18957, 16),
22998 => conv_std_logic_vector(19046, 16),
22999 => conv_std_logic_vector(19135, 16),
23000 => conv_std_logic_vector(19224, 16),
23001 => conv_std_logic_vector(19313, 16),
23002 => conv_std_logic_vector(19402, 16),
23003 => conv_std_logic_vector(19491, 16),
23004 => conv_std_logic_vector(19580, 16),
23005 => conv_std_logic_vector(19669, 16),
23006 => conv_std_logic_vector(19758, 16),
23007 => conv_std_logic_vector(19847, 16),
23008 => conv_std_logic_vector(19936, 16),
23009 => conv_std_logic_vector(20025, 16),
23010 => conv_std_logic_vector(20114, 16),
23011 => conv_std_logic_vector(20203, 16),
23012 => conv_std_logic_vector(20292, 16),
23013 => conv_std_logic_vector(20381, 16),
23014 => conv_std_logic_vector(20470, 16),
23015 => conv_std_logic_vector(20559, 16),
23016 => conv_std_logic_vector(20648, 16),
23017 => conv_std_logic_vector(20737, 16),
23018 => conv_std_logic_vector(20826, 16),
23019 => conv_std_logic_vector(20915, 16),
23020 => conv_std_logic_vector(21004, 16),
23021 => conv_std_logic_vector(21093, 16),
23022 => conv_std_logic_vector(21182, 16),
23023 => conv_std_logic_vector(21271, 16),
23024 => conv_std_logic_vector(21360, 16),
23025 => conv_std_logic_vector(21449, 16),
23026 => conv_std_logic_vector(21538, 16),
23027 => conv_std_logic_vector(21627, 16),
23028 => conv_std_logic_vector(21716, 16),
23029 => conv_std_logic_vector(21805, 16),
23030 => conv_std_logic_vector(21894, 16),
23031 => conv_std_logic_vector(21983, 16),
23032 => conv_std_logic_vector(22072, 16),
23033 => conv_std_logic_vector(22161, 16),
23034 => conv_std_logic_vector(22250, 16),
23035 => conv_std_logic_vector(22339, 16),
23036 => conv_std_logic_vector(22428, 16),
23037 => conv_std_logic_vector(22517, 16),
23038 => conv_std_logic_vector(22606, 16),
23039 => conv_std_logic_vector(22695, 16),
23040 => conv_std_logic_vector(0, 16),
23041 => conv_std_logic_vector(90, 16),
23042 => conv_std_logic_vector(180, 16),
23043 => conv_std_logic_vector(270, 16),
23044 => conv_std_logic_vector(360, 16),
23045 => conv_std_logic_vector(450, 16),
23046 => conv_std_logic_vector(540, 16),
23047 => conv_std_logic_vector(630, 16),
23048 => conv_std_logic_vector(720, 16),
23049 => conv_std_logic_vector(810, 16),
23050 => conv_std_logic_vector(900, 16),
23051 => conv_std_logic_vector(990, 16),
23052 => conv_std_logic_vector(1080, 16),
23053 => conv_std_logic_vector(1170, 16),
23054 => conv_std_logic_vector(1260, 16),
23055 => conv_std_logic_vector(1350, 16),
23056 => conv_std_logic_vector(1440, 16),
23057 => conv_std_logic_vector(1530, 16),
23058 => conv_std_logic_vector(1620, 16),
23059 => conv_std_logic_vector(1710, 16),
23060 => conv_std_logic_vector(1800, 16),
23061 => conv_std_logic_vector(1890, 16),
23062 => conv_std_logic_vector(1980, 16),
23063 => conv_std_logic_vector(2070, 16),
23064 => conv_std_logic_vector(2160, 16),
23065 => conv_std_logic_vector(2250, 16),
23066 => conv_std_logic_vector(2340, 16),
23067 => conv_std_logic_vector(2430, 16),
23068 => conv_std_logic_vector(2520, 16),
23069 => conv_std_logic_vector(2610, 16),
23070 => conv_std_logic_vector(2700, 16),
23071 => conv_std_logic_vector(2790, 16),
23072 => conv_std_logic_vector(2880, 16),
23073 => conv_std_logic_vector(2970, 16),
23074 => conv_std_logic_vector(3060, 16),
23075 => conv_std_logic_vector(3150, 16),
23076 => conv_std_logic_vector(3240, 16),
23077 => conv_std_logic_vector(3330, 16),
23078 => conv_std_logic_vector(3420, 16),
23079 => conv_std_logic_vector(3510, 16),
23080 => conv_std_logic_vector(3600, 16),
23081 => conv_std_logic_vector(3690, 16),
23082 => conv_std_logic_vector(3780, 16),
23083 => conv_std_logic_vector(3870, 16),
23084 => conv_std_logic_vector(3960, 16),
23085 => conv_std_logic_vector(4050, 16),
23086 => conv_std_logic_vector(4140, 16),
23087 => conv_std_logic_vector(4230, 16),
23088 => conv_std_logic_vector(4320, 16),
23089 => conv_std_logic_vector(4410, 16),
23090 => conv_std_logic_vector(4500, 16),
23091 => conv_std_logic_vector(4590, 16),
23092 => conv_std_logic_vector(4680, 16),
23093 => conv_std_logic_vector(4770, 16),
23094 => conv_std_logic_vector(4860, 16),
23095 => conv_std_logic_vector(4950, 16),
23096 => conv_std_logic_vector(5040, 16),
23097 => conv_std_logic_vector(5130, 16),
23098 => conv_std_logic_vector(5220, 16),
23099 => conv_std_logic_vector(5310, 16),
23100 => conv_std_logic_vector(5400, 16),
23101 => conv_std_logic_vector(5490, 16),
23102 => conv_std_logic_vector(5580, 16),
23103 => conv_std_logic_vector(5670, 16),
23104 => conv_std_logic_vector(5760, 16),
23105 => conv_std_logic_vector(5850, 16),
23106 => conv_std_logic_vector(5940, 16),
23107 => conv_std_logic_vector(6030, 16),
23108 => conv_std_logic_vector(6120, 16),
23109 => conv_std_logic_vector(6210, 16),
23110 => conv_std_logic_vector(6300, 16),
23111 => conv_std_logic_vector(6390, 16),
23112 => conv_std_logic_vector(6480, 16),
23113 => conv_std_logic_vector(6570, 16),
23114 => conv_std_logic_vector(6660, 16),
23115 => conv_std_logic_vector(6750, 16),
23116 => conv_std_logic_vector(6840, 16),
23117 => conv_std_logic_vector(6930, 16),
23118 => conv_std_logic_vector(7020, 16),
23119 => conv_std_logic_vector(7110, 16),
23120 => conv_std_logic_vector(7200, 16),
23121 => conv_std_logic_vector(7290, 16),
23122 => conv_std_logic_vector(7380, 16),
23123 => conv_std_logic_vector(7470, 16),
23124 => conv_std_logic_vector(7560, 16),
23125 => conv_std_logic_vector(7650, 16),
23126 => conv_std_logic_vector(7740, 16),
23127 => conv_std_logic_vector(7830, 16),
23128 => conv_std_logic_vector(7920, 16),
23129 => conv_std_logic_vector(8010, 16),
23130 => conv_std_logic_vector(8100, 16),
23131 => conv_std_logic_vector(8190, 16),
23132 => conv_std_logic_vector(8280, 16),
23133 => conv_std_logic_vector(8370, 16),
23134 => conv_std_logic_vector(8460, 16),
23135 => conv_std_logic_vector(8550, 16),
23136 => conv_std_logic_vector(8640, 16),
23137 => conv_std_logic_vector(8730, 16),
23138 => conv_std_logic_vector(8820, 16),
23139 => conv_std_logic_vector(8910, 16),
23140 => conv_std_logic_vector(9000, 16),
23141 => conv_std_logic_vector(9090, 16),
23142 => conv_std_logic_vector(9180, 16),
23143 => conv_std_logic_vector(9270, 16),
23144 => conv_std_logic_vector(9360, 16),
23145 => conv_std_logic_vector(9450, 16),
23146 => conv_std_logic_vector(9540, 16),
23147 => conv_std_logic_vector(9630, 16),
23148 => conv_std_logic_vector(9720, 16),
23149 => conv_std_logic_vector(9810, 16),
23150 => conv_std_logic_vector(9900, 16),
23151 => conv_std_logic_vector(9990, 16),
23152 => conv_std_logic_vector(10080, 16),
23153 => conv_std_logic_vector(10170, 16),
23154 => conv_std_logic_vector(10260, 16),
23155 => conv_std_logic_vector(10350, 16),
23156 => conv_std_logic_vector(10440, 16),
23157 => conv_std_logic_vector(10530, 16),
23158 => conv_std_logic_vector(10620, 16),
23159 => conv_std_logic_vector(10710, 16),
23160 => conv_std_logic_vector(10800, 16),
23161 => conv_std_logic_vector(10890, 16),
23162 => conv_std_logic_vector(10980, 16),
23163 => conv_std_logic_vector(11070, 16),
23164 => conv_std_logic_vector(11160, 16),
23165 => conv_std_logic_vector(11250, 16),
23166 => conv_std_logic_vector(11340, 16),
23167 => conv_std_logic_vector(11430, 16),
23168 => conv_std_logic_vector(11520, 16),
23169 => conv_std_logic_vector(11610, 16),
23170 => conv_std_logic_vector(11700, 16),
23171 => conv_std_logic_vector(11790, 16),
23172 => conv_std_logic_vector(11880, 16),
23173 => conv_std_logic_vector(11970, 16),
23174 => conv_std_logic_vector(12060, 16),
23175 => conv_std_logic_vector(12150, 16),
23176 => conv_std_logic_vector(12240, 16),
23177 => conv_std_logic_vector(12330, 16),
23178 => conv_std_logic_vector(12420, 16),
23179 => conv_std_logic_vector(12510, 16),
23180 => conv_std_logic_vector(12600, 16),
23181 => conv_std_logic_vector(12690, 16),
23182 => conv_std_logic_vector(12780, 16),
23183 => conv_std_logic_vector(12870, 16),
23184 => conv_std_logic_vector(12960, 16),
23185 => conv_std_logic_vector(13050, 16),
23186 => conv_std_logic_vector(13140, 16),
23187 => conv_std_logic_vector(13230, 16),
23188 => conv_std_logic_vector(13320, 16),
23189 => conv_std_logic_vector(13410, 16),
23190 => conv_std_logic_vector(13500, 16),
23191 => conv_std_logic_vector(13590, 16),
23192 => conv_std_logic_vector(13680, 16),
23193 => conv_std_logic_vector(13770, 16),
23194 => conv_std_logic_vector(13860, 16),
23195 => conv_std_logic_vector(13950, 16),
23196 => conv_std_logic_vector(14040, 16),
23197 => conv_std_logic_vector(14130, 16),
23198 => conv_std_logic_vector(14220, 16),
23199 => conv_std_logic_vector(14310, 16),
23200 => conv_std_logic_vector(14400, 16),
23201 => conv_std_logic_vector(14490, 16),
23202 => conv_std_logic_vector(14580, 16),
23203 => conv_std_logic_vector(14670, 16),
23204 => conv_std_logic_vector(14760, 16),
23205 => conv_std_logic_vector(14850, 16),
23206 => conv_std_logic_vector(14940, 16),
23207 => conv_std_logic_vector(15030, 16),
23208 => conv_std_logic_vector(15120, 16),
23209 => conv_std_logic_vector(15210, 16),
23210 => conv_std_logic_vector(15300, 16),
23211 => conv_std_logic_vector(15390, 16),
23212 => conv_std_logic_vector(15480, 16),
23213 => conv_std_logic_vector(15570, 16),
23214 => conv_std_logic_vector(15660, 16),
23215 => conv_std_logic_vector(15750, 16),
23216 => conv_std_logic_vector(15840, 16),
23217 => conv_std_logic_vector(15930, 16),
23218 => conv_std_logic_vector(16020, 16),
23219 => conv_std_logic_vector(16110, 16),
23220 => conv_std_logic_vector(16200, 16),
23221 => conv_std_logic_vector(16290, 16),
23222 => conv_std_logic_vector(16380, 16),
23223 => conv_std_logic_vector(16470, 16),
23224 => conv_std_logic_vector(16560, 16),
23225 => conv_std_logic_vector(16650, 16),
23226 => conv_std_logic_vector(16740, 16),
23227 => conv_std_logic_vector(16830, 16),
23228 => conv_std_logic_vector(16920, 16),
23229 => conv_std_logic_vector(17010, 16),
23230 => conv_std_logic_vector(17100, 16),
23231 => conv_std_logic_vector(17190, 16),
23232 => conv_std_logic_vector(17280, 16),
23233 => conv_std_logic_vector(17370, 16),
23234 => conv_std_logic_vector(17460, 16),
23235 => conv_std_logic_vector(17550, 16),
23236 => conv_std_logic_vector(17640, 16),
23237 => conv_std_logic_vector(17730, 16),
23238 => conv_std_logic_vector(17820, 16),
23239 => conv_std_logic_vector(17910, 16),
23240 => conv_std_logic_vector(18000, 16),
23241 => conv_std_logic_vector(18090, 16),
23242 => conv_std_logic_vector(18180, 16),
23243 => conv_std_logic_vector(18270, 16),
23244 => conv_std_logic_vector(18360, 16),
23245 => conv_std_logic_vector(18450, 16),
23246 => conv_std_logic_vector(18540, 16),
23247 => conv_std_logic_vector(18630, 16),
23248 => conv_std_logic_vector(18720, 16),
23249 => conv_std_logic_vector(18810, 16),
23250 => conv_std_logic_vector(18900, 16),
23251 => conv_std_logic_vector(18990, 16),
23252 => conv_std_logic_vector(19080, 16),
23253 => conv_std_logic_vector(19170, 16),
23254 => conv_std_logic_vector(19260, 16),
23255 => conv_std_logic_vector(19350, 16),
23256 => conv_std_logic_vector(19440, 16),
23257 => conv_std_logic_vector(19530, 16),
23258 => conv_std_logic_vector(19620, 16),
23259 => conv_std_logic_vector(19710, 16),
23260 => conv_std_logic_vector(19800, 16),
23261 => conv_std_logic_vector(19890, 16),
23262 => conv_std_logic_vector(19980, 16),
23263 => conv_std_logic_vector(20070, 16),
23264 => conv_std_logic_vector(20160, 16),
23265 => conv_std_logic_vector(20250, 16),
23266 => conv_std_logic_vector(20340, 16),
23267 => conv_std_logic_vector(20430, 16),
23268 => conv_std_logic_vector(20520, 16),
23269 => conv_std_logic_vector(20610, 16),
23270 => conv_std_logic_vector(20700, 16),
23271 => conv_std_logic_vector(20790, 16),
23272 => conv_std_logic_vector(20880, 16),
23273 => conv_std_logic_vector(20970, 16),
23274 => conv_std_logic_vector(21060, 16),
23275 => conv_std_logic_vector(21150, 16),
23276 => conv_std_logic_vector(21240, 16),
23277 => conv_std_logic_vector(21330, 16),
23278 => conv_std_logic_vector(21420, 16),
23279 => conv_std_logic_vector(21510, 16),
23280 => conv_std_logic_vector(21600, 16),
23281 => conv_std_logic_vector(21690, 16),
23282 => conv_std_logic_vector(21780, 16),
23283 => conv_std_logic_vector(21870, 16),
23284 => conv_std_logic_vector(21960, 16),
23285 => conv_std_logic_vector(22050, 16),
23286 => conv_std_logic_vector(22140, 16),
23287 => conv_std_logic_vector(22230, 16),
23288 => conv_std_logic_vector(22320, 16),
23289 => conv_std_logic_vector(22410, 16),
23290 => conv_std_logic_vector(22500, 16),
23291 => conv_std_logic_vector(22590, 16),
23292 => conv_std_logic_vector(22680, 16),
23293 => conv_std_logic_vector(22770, 16),
23294 => conv_std_logic_vector(22860, 16),
23295 => conv_std_logic_vector(22950, 16),
23296 => conv_std_logic_vector(0, 16),
23297 => conv_std_logic_vector(91, 16),
23298 => conv_std_logic_vector(182, 16),
23299 => conv_std_logic_vector(273, 16),
23300 => conv_std_logic_vector(364, 16),
23301 => conv_std_logic_vector(455, 16),
23302 => conv_std_logic_vector(546, 16),
23303 => conv_std_logic_vector(637, 16),
23304 => conv_std_logic_vector(728, 16),
23305 => conv_std_logic_vector(819, 16),
23306 => conv_std_logic_vector(910, 16),
23307 => conv_std_logic_vector(1001, 16),
23308 => conv_std_logic_vector(1092, 16),
23309 => conv_std_logic_vector(1183, 16),
23310 => conv_std_logic_vector(1274, 16),
23311 => conv_std_logic_vector(1365, 16),
23312 => conv_std_logic_vector(1456, 16),
23313 => conv_std_logic_vector(1547, 16),
23314 => conv_std_logic_vector(1638, 16),
23315 => conv_std_logic_vector(1729, 16),
23316 => conv_std_logic_vector(1820, 16),
23317 => conv_std_logic_vector(1911, 16),
23318 => conv_std_logic_vector(2002, 16),
23319 => conv_std_logic_vector(2093, 16),
23320 => conv_std_logic_vector(2184, 16),
23321 => conv_std_logic_vector(2275, 16),
23322 => conv_std_logic_vector(2366, 16),
23323 => conv_std_logic_vector(2457, 16),
23324 => conv_std_logic_vector(2548, 16),
23325 => conv_std_logic_vector(2639, 16),
23326 => conv_std_logic_vector(2730, 16),
23327 => conv_std_logic_vector(2821, 16),
23328 => conv_std_logic_vector(2912, 16),
23329 => conv_std_logic_vector(3003, 16),
23330 => conv_std_logic_vector(3094, 16),
23331 => conv_std_logic_vector(3185, 16),
23332 => conv_std_logic_vector(3276, 16),
23333 => conv_std_logic_vector(3367, 16),
23334 => conv_std_logic_vector(3458, 16),
23335 => conv_std_logic_vector(3549, 16),
23336 => conv_std_logic_vector(3640, 16),
23337 => conv_std_logic_vector(3731, 16),
23338 => conv_std_logic_vector(3822, 16),
23339 => conv_std_logic_vector(3913, 16),
23340 => conv_std_logic_vector(4004, 16),
23341 => conv_std_logic_vector(4095, 16),
23342 => conv_std_logic_vector(4186, 16),
23343 => conv_std_logic_vector(4277, 16),
23344 => conv_std_logic_vector(4368, 16),
23345 => conv_std_logic_vector(4459, 16),
23346 => conv_std_logic_vector(4550, 16),
23347 => conv_std_logic_vector(4641, 16),
23348 => conv_std_logic_vector(4732, 16),
23349 => conv_std_logic_vector(4823, 16),
23350 => conv_std_logic_vector(4914, 16),
23351 => conv_std_logic_vector(5005, 16),
23352 => conv_std_logic_vector(5096, 16),
23353 => conv_std_logic_vector(5187, 16),
23354 => conv_std_logic_vector(5278, 16),
23355 => conv_std_logic_vector(5369, 16),
23356 => conv_std_logic_vector(5460, 16),
23357 => conv_std_logic_vector(5551, 16),
23358 => conv_std_logic_vector(5642, 16),
23359 => conv_std_logic_vector(5733, 16),
23360 => conv_std_logic_vector(5824, 16),
23361 => conv_std_logic_vector(5915, 16),
23362 => conv_std_logic_vector(6006, 16),
23363 => conv_std_logic_vector(6097, 16),
23364 => conv_std_logic_vector(6188, 16),
23365 => conv_std_logic_vector(6279, 16),
23366 => conv_std_logic_vector(6370, 16),
23367 => conv_std_logic_vector(6461, 16),
23368 => conv_std_logic_vector(6552, 16),
23369 => conv_std_logic_vector(6643, 16),
23370 => conv_std_logic_vector(6734, 16),
23371 => conv_std_logic_vector(6825, 16),
23372 => conv_std_logic_vector(6916, 16),
23373 => conv_std_logic_vector(7007, 16),
23374 => conv_std_logic_vector(7098, 16),
23375 => conv_std_logic_vector(7189, 16),
23376 => conv_std_logic_vector(7280, 16),
23377 => conv_std_logic_vector(7371, 16),
23378 => conv_std_logic_vector(7462, 16),
23379 => conv_std_logic_vector(7553, 16),
23380 => conv_std_logic_vector(7644, 16),
23381 => conv_std_logic_vector(7735, 16),
23382 => conv_std_logic_vector(7826, 16),
23383 => conv_std_logic_vector(7917, 16),
23384 => conv_std_logic_vector(8008, 16),
23385 => conv_std_logic_vector(8099, 16),
23386 => conv_std_logic_vector(8190, 16),
23387 => conv_std_logic_vector(8281, 16),
23388 => conv_std_logic_vector(8372, 16),
23389 => conv_std_logic_vector(8463, 16),
23390 => conv_std_logic_vector(8554, 16),
23391 => conv_std_logic_vector(8645, 16),
23392 => conv_std_logic_vector(8736, 16),
23393 => conv_std_logic_vector(8827, 16),
23394 => conv_std_logic_vector(8918, 16),
23395 => conv_std_logic_vector(9009, 16),
23396 => conv_std_logic_vector(9100, 16),
23397 => conv_std_logic_vector(9191, 16),
23398 => conv_std_logic_vector(9282, 16),
23399 => conv_std_logic_vector(9373, 16),
23400 => conv_std_logic_vector(9464, 16),
23401 => conv_std_logic_vector(9555, 16),
23402 => conv_std_logic_vector(9646, 16),
23403 => conv_std_logic_vector(9737, 16),
23404 => conv_std_logic_vector(9828, 16),
23405 => conv_std_logic_vector(9919, 16),
23406 => conv_std_logic_vector(10010, 16),
23407 => conv_std_logic_vector(10101, 16),
23408 => conv_std_logic_vector(10192, 16),
23409 => conv_std_logic_vector(10283, 16),
23410 => conv_std_logic_vector(10374, 16),
23411 => conv_std_logic_vector(10465, 16),
23412 => conv_std_logic_vector(10556, 16),
23413 => conv_std_logic_vector(10647, 16),
23414 => conv_std_logic_vector(10738, 16),
23415 => conv_std_logic_vector(10829, 16),
23416 => conv_std_logic_vector(10920, 16),
23417 => conv_std_logic_vector(11011, 16),
23418 => conv_std_logic_vector(11102, 16),
23419 => conv_std_logic_vector(11193, 16),
23420 => conv_std_logic_vector(11284, 16),
23421 => conv_std_logic_vector(11375, 16),
23422 => conv_std_logic_vector(11466, 16),
23423 => conv_std_logic_vector(11557, 16),
23424 => conv_std_logic_vector(11648, 16),
23425 => conv_std_logic_vector(11739, 16),
23426 => conv_std_logic_vector(11830, 16),
23427 => conv_std_logic_vector(11921, 16),
23428 => conv_std_logic_vector(12012, 16),
23429 => conv_std_logic_vector(12103, 16),
23430 => conv_std_logic_vector(12194, 16),
23431 => conv_std_logic_vector(12285, 16),
23432 => conv_std_logic_vector(12376, 16),
23433 => conv_std_logic_vector(12467, 16),
23434 => conv_std_logic_vector(12558, 16),
23435 => conv_std_logic_vector(12649, 16),
23436 => conv_std_logic_vector(12740, 16),
23437 => conv_std_logic_vector(12831, 16),
23438 => conv_std_logic_vector(12922, 16),
23439 => conv_std_logic_vector(13013, 16),
23440 => conv_std_logic_vector(13104, 16),
23441 => conv_std_logic_vector(13195, 16),
23442 => conv_std_logic_vector(13286, 16),
23443 => conv_std_logic_vector(13377, 16),
23444 => conv_std_logic_vector(13468, 16),
23445 => conv_std_logic_vector(13559, 16),
23446 => conv_std_logic_vector(13650, 16),
23447 => conv_std_logic_vector(13741, 16),
23448 => conv_std_logic_vector(13832, 16),
23449 => conv_std_logic_vector(13923, 16),
23450 => conv_std_logic_vector(14014, 16),
23451 => conv_std_logic_vector(14105, 16),
23452 => conv_std_logic_vector(14196, 16),
23453 => conv_std_logic_vector(14287, 16),
23454 => conv_std_logic_vector(14378, 16),
23455 => conv_std_logic_vector(14469, 16),
23456 => conv_std_logic_vector(14560, 16),
23457 => conv_std_logic_vector(14651, 16),
23458 => conv_std_logic_vector(14742, 16),
23459 => conv_std_logic_vector(14833, 16),
23460 => conv_std_logic_vector(14924, 16),
23461 => conv_std_logic_vector(15015, 16),
23462 => conv_std_logic_vector(15106, 16),
23463 => conv_std_logic_vector(15197, 16),
23464 => conv_std_logic_vector(15288, 16),
23465 => conv_std_logic_vector(15379, 16),
23466 => conv_std_logic_vector(15470, 16),
23467 => conv_std_logic_vector(15561, 16),
23468 => conv_std_logic_vector(15652, 16),
23469 => conv_std_logic_vector(15743, 16),
23470 => conv_std_logic_vector(15834, 16),
23471 => conv_std_logic_vector(15925, 16),
23472 => conv_std_logic_vector(16016, 16),
23473 => conv_std_logic_vector(16107, 16),
23474 => conv_std_logic_vector(16198, 16),
23475 => conv_std_logic_vector(16289, 16),
23476 => conv_std_logic_vector(16380, 16),
23477 => conv_std_logic_vector(16471, 16),
23478 => conv_std_logic_vector(16562, 16),
23479 => conv_std_logic_vector(16653, 16),
23480 => conv_std_logic_vector(16744, 16),
23481 => conv_std_logic_vector(16835, 16),
23482 => conv_std_logic_vector(16926, 16),
23483 => conv_std_logic_vector(17017, 16),
23484 => conv_std_logic_vector(17108, 16),
23485 => conv_std_logic_vector(17199, 16),
23486 => conv_std_logic_vector(17290, 16),
23487 => conv_std_logic_vector(17381, 16),
23488 => conv_std_logic_vector(17472, 16),
23489 => conv_std_logic_vector(17563, 16),
23490 => conv_std_logic_vector(17654, 16),
23491 => conv_std_logic_vector(17745, 16),
23492 => conv_std_logic_vector(17836, 16),
23493 => conv_std_logic_vector(17927, 16),
23494 => conv_std_logic_vector(18018, 16),
23495 => conv_std_logic_vector(18109, 16),
23496 => conv_std_logic_vector(18200, 16),
23497 => conv_std_logic_vector(18291, 16),
23498 => conv_std_logic_vector(18382, 16),
23499 => conv_std_logic_vector(18473, 16),
23500 => conv_std_logic_vector(18564, 16),
23501 => conv_std_logic_vector(18655, 16),
23502 => conv_std_logic_vector(18746, 16),
23503 => conv_std_logic_vector(18837, 16),
23504 => conv_std_logic_vector(18928, 16),
23505 => conv_std_logic_vector(19019, 16),
23506 => conv_std_logic_vector(19110, 16),
23507 => conv_std_logic_vector(19201, 16),
23508 => conv_std_logic_vector(19292, 16),
23509 => conv_std_logic_vector(19383, 16),
23510 => conv_std_logic_vector(19474, 16),
23511 => conv_std_logic_vector(19565, 16),
23512 => conv_std_logic_vector(19656, 16),
23513 => conv_std_logic_vector(19747, 16),
23514 => conv_std_logic_vector(19838, 16),
23515 => conv_std_logic_vector(19929, 16),
23516 => conv_std_logic_vector(20020, 16),
23517 => conv_std_logic_vector(20111, 16),
23518 => conv_std_logic_vector(20202, 16),
23519 => conv_std_logic_vector(20293, 16),
23520 => conv_std_logic_vector(20384, 16),
23521 => conv_std_logic_vector(20475, 16),
23522 => conv_std_logic_vector(20566, 16),
23523 => conv_std_logic_vector(20657, 16),
23524 => conv_std_logic_vector(20748, 16),
23525 => conv_std_logic_vector(20839, 16),
23526 => conv_std_logic_vector(20930, 16),
23527 => conv_std_logic_vector(21021, 16),
23528 => conv_std_logic_vector(21112, 16),
23529 => conv_std_logic_vector(21203, 16),
23530 => conv_std_logic_vector(21294, 16),
23531 => conv_std_logic_vector(21385, 16),
23532 => conv_std_logic_vector(21476, 16),
23533 => conv_std_logic_vector(21567, 16),
23534 => conv_std_logic_vector(21658, 16),
23535 => conv_std_logic_vector(21749, 16),
23536 => conv_std_logic_vector(21840, 16),
23537 => conv_std_logic_vector(21931, 16),
23538 => conv_std_logic_vector(22022, 16),
23539 => conv_std_logic_vector(22113, 16),
23540 => conv_std_logic_vector(22204, 16),
23541 => conv_std_logic_vector(22295, 16),
23542 => conv_std_logic_vector(22386, 16),
23543 => conv_std_logic_vector(22477, 16),
23544 => conv_std_logic_vector(22568, 16),
23545 => conv_std_logic_vector(22659, 16),
23546 => conv_std_logic_vector(22750, 16),
23547 => conv_std_logic_vector(22841, 16),
23548 => conv_std_logic_vector(22932, 16),
23549 => conv_std_logic_vector(23023, 16),
23550 => conv_std_logic_vector(23114, 16),
23551 => conv_std_logic_vector(23205, 16),
23552 => conv_std_logic_vector(0, 16),
23553 => conv_std_logic_vector(92, 16),
23554 => conv_std_logic_vector(184, 16),
23555 => conv_std_logic_vector(276, 16),
23556 => conv_std_logic_vector(368, 16),
23557 => conv_std_logic_vector(460, 16),
23558 => conv_std_logic_vector(552, 16),
23559 => conv_std_logic_vector(644, 16),
23560 => conv_std_logic_vector(736, 16),
23561 => conv_std_logic_vector(828, 16),
23562 => conv_std_logic_vector(920, 16),
23563 => conv_std_logic_vector(1012, 16),
23564 => conv_std_logic_vector(1104, 16),
23565 => conv_std_logic_vector(1196, 16),
23566 => conv_std_logic_vector(1288, 16),
23567 => conv_std_logic_vector(1380, 16),
23568 => conv_std_logic_vector(1472, 16),
23569 => conv_std_logic_vector(1564, 16),
23570 => conv_std_logic_vector(1656, 16),
23571 => conv_std_logic_vector(1748, 16),
23572 => conv_std_logic_vector(1840, 16),
23573 => conv_std_logic_vector(1932, 16),
23574 => conv_std_logic_vector(2024, 16),
23575 => conv_std_logic_vector(2116, 16),
23576 => conv_std_logic_vector(2208, 16),
23577 => conv_std_logic_vector(2300, 16),
23578 => conv_std_logic_vector(2392, 16),
23579 => conv_std_logic_vector(2484, 16),
23580 => conv_std_logic_vector(2576, 16),
23581 => conv_std_logic_vector(2668, 16),
23582 => conv_std_logic_vector(2760, 16),
23583 => conv_std_logic_vector(2852, 16),
23584 => conv_std_logic_vector(2944, 16),
23585 => conv_std_logic_vector(3036, 16),
23586 => conv_std_logic_vector(3128, 16),
23587 => conv_std_logic_vector(3220, 16),
23588 => conv_std_logic_vector(3312, 16),
23589 => conv_std_logic_vector(3404, 16),
23590 => conv_std_logic_vector(3496, 16),
23591 => conv_std_logic_vector(3588, 16),
23592 => conv_std_logic_vector(3680, 16),
23593 => conv_std_logic_vector(3772, 16),
23594 => conv_std_logic_vector(3864, 16),
23595 => conv_std_logic_vector(3956, 16),
23596 => conv_std_logic_vector(4048, 16),
23597 => conv_std_logic_vector(4140, 16),
23598 => conv_std_logic_vector(4232, 16),
23599 => conv_std_logic_vector(4324, 16),
23600 => conv_std_logic_vector(4416, 16),
23601 => conv_std_logic_vector(4508, 16),
23602 => conv_std_logic_vector(4600, 16),
23603 => conv_std_logic_vector(4692, 16),
23604 => conv_std_logic_vector(4784, 16),
23605 => conv_std_logic_vector(4876, 16),
23606 => conv_std_logic_vector(4968, 16),
23607 => conv_std_logic_vector(5060, 16),
23608 => conv_std_logic_vector(5152, 16),
23609 => conv_std_logic_vector(5244, 16),
23610 => conv_std_logic_vector(5336, 16),
23611 => conv_std_logic_vector(5428, 16),
23612 => conv_std_logic_vector(5520, 16),
23613 => conv_std_logic_vector(5612, 16),
23614 => conv_std_logic_vector(5704, 16),
23615 => conv_std_logic_vector(5796, 16),
23616 => conv_std_logic_vector(5888, 16),
23617 => conv_std_logic_vector(5980, 16),
23618 => conv_std_logic_vector(6072, 16),
23619 => conv_std_logic_vector(6164, 16),
23620 => conv_std_logic_vector(6256, 16),
23621 => conv_std_logic_vector(6348, 16),
23622 => conv_std_logic_vector(6440, 16),
23623 => conv_std_logic_vector(6532, 16),
23624 => conv_std_logic_vector(6624, 16),
23625 => conv_std_logic_vector(6716, 16),
23626 => conv_std_logic_vector(6808, 16),
23627 => conv_std_logic_vector(6900, 16),
23628 => conv_std_logic_vector(6992, 16),
23629 => conv_std_logic_vector(7084, 16),
23630 => conv_std_logic_vector(7176, 16),
23631 => conv_std_logic_vector(7268, 16),
23632 => conv_std_logic_vector(7360, 16),
23633 => conv_std_logic_vector(7452, 16),
23634 => conv_std_logic_vector(7544, 16),
23635 => conv_std_logic_vector(7636, 16),
23636 => conv_std_logic_vector(7728, 16),
23637 => conv_std_logic_vector(7820, 16),
23638 => conv_std_logic_vector(7912, 16),
23639 => conv_std_logic_vector(8004, 16),
23640 => conv_std_logic_vector(8096, 16),
23641 => conv_std_logic_vector(8188, 16),
23642 => conv_std_logic_vector(8280, 16),
23643 => conv_std_logic_vector(8372, 16),
23644 => conv_std_logic_vector(8464, 16),
23645 => conv_std_logic_vector(8556, 16),
23646 => conv_std_logic_vector(8648, 16),
23647 => conv_std_logic_vector(8740, 16),
23648 => conv_std_logic_vector(8832, 16),
23649 => conv_std_logic_vector(8924, 16),
23650 => conv_std_logic_vector(9016, 16),
23651 => conv_std_logic_vector(9108, 16),
23652 => conv_std_logic_vector(9200, 16),
23653 => conv_std_logic_vector(9292, 16),
23654 => conv_std_logic_vector(9384, 16),
23655 => conv_std_logic_vector(9476, 16),
23656 => conv_std_logic_vector(9568, 16),
23657 => conv_std_logic_vector(9660, 16),
23658 => conv_std_logic_vector(9752, 16),
23659 => conv_std_logic_vector(9844, 16),
23660 => conv_std_logic_vector(9936, 16),
23661 => conv_std_logic_vector(10028, 16),
23662 => conv_std_logic_vector(10120, 16),
23663 => conv_std_logic_vector(10212, 16),
23664 => conv_std_logic_vector(10304, 16),
23665 => conv_std_logic_vector(10396, 16),
23666 => conv_std_logic_vector(10488, 16),
23667 => conv_std_logic_vector(10580, 16),
23668 => conv_std_logic_vector(10672, 16),
23669 => conv_std_logic_vector(10764, 16),
23670 => conv_std_logic_vector(10856, 16),
23671 => conv_std_logic_vector(10948, 16),
23672 => conv_std_logic_vector(11040, 16),
23673 => conv_std_logic_vector(11132, 16),
23674 => conv_std_logic_vector(11224, 16),
23675 => conv_std_logic_vector(11316, 16),
23676 => conv_std_logic_vector(11408, 16),
23677 => conv_std_logic_vector(11500, 16),
23678 => conv_std_logic_vector(11592, 16),
23679 => conv_std_logic_vector(11684, 16),
23680 => conv_std_logic_vector(11776, 16),
23681 => conv_std_logic_vector(11868, 16),
23682 => conv_std_logic_vector(11960, 16),
23683 => conv_std_logic_vector(12052, 16),
23684 => conv_std_logic_vector(12144, 16),
23685 => conv_std_logic_vector(12236, 16),
23686 => conv_std_logic_vector(12328, 16),
23687 => conv_std_logic_vector(12420, 16),
23688 => conv_std_logic_vector(12512, 16),
23689 => conv_std_logic_vector(12604, 16),
23690 => conv_std_logic_vector(12696, 16),
23691 => conv_std_logic_vector(12788, 16),
23692 => conv_std_logic_vector(12880, 16),
23693 => conv_std_logic_vector(12972, 16),
23694 => conv_std_logic_vector(13064, 16),
23695 => conv_std_logic_vector(13156, 16),
23696 => conv_std_logic_vector(13248, 16),
23697 => conv_std_logic_vector(13340, 16),
23698 => conv_std_logic_vector(13432, 16),
23699 => conv_std_logic_vector(13524, 16),
23700 => conv_std_logic_vector(13616, 16),
23701 => conv_std_logic_vector(13708, 16),
23702 => conv_std_logic_vector(13800, 16),
23703 => conv_std_logic_vector(13892, 16),
23704 => conv_std_logic_vector(13984, 16),
23705 => conv_std_logic_vector(14076, 16),
23706 => conv_std_logic_vector(14168, 16),
23707 => conv_std_logic_vector(14260, 16),
23708 => conv_std_logic_vector(14352, 16),
23709 => conv_std_logic_vector(14444, 16),
23710 => conv_std_logic_vector(14536, 16),
23711 => conv_std_logic_vector(14628, 16),
23712 => conv_std_logic_vector(14720, 16),
23713 => conv_std_logic_vector(14812, 16),
23714 => conv_std_logic_vector(14904, 16),
23715 => conv_std_logic_vector(14996, 16),
23716 => conv_std_logic_vector(15088, 16),
23717 => conv_std_logic_vector(15180, 16),
23718 => conv_std_logic_vector(15272, 16),
23719 => conv_std_logic_vector(15364, 16),
23720 => conv_std_logic_vector(15456, 16),
23721 => conv_std_logic_vector(15548, 16),
23722 => conv_std_logic_vector(15640, 16),
23723 => conv_std_logic_vector(15732, 16),
23724 => conv_std_logic_vector(15824, 16),
23725 => conv_std_logic_vector(15916, 16),
23726 => conv_std_logic_vector(16008, 16),
23727 => conv_std_logic_vector(16100, 16),
23728 => conv_std_logic_vector(16192, 16),
23729 => conv_std_logic_vector(16284, 16),
23730 => conv_std_logic_vector(16376, 16),
23731 => conv_std_logic_vector(16468, 16),
23732 => conv_std_logic_vector(16560, 16),
23733 => conv_std_logic_vector(16652, 16),
23734 => conv_std_logic_vector(16744, 16),
23735 => conv_std_logic_vector(16836, 16),
23736 => conv_std_logic_vector(16928, 16),
23737 => conv_std_logic_vector(17020, 16),
23738 => conv_std_logic_vector(17112, 16),
23739 => conv_std_logic_vector(17204, 16),
23740 => conv_std_logic_vector(17296, 16),
23741 => conv_std_logic_vector(17388, 16),
23742 => conv_std_logic_vector(17480, 16),
23743 => conv_std_logic_vector(17572, 16),
23744 => conv_std_logic_vector(17664, 16),
23745 => conv_std_logic_vector(17756, 16),
23746 => conv_std_logic_vector(17848, 16),
23747 => conv_std_logic_vector(17940, 16),
23748 => conv_std_logic_vector(18032, 16),
23749 => conv_std_logic_vector(18124, 16),
23750 => conv_std_logic_vector(18216, 16),
23751 => conv_std_logic_vector(18308, 16),
23752 => conv_std_logic_vector(18400, 16),
23753 => conv_std_logic_vector(18492, 16),
23754 => conv_std_logic_vector(18584, 16),
23755 => conv_std_logic_vector(18676, 16),
23756 => conv_std_logic_vector(18768, 16),
23757 => conv_std_logic_vector(18860, 16),
23758 => conv_std_logic_vector(18952, 16),
23759 => conv_std_logic_vector(19044, 16),
23760 => conv_std_logic_vector(19136, 16),
23761 => conv_std_logic_vector(19228, 16),
23762 => conv_std_logic_vector(19320, 16),
23763 => conv_std_logic_vector(19412, 16),
23764 => conv_std_logic_vector(19504, 16),
23765 => conv_std_logic_vector(19596, 16),
23766 => conv_std_logic_vector(19688, 16),
23767 => conv_std_logic_vector(19780, 16),
23768 => conv_std_logic_vector(19872, 16),
23769 => conv_std_logic_vector(19964, 16),
23770 => conv_std_logic_vector(20056, 16),
23771 => conv_std_logic_vector(20148, 16),
23772 => conv_std_logic_vector(20240, 16),
23773 => conv_std_logic_vector(20332, 16),
23774 => conv_std_logic_vector(20424, 16),
23775 => conv_std_logic_vector(20516, 16),
23776 => conv_std_logic_vector(20608, 16),
23777 => conv_std_logic_vector(20700, 16),
23778 => conv_std_logic_vector(20792, 16),
23779 => conv_std_logic_vector(20884, 16),
23780 => conv_std_logic_vector(20976, 16),
23781 => conv_std_logic_vector(21068, 16),
23782 => conv_std_logic_vector(21160, 16),
23783 => conv_std_logic_vector(21252, 16),
23784 => conv_std_logic_vector(21344, 16),
23785 => conv_std_logic_vector(21436, 16),
23786 => conv_std_logic_vector(21528, 16),
23787 => conv_std_logic_vector(21620, 16),
23788 => conv_std_logic_vector(21712, 16),
23789 => conv_std_logic_vector(21804, 16),
23790 => conv_std_logic_vector(21896, 16),
23791 => conv_std_logic_vector(21988, 16),
23792 => conv_std_logic_vector(22080, 16),
23793 => conv_std_logic_vector(22172, 16),
23794 => conv_std_logic_vector(22264, 16),
23795 => conv_std_logic_vector(22356, 16),
23796 => conv_std_logic_vector(22448, 16),
23797 => conv_std_logic_vector(22540, 16),
23798 => conv_std_logic_vector(22632, 16),
23799 => conv_std_logic_vector(22724, 16),
23800 => conv_std_logic_vector(22816, 16),
23801 => conv_std_logic_vector(22908, 16),
23802 => conv_std_logic_vector(23000, 16),
23803 => conv_std_logic_vector(23092, 16),
23804 => conv_std_logic_vector(23184, 16),
23805 => conv_std_logic_vector(23276, 16),
23806 => conv_std_logic_vector(23368, 16),
23807 => conv_std_logic_vector(23460, 16),
23808 => conv_std_logic_vector(0, 16),
23809 => conv_std_logic_vector(93, 16),
23810 => conv_std_logic_vector(186, 16),
23811 => conv_std_logic_vector(279, 16),
23812 => conv_std_logic_vector(372, 16),
23813 => conv_std_logic_vector(465, 16),
23814 => conv_std_logic_vector(558, 16),
23815 => conv_std_logic_vector(651, 16),
23816 => conv_std_logic_vector(744, 16),
23817 => conv_std_logic_vector(837, 16),
23818 => conv_std_logic_vector(930, 16),
23819 => conv_std_logic_vector(1023, 16),
23820 => conv_std_logic_vector(1116, 16),
23821 => conv_std_logic_vector(1209, 16),
23822 => conv_std_logic_vector(1302, 16),
23823 => conv_std_logic_vector(1395, 16),
23824 => conv_std_logic_vector(1488, 16),
23825 => conv_std_logic_vector(1581, 16),
23826 => conv_std_logic_vector(1674, 16),
23827 => conv_std_logic_vector(1767, 16),
23828 => conv_std_logic_vector(1860, 16),
23829 => conv_std_logic_vector(1953, 16),
23830 => conv_std_logic_vector(2046, 16),
23831 => conv_std_logic_vector(2139, 16),
23832 => conv_std_logic_vector(2232, 16),
23833 => conv_std_logic_vector(2325, 16),
23834 => conv_std_logic_vector(2418, 16),
23835 => conv_std_logic_vector(2511, 16),
23836 => conv_std_logic_vector(2604, 16),
23837 => conv_std_logic_vector(2697, 16),
23838 => conv_std_logic_vector(2790, 16),
23839 => conv_std_logic_vector(2883, 16),
23840 => conv_std_logic_vector(2976, 16),
23841 => conv_std_logic_vector(3069, 16),
23842 => conv_std_logic_vector(3162, 16),
23843 => conv_std_logic_vector(3255, 16),
23844 => conv_std_logic_vector(3348, 16),
23845 => conv_std_logic_vector(3441, 16),
23846 => conv_std_logic_vector(3534, 16),
23847 => conv_std_logic_vector(3627, 16),
23848 => conv_std_logic_vector(3720, 16),
23849 => conv_std_logic_vector(3813, 16),
23850 => conv_std_logic_vector(3906, 16),
23851 => conv_std_logic_vector(3999, 16),
23852 => conv_std_logic_vector(4092, 16),
23853 => conv_std_logic_vector(4185, 16),
23854 => conv_std_logic_vector(4278, 16),
23855 => conv_std_logic_vector(4371, 16),
23856 => conv_std_logic_vector(4464, 16),
23857 => conv_std_logic_vector(4557, 16),
23858 => conv_std_logic_vector(4650, 16),
23859 => conv_std_logic_vector(4743, 16),
23860 => conv_std_logic_vector(4836, 16),
23861 => conv_std_logic_vector(4929, 16),
23862 => conv_std_logic_vector(5022, 16),
23863 => conv_std_logic_vector(5115, 16),
23864 => conv_std_logic_vector(5208, 16),
23865 => conv_std_logic_vector(5301, 16),
23866 => conv_std_logic_vector(5394, 16),
23867 => conv_std_logic_vector(5487, 16),
23868 => conv_std_logic_vector(5580, 16),
23869 => conv_std_logic_vector(5673, 16),
23870 => conv_std_logic_vector(5766, 16),
23871 => conv_std_logic_vector(5859, 16),
23872 => conv_std_logic_vector(5952, 16),
23873 => conv_std_logic_vector(6045, 16),
23874 => conv_std_logic_vector(6138, 16),
23875 => conv_std_logic_vector(6231, 16),
23876 => conv_std_logic_vector(6324, 16),
23877 => conv_std_logic_vector(6417, 16),
23878 => conv_std_logic_vector(6510, 16),
23879 => conv_std_logic_vector(6603, 16),
23880 => conv_std_logic_vector(6696, 16),
23881 => conv_std_logic_vector(6789, 16),
23882 => conv_std_logic_vector(6882, 16),
23883 => conv_std_logic_vector(6975, 16),
23884 => conv_std_logic_vector(7068, 16),
23885 => conv_std_logic_vector(7161, 16),
23886 => conv_std_logic_vector(7254, 16),
23887 => conv_std_logic_vector(7347, 16),
23888 => conv_std_logic_vector(7440, 16),
23889 => conv_std_logic_vector(7533, 16),
23890 => conv_std_logic_vector(7626, 16),
23891 => conv_std_logic_vector(7719, 16),
23892 => conv_std_logic_vector(7812, 16),
23893 => conv_std_logic_vector(7905, 16),
23894 => conv_std_logic_vector(7998, 16),
23895 => conv_std_logic_vector(8091, 16),
23896 => conv_std_logic_vector(8184, 16),
23897 => conv_std_logic_vector(8277, 16),
23898 => conv_std_logic_vector(8370, 16),
23899 => conv_std_logic_vector(8463, 16),
23900 => conv_std_logic_vector(8556, 16),
23901 => conv_std_logic_vector(8649, 16),
23902 => conv_std_logic_vector(8742, 16),
23903 => conv_std_logic_vector(8835, 16),
23904 => conv_std_logic_vector(8928, 16),
23905 => conv_std_logic_vector(9021, 16),
23906 => conv_std_logic_vector(9114, 16),
23907 => conv_std_logic_vector(9207, 16),
23908 => conv_std_logic_vector(9300, 16),
23909 => conv_std_logic_vector(9393, 16),
23910 => conv_std_logic_vector(9486, 16),
23911 => conv_std_logic_vector(9579, 16),
23912 => conv_std_logic_vector(9672, 16),
23913 => conv_std_logic_vector(9765, 16),
23914 => conv_std_logic_vector(9858, 16),
23915 => conv_std_logic_vector(9951, 16),
23916 => conv_std_logic_vector(10044, 16),
23917 => conv_std_logic_vector(10137, 16),
23918 => conv_std_logic_vector(10230, 16),
23919 => conv_std_logic_vector(10323, 16),
23920 => conv_std_logic_vector(10416, 16),
23921 => conv_std_logic_vector(10509, 16),
23922 => conv_std_logic_vector(10602, 16),
23923 => conv_std_logic_vector(10695, 16),
23924 => conv_std_logic_vector(10788, 16),
23925 => conv_std_logic_vector(10881, 16),
23926 => conv_std_logic_vector(10974, 16),
23927 => conv_std_logic_vector(11067, 16),
23928 => conv_std_logic_vector(11160, 16),
23929 => conv_std_logic_vector(11253, 16),
23930 => conv_std_logic_vector(11346, 16),
23931 => conv_std_logic_vector(11439, 16),
23932 => conv_std_logic_vector(11532, 16),
23933 => conv_std_logic_vector(11625, 16),
23934 => conv_std_logic_vector(11718, 16),
23935 => conv_std_logic_vector(11811, 16),
23936 => conv_std_logic_vector(11904, 16),
23937 => conv_std_logic_vector(11997, 16),
23938 => conv_std_logic_vector(12090, 16),
23939 => conv_std_logic_vector(12183, 16),
23940 => conv_std_logic_vector(12276, 16),
23941 => conv_std_logic_vector(12369, 16),
23942 => conv_std_logic_vector(12462, 16),
23943 => conv_std_logic_vector(12555, 16),
23944 => conv_std_logic_vector(12648, 16),
23945 => conv_std_logic_vector(12741, 16),
23946 => conv_std_logic_vector(12834, 16),
23947 => conv_std_logic_vector(12927, 16),
23948 => conv_std_logic_vector(13020, 16),
23949 => conv_std_logic_vector(13113, 16),
23950 => conv_std_logic_vector(13206, 16),
23951 => conv_std_logic_vector(13299, 16),
23952 => conv_std_logic_vector(13392, 16),
23953 => conv_std_logic_vector(13485, 16),
23954 => conv_std_logic_vector(13578, 16),
23955 => conv_std_logic_vector(13671, 16),
23956 => conv_std_logic_vector(13764, 16),
23957 => conv_std_logic_vector(13857, 16),
23958 => conv_std_logic_vector(13950, 16),
23959 => conv_std_logic_vector(14043, 16),
23960 => conv_std_logic_vector(14136, 16),
23961 => conv_std_logic_vector(14229, 16),
23962 => conv_std_logic_vector(14322, 16),
23963 => conv_std_logic_vector(14415, 16),
23964 => conv_std_logic_vector(14508, 16),
23965 => conv_std_logic_vector(14601, 16),
23966 => conv_std_logic_vector(14694, 16),
23967 => conv_std_logic_vector(14787, 16),
23968 => conv_std_logic_vector(14880, 16),
23969 => conv_std_logic_vector(14973, 16),
23970 => conv_std_logic_vector(15066, 16),
23971 => conv_std_logic_vector(15159, 16),
23972 => conv_std_logic_vector(15252, 16),
23973 => conv_std_logic_vector(15345, 16),
23974 => conv_std_logic_vector(15438, 16),
23975 => conv_std_logic_vector(15531, 16),
23976 => conv_std_logic_vector(15624, 16),
23977 => conv_std_logic_vector(15717, 16),
23978 => conv_std_logic_vector(15810, 16),
23979 => conv_std_logic_vector(15903, 16),
23980 => conv_std_logic_vector(15996, 16),
23981 => conv_std_logic_vector(16089, 16),
23982 => conv_std_logic_vector(16182, 16),
23983 => conv_std_logic_vector(16275, 16),
23984 => conv_std_logic_vector(16368, 16),
23985 => conv_std_logic_vector(16461, 16),
23986 => conv_std_logic_vector(16554, 16),
23987 => conv_std_logic_vector(16647, 16),
23988 => conv_std_logic_vector(16740, 16),
23989 => conv_std_logic_vector(16833, 16),
23990 => conv_std_logic_vector(16926, 16),
23991 => conv_std_logic_vector(17019, 16),
23992 => conv_std_logic_vector(17112, 16),
23993 => conv_std_logic_vector(17205, 16),
23994 => conv_std_logic_vector(17298, 16),
23995 => conv_std_logic_vector(17391, 16),
23996 => conv_std_logic_vector(17484, 16),
23997 => conv_std_logic_vector(17577, 16),
23998 => conv_std_logic_vector(17670, 16),
23999 => conv_std_logic_vector(17763, 16),
24000 => conv_std_logic_vector(17856, 16),
24001 => conv_std_logic_vector(17949, 16),
24002 => conv_std_logic_vector(18042, 16),
24003 => conv_std_logic_vector(18135, 16),
24004 => conv_std_logic_vector(18228, 16),
24005 => conv_std_logic_vector(18321, 16),
24006 => conv_std_logic_vector(18414, 16),
24007 => conv_std_logic_vector(18507, 16),
24008 => conv_std_logic_vector(18600, 16),
24009 => conv_std_logic_vector(18693, 16),
24010 => conv_std_logic_vector(18786, 16),
24011 => conv_std_logic_vector(18879, 16),
24012 => conv_std_logic_vector(18972, 16),
24013 => conv_std_logic_vector(19065, 16),
24014 => conv_std_logic_vector(19158, 16),
24015 => conv_std_logic_vector(19251, 16),
24016 => conv_std_logic_vector(19344, 16),
24017 => conv_std_logic_vector(19437, 16),
24018 => conv_std_logic_vector(19530, 16),
24019 => conv_std_logic_vector(19623, 16),
24020 => conv_std_logic_vector(19716, 16),
24021 => conv_std_logic_vector(19809, 16),
24022 => conv_std_logic_vector(19902, 16),
24023 => conv_std_logic_vector(19995, 16),
24024 => conv_std_logic_vector(20088, 16),
24025 => conv_std_logic_vector(20181, 16),
24026 => conv_std_logic_vector(20274, 16),
24027 => conv_std_logic_vector(20367, 16),
24028 => conv_std_logic_vector(20460, 16),
24029 => conv_std_logic_vector(20553, 16),
24030 => conv_std_logic_vector(20646, 16),
24031 => conv_std_logic_vector(20739, 16),
24032 => conv_std_logic_vector(20832, 16),
24033 => conv_std_logic_vector(20925, 16),
24034 => conv_std_logic_vector(21018, 16),
24035 => conv_std_logic_vector(21111, 16),
24036 => conv_std_logic_vector(21204, 16),
24037 => conv_std_logic_vector(21297, 16),
24038 => conv_std_logic_vector(21390, 16),
24039 => conv_std_logic_vector(21483, 16),
24040 => conv_std_logic_vector(21576, 16),
24041 => conv_std_logic_vector(21669, 16),
24042 => conv_std_logic_vector(21762, 16),
24043 => conv_std_logic_vector(21855, 16),
24044 => conv_std_logic_vector(21948, 16),
24045 => conv_std_logic_vector(22041, 16),
24046 => conv_std_logic_vector(22134, 16),
24047 => conv_std_logic_vector(22227, 16),
24048 => conv_std_logic_vector(22320, 16),
24049 => conv_std_logic_vector(22413, 16),
24050 => conv_std_logic_vector(22506, 16),
24051 => conv_std_logic_vector(22599, 16),
24052 => conv_std_logic_vector(22692, 16),
24053 => conv_std_logic_vector(22785, 16),
24054 => conv_std_logic_vector(22878, 16),
24055 => conv_std_logic_vector(22971, 16),
24056 => conv_std_logic_vector(23064, 16),
24057 => conv_std_logic_vector(23157, 16),
24058 => conv_std_logic_vector(23250, 16),
24059 => conv_std_logic_vector(23343, 16),
24060 => conv_std_logic_vector(23436, 16),
24061 => conv_std_logic_vector(23529, 16),
24062 => conv_std_logic_vector(23622, 16),
24063 => conv_std_logic_vector(23715, 16),
24064 => conv_std_logic_vector(0, 16),
24065 => conv_std_logic_vector(94, 16),
24066 => conv_std_logic_vector(188, 16),
24067 => conv_std_logic_vector(282, 16),
24068 => conv_std_logic_vector(376, 16),
24069 => conv_std_logic_vector(470, 16),
24070 => conv_std_logic_vector(564, 16),
24071 => conv_std_logic_vector(658, 16),
24072 => conv_std_logic_vector(752, 16),
24073 => conv_std_logic_vector(846, 16),
24074 => conv_std_logic_vector(940, 16),
24075 => conv_std_logic_vector(1034, 16),
24076 => conv_std_logic_vector(1128, 16),
24077 => conv_std_logic_vector(1222, 16),
24078 => conv_std_logic_vector(1316, 16),
24079 => conv_std_logic_vector(1410, 16),
24080 => conv_std_logic_vector(1504, 16),
24081 => conv_std_logic_vector(1598, 16),
24082 => conv_std_logic_vector(1692, 16),
24083 => conv_std_logic_vector(1786, 16),
24084 => conv_std_logic_vector(1880, 16),
24085 => conv_std_logic_vector(1974, 16),
24086 => conv_std_logic_vector(2068, 16),
24087 => conv_std_logic_vector(2162, 16),
24088 => conv_std_logic_vector(2256, 16),
24089 => conv_std_logic_vector(2350, 16),
24090 => conv_std_logic_vector(2444, 16),
24091 => conv_std_logic_vector(2538, 16),
24092 => conv_std_logic_vector(2632, 16),
24093 => conv_std_logic_vector(2726, 16),
24094 => conv_std_logic_vector(2820, 16),
24095 => conv_std_logic_vector(2914, 16),
24096 => conv_std_logic_vector(3008, 16),
24097 => conv_std_logic_vector(3102, 16),
24098 => conv_std_logic_vector(3196, 16),
24099 => conv_std_logic_vector(3290, 16),
24100 => conv_std_logic_vector(3384, 16),
24101 => conv_std_logic_vector(3478, 16),
24102 => conv_std_logic_vector(3572, 16),
24103 => conv_std_logic_vector(3666, 16),
24104 => conv_std_logic_vector(3760, 16),
24105 => conv_std_logic_vector(3854, 16),
24106 => conv_std_logic_vector(3948, 16),
24107 => conv_std_logic_vector(4042, 16),
24108 => conv_std_logic_vector(4136, 16),
24109 => conv_std_logic_vector(4230, 16),
24110 => conv_std_logic_vector(4324, 16),
24111 => conv_std_logic_vector(4418, 16),
24112 => conv_std_logic_vector(4512, 16),
24113 => conv_std_logic_vector(4606, 16),
24114 => conv_std_logic_vector(4700, 16),
24115 => conv_std_logic_vector(4794, 16),
24116 => conv_std_logic_vector(4888, 16),
24117 => conv_std_logic_vector(4982, 16),
24118 => conv_std_logic_vector(5076, 16),
24119 => conv_std_logic_vector(5170, 16),
24120 => conv_std_logic_vector(5264, 16),
24121 => conv_std_logic_vector(5358, 16),
24122 => conv_std_logic_vector(5452, 16),
24123 => conv_std_logic_vector(5546, 16),
24124 => conv_std_logic_vector(5640, 16),
24125 => conv_std_logic_vector(5734, 16),
24126 => conv_std_logic_vector(5828, 16),
24127 => conv_std_logic_vector(5922, 16),
24128 => conv_std_logic_vector(6016, 16),
24129 => conv_std_logic_vector(6110, 16),
24130 => conv_std_logic_vector(6204, 16),
24131 => conv_std_logic_vector(6298, 16),
24132 => conv_std_logic_vector(6392, 16),
24133 => conv_std_logic_vector(6486, 16),
24134 => conv_std_logic_vector(6580, 16),
24135 => conv_std_logic_vector(6674, 16),
24136 => conv_std_logic_vector(6768, 16),
24137 => conv_std_logic_vector(6862, 16),
24138 => conv_std_logic_vector(6956, 16),
24139 => conv_std_logic_vector(7050, 16),
24140 => conv_std_logic_vector(7144, 16),
24141 => conv_std_logic_vector(7238, 16),
24142 => conv_std_logic_vector(7332, 16),
24143 => conv_std_logic_vector(7426, 16),
24144 => conv_std_logic_vector(7520, 16),
24145 => conv_std_logic_vector(7614, 16),
24146 => conv_std_logic_vector(7708, 16),
24147 => conv_std_logic_vector(7802, 16),
24148 => conv_std_logic_vector(7896, 16),
24149 => conv_std_logic_vector(7990, 16),
24150 => conv_std_logic_vector(8084, 16),
24151 => conv_std_logic_vector(8178, 16),
24152 => conv_std_logic_vector(8272, 16),
24153 => conv_std_logic_vector(8366, 16),
24154 => conv_std_logic_vector(8460, 16),
24155 => conv_std_logic_vector(8554, 16),
24156 => conv_std_logic_vector(8648, 16),
24157 => conv_std_logic_vector(8742, 16),
24158 => conv_std_logic_vector(8836, 16),
24159 => conv_std_logic_vector(8930, 16),
24160 => conv_std_logic_vector(9024, 16),
24161 => conv_std_logic_vector(9118, 16),
24162 => conv_std_logic_vector(9212, 16),
24163 => conv_std_logic_vector(9306, 16),
24164 => conv_std_logic_vector(9400, 16),
24165 => conv_std_logic_vector(9494, 16),
24166 => conv_std_logic_vector(9588, 16),
24167 => conv_std_logic_vector(9682, 16),
24168 => conv_std_logic_vector(9776, 16),
24169 => conv_std_logic_vector(9870, 16),
24170 => conv_std_logic_vector(9964, 16),
24171 => conv_std_logic_vector(10058, 16),
24172 => conv_std_logic_vector(10152, 16),
24173 => conv_std_logic_vector(10246, 16),
24174 => conv_std_logic_vector(10340, 16),
24175 => conv_std_logic_vector(10434, 16),
24176 => conv_std_logic_vector(10528, 16),
24177 => conv_std_logic_vector(10622, 16),
24178 => conv_std_logic_vector(10716, 16),
24179 => conv_std_logic_vector(10810, 16),
24180 => conv_std_logic_vector(10904, 16),
24181 => conv_std_logic_vector(10998, 16),
24182 => conv_std_logic_vector(11092, 16),
24183 => conv_std_logic_vector(11186, 16),
24184 => conv_std_logic_vector(11280, 16),
24185 => conv_std_logic_vector(11374, 16),
24186 => conv_std_logic_vector(11468, 16),
24187 => conv_std_logic_vector(11562, 16),
24188 => conv_std_logic_vector(11656, 16),
24189 => conv_std_logic_vector(11750, 16),
24190 => conv_std_logic_vector(11844, 16),
24191 => conv_std_logic_vector(11938, 16),
24192 => conv_std_logic_vector(12032, 16),
24193 => conv_std_logic_vector(12126, 16),
24194 => conv_std_logic_vector(12220, 16),
24195 => conv_std_logic_vector(12314, 16),
24196 => conv_std_logic_vector(12408, 16),
24197 => conv_std_logic_vector(12502, 16),
24198 => conv_std_logic_vector(12596, 16),
24199 => conv_std_logic_vector(12690, 16),
24200 => conv_std_logic_vector(12784, 16),
24201 => conv_std_logic_vector(12878, 16),
24202 => conv_std_logic_vector(12972, 16),
24203 => conv_std_logic_vector(13066, 16),
24204 => conv_std_logic_vector(13160, 16),
24205 => conv_std_logic_vector(13254, 16),
24206 => conv_std_logic_vector(13348, 16),
24207 => conv_std_logic_vector(13442, 16),
24208 => conv_std_logic_vector(13536, 16),
24209 => conv_std_logic_vector(13630, 16),
24210 => conv_std_logic_vector(13724, 16),
24211 => conv_std_logic_vector(13818, 16),
24212 => conv_std_logic_vector(13912, 16),
24213 => conv_std_logic_vector(14006, 16),
24214 => conv_std_logic_vector(14100, 16),
24215 => conv_std_logic_vector(14194, 16),
24216 => conv_std_logic_vector(14288, 16),
24217 => conv_std_logic_vector(14382, 16),
24218 => conv_std_logic_vector(14476, 16),
24219 => conv_std_logic_vector(14570, 16),
24220 => conv_std_logic_vector(14664, 16),
24221 => conv_std_logic_vector(14758, 16),
24222 => conv_std_logic_vector(14852, 16),
24223 => conv_std_logic_vector(14946, 16),
24224 => conv_std_logic_vector(15040, 16),
24225 => conv_std_logic_vector(15134, 16),
24226 => conv_std_logic_vector(15228, 16),
24227 => conv_std_logic_vector(15322, 16),
24228 => conv_std_logic_vector(15416, 16),
24229 => conv_std_logic_vector(15510, 16),
24230 => conv_std_logic_vector(15604, 16),
24231 => conv_std_logic_vector(15698, 16),
24232 => conv_std_logic_vector(15792, 16),
24233 => conv_std_logic_vector(15886, 16),
24234 => conv_std_logic_vector(15980, 16),
24235 => conv_std_logic_vector(16074, 16),
24236 => conv_std_logic_vector(16168, 16),
24237 => conv_std_logic_vector(16262, 16),
24238 => conv_std_logic_vector(16356, 16),
24239 => conv_std_logic_vector(16450, 16),
24240 => conv_std_logic_vector(16544, 16),
24241 => conv_std_logic_vector(16638, 16),
24242 => conv_std_logic_vector(16732, 16),
24243 => conv_std_logic_vector(16826, 16),
24244 => conv_std_logic_vector(16920, 16),
24245 => conv_std_logic_vector(17014, 16),
24246 => conv_std_logic_vector(17108, 16),
24247 => conv_std_logic_vector(17202, 16),
24248 => conv_std_logic_vector(17296, 16),
24249 => conv_std_logic_vector(17390, 16),
24250 => conv_std_logic_vector(17484, 16),
24251 => conv_std_logic_vector(17578, 16),
24252 => conv_std_logic_vector(17672, 16),
24253 => conv_std_logic_vector(17766, 16),
24254 => conv_std_logic_vector(17860, 16),
24255 => conv_std_logic_vector(17954, 16),
24256 => conv_std_logic_vector(18048, 16),
24257 => conv_std_logic_vector(18142, 16),
24258 => conv_std_logic_vector(18236, 16),
24259 => conv_std_logic_vector(18330, 16),
24260 => conv_std_logic_vector(18424, 16),
24261 => conv_std_logic_vector(18518, 16),
24262 => conv_std_logic_vector(18612, 16),
24263 => conv_std_logic_vector(18706, 16),
24264 => conv_std_logic_vector(18800, 16),
24265 => conv_std_logic_vector(18894, 16),
24266 => conv_std_logic_vector(18988, 16),
24267 => conv_std_logic_vector(19082, 16),
24268 => conv_std_logic_vector(19176, 16),
24269 => conv_std_logic_vector(19270, 16),
24270 => conv_std_logic_vector(19364, 16),
24271 => conv_std_logic_vector(19458, 16),
24272 => conv_std_logic_vector(19552, 16),
24273 => conv_std_logic_vector(19646, 16),
24274 => conv_std_logic_vector(19740, 16),
24275 => conv_std_logic_vector(19834, 16),
24276 => conv_std_logic_vector(19928, 16),
24277 => conv_std_logic_vector(20022, 16),
24278 => conv_std_logic_vector(20116, 16),
24279 => conv_std_logic_vector(20210, 16),
24280 => conv_std_logic_vector(20304, 16),
24281 => conv_std_logic_vector(20398, 16),
24282 => conv_std_logic_vector(20492, 16),
24283 => conv_std_logic_vector(20586, 16),
24284 => conv_std_logic_vector(20680, 16),
24285 => conv_std_logic_vector(20774, 16),
24286 => conv_std_logic_vector(20868, 16),
24287 => conv_std_logic_vector(20962, 16),
24288 => conv_std_logic_vector(21056, 16),
24289 => conv_std_logic_vector(21150, 16),
24290 => conv_std_logic_vector(21244, 16),
24291 => conv_std_logic_vector(21338, 16),
24292 => conv_std_logic_vector(21432, 16),
24293 => conv_std_logic_vector(21526, 16),
24294 => conv_std_logic_vector(21620, 16),
24295 => conv_std_logic_vector(21714, 16),
24296 => conv_std_logic_vector(21808, 16),
24297 => conv_std_logic_vector(21902, 16),
24298 => conv_std_logic_vector(21996, 16),
24299 => conv_std_logic_vector(22090, 16),
24300 => conv_std_logic_vector(22184, 16),
24301 => conv_std_logic_vector(22278, 16),
24302 => conv_std_logic_vector(22372, 16),
24303 => conv_std_logic_vector(22466, 16),
24304 => conv_std_logic_vector(22560, 16),
24305 => conv_std_logic_vector(22654, 16),
24306 => conv_std_logic_vector(22748, 16),
24307 => conv_std_logic_vector(22842, 16),
24308 => conv_std_logic_vector(22936, 16),
24309 => conv_std_logic_vector(23030, 16),
24310 => conv_std_logic_vector(23124, 16),
24311 => conv_std_logic_vector(23218, 16),
24312 => conv_std_logic_vector(23312, 16),
24313 => conv_std_logic_vector(23406, 16),
24314 => conv_std_logic_vector(23500, 16),
24315 => conv_std_logic_vector(23594, 16),
24316 => conv_std_logic_vector(23688, 16),
24317 => conv_std_logic_vector(23782, 16),
24318 => conv_std_logic_vector(23876, 16),
24319 => conv_std_logic_vector(23970, 16),
24320 => conv_std_logic_vector(0, 16),
24321 => conv_std_logic_vector(95, 16),
24322 => conv_std_logic_vector(190, 16),
24323 => conv_std_logic_vector(285, 16),
24324 => conv_std_logic_vector(380, 16),
24325 => conv_std_logic_vector(475, 16),
24326 => conv_std_logic_vector(570, 16),
24327 => conv_std_logic_vector(665, 16),
24328 => conv_std_logic_vector(760, 16),
24329 => conv_std_logic_vector(855, 16),
24330 => conv_std_logic_vector(950, 16),
24331 => conv_std_logic_vector(1045, 16),
24332 => conv_std_logic_vector(1140, 16),
24333 => conv_std_logic_vector(1235, 16),
24334 => conv_std_logic_vector(1330, 16),
24335 => conv_std_logic_vector(1425, 16),
24336 => conv_std_logic_vector(1520, 16),
24337 => conv_std_logic_vector(1615, 16),
24338 => conv_std_logic_vector(1710, 16),
24339 => conv_std_logic_vector(1805, 16),
24340 => conv_std_logic_vector(1900, 16),
24341 => conv_std_logic_vector(1995, 16),
24342 => conv_std_logic_vector(2090, 16),
24343 => conv_std_logic_vector(2185, 16),
24344 => conv_std_logic_vector(2280, 16),
24345 => conv_std_logic_vector(2375, 16),
24346 => conv_std_logic_vector(2470, 16),
24347 => conv_std_logic_vector(2565, 16),
24348 => conv_std_logic_vector(2660, 16),
24349 => conv_std_logic_vector(2755, 16),
24350 => conv_std_logic_vector(2850, 16),
24351 => conv_std_logic_vector(2945, 16),
24352 => conv_std_logic_vector(3040, 16),
24353 => conv_std_logic_vector(3135, 16),
24354 => conv_std_logic_vector(3230, 16),
24355 => conv_std_logic_vector(3325, 16),
24356 => conv_std_logic_vector(3420, 16),
24357 => conv_std_logic_vector(3515, 16),
24358 => conv_std_logic_vector(3610, 16),
24359 => conv_std_logic_vector(3705, 16),
24360 => conv_std_logic_vector(3800, 16),
24361 => conv_std_logic_vector(3895, 16),
24362 => conv_std_logic_vector(3990, 16),
24363 => conv_std_logic_vector(4085, 16),
24364 => conv_std_logic_vector(4180, 16),
24365 => conv_std_logic_vector(4275, 16),
24366 => conv_std_logic_vector(4370, 16),
24367 => conv_std_logic_vector(4465, 16),
24368 => conv_std_logic_vector(4560, 16),
24369 => conv_std_logic_vector(4655, 16),
24370 => conv_std_logic_vector(4750, 16),
24371 => conv_std_logic_vector(4845, 16),
24372 => conv_std_logic_vector(4940, 16),
24373 => conv_std_logic_vector(5035, 16),
24374 => conv_std_logic_vector(5130, 16),
24375 => conv_std_logic_vector(5225, 16),
24376 => conv_std_logic_vector(5320, 16),
24377 => conv_std_logic_vector(5415, 16),
24378 => conv_std_logic_vector(5510, 16),
24379 => conv_std_logic_vector(5605, 16),
24380 => conv_std_logic_vector(5700, 16),
24381 => conv_std_logic_vector(5795, 16),
24382 => conv_std_logic_vector(5890, 16),
24383 => conv_std_logic_vector(5985, 16),
24384 => conv_std_logic_vector(6080, 16),
24385 => conv_std_logic_vector(6175, 16),
24386 => conv_std_logic_vector(6270, 16),
24387 => conv_std_logic_vector(6365, 16),
24388 => conv_std_logic_vector(6460, 16),
24389 => conv_std_logic_vector(6555, 16),
24390 => conv_std_logic_vector(6650, 16),
24391 => conv_std_logic_vector(6745, 16),
24392 => conv_std_logic_vector(6840, 16),
24393 => conv_std_logic_vector(6935, 16),
24394 => conv_std_logic_vector(7030, 16),
24395 => conv_std_logic_vector(7125, 16),
24396 => conv_std_logic_vector(7220, 16),
24397 => conv_std_logic_vector(7315, 16),
24398 => conv_std_logic_vector(7410, 16),
24399 => conv_std_logic_vector(7505, 16),
24400 => conv_std_logic_vector(7600, 16),
24401 => conv_std_logic_vector(7695, 16),
24402 => conv_std_logic_vector(7790, 16),
24403 => conv_std_logic_vector(7885, 16),
24404 => conv_std_logic_vector(7980, 16),
24405 => conv_std_logic_vector(8075, 16),
24406 => conv_std_logic_vector(8170, 16),
24407 => conv_std_logic_vector(8265, 16),
24408 => conv_std_logic_vector(8360, 16),
24409 => conv_std_logic_vector(8455, 16),
24410 => conv_std_logic_vector(8550, 16),
24411 => conv_std_logic_vector(8645, 16),
24412 => conv_std_logic_vector(8740, 16),
24413 => conv_std_logic_vector(8835, 16),
24414 => conv_std_logic_vector(8930, 16),
24415 => conv_std_logic_vector(9025, 16),
24416 => conv_std_logic_vector(9120, 16),
24417 => conv_std_logic_vector(9215, 16),
24418 => conv_std_logic_vector(9310, 16),
24419 => conv_std_logic_vector(9405, 16),
24420 => conv_std_logic_vector(9500, 16),
24421 => conv_std_logic_vector(9595, 16),
24422 => conv_std_logic_vector(9690, 16),
24423 => conv_std_logic_vector(9785, 16),
24424 => conv_std_logic_vector(9880, 16),
24425 => conv_std_logic_vector(9975, 16),
24426 => conv_std_logic_vector(10070, 16),
24427 => conv_std_logic_vector(10165, 16),
24428 => conv_std_logic_vector(10260, 16),
24429 => conv_std_logic_vector(10355, 16),
24430 => conv_std_logic_vector(10450, 16),
24431 => conv_std_logic_vector(10545, 16),
24432 => conv_std_logic_vector(10640, 16),
24433 => conv_std_logic_vector(10735, 16),
24434 => conv_std_logic_vector(10830, 16),
24435 => conv_std_logic_vector(10925, 16),
24436 => conv_std_logic_vector(11020, 16),
24437 => conv_std_logic_vector(11115, 16),
24438 => conv_std_logic_vector(11210, 16),
24439 => conv_std_logic_vector(11305, 16),
24440 => conv_std_logic_vector(11400, 16),
24441 => conv_std_logic_vector(11495, 16),
24442 => conv_std_logic_vector(11590, 16),
24443 => conv_std_logic_vector(11685, 16),
24444 => conv_std_logic_vector(11780, 16),
24445 => conv_std_logic_vector(11875, 16),
24446 => conv_std_logic_vector(11970, 16),
24447 => conv_std_logic_vector(12065, 16),
24448 => conv_std_logic_vector(12160, 16),
24449 => conv_std_logic_vector(12255, 16),
24450 => conv_std_logic_vector(12350, 16),
24451 => conv_std_logic_vector(12445, 16),
24452 => conv_std_logic_vector(12540, 16),
24453 => conv_std_logic_vector(12635, 16),
24454 => conv_std_logic_vector(12730, 16),
24455 => conv_std_logic_vector(12825, 16),
24456 => conv_std_logic_vector(12920, 16),
24457 => conv_std_logic_vector(13015, 16),
24458 => conv_std_logic_vector(13110, 16),
24459 => conv_std_logic_vector(13205, 16),
24460 => conv_std_logic_vector(13300, 16),
24461 => conv_std_logic_vector(13395, 16),
24462 => conv_std_logic_vector(13490, 16),
24463 => conv_std_logic_vector(13585, 16),
24464 => conv_std_logic_vector(13680, 16),
24465 => conv_std_logic_vector(13775, 16),
24466 => conv_std_logic_vector(13870, 16),
24467 => conv_std_logic_vector(13965, 16),
24468 => conv_std_logic_vector(14060, 16),
24469 => conv_std_logic_vector(14155, 16),
24470 => conv_std_logic_vector(14250, 16),
24471 => conv_std_logic_vector(14345, 16),
24472 => conv_std_logic_vector(14440, 16),
24473 => conv_std_logic_vector(14535, 16),
24474 => conv_std_logic_vector(14630, 16),
24475 => conv_std_logic_vector(14725, 16),
24476 => conv_std_logic_vector(14820, 16),
24477 => conv_std_logic_vector(14915, 16),
24478 => conv_std_logic_vector(15010, 16),
24479 => conv_std_logic_vector(15105, 16),
24480 => conv_std_logic_vector(15200, 16),
24481 => conv_std_logic_vector(15295, 16),
24482 => conv_std_logic_vector(15390, 16),
24483 => conv_std_logic_vector(15485, 16),
24484 => conv_std_logic_vector(15580, 16),
24485 => conv_std_logic_vector(15675, 16),
24486 => conv_std_logic_vector(15770, 16),
24487 => conv_std_logic_vector(15865, 16),
24488 => conv_std_logic_vector(15960, 16),
24489 => conv_std_logic_vector(16055, 16),
24490 => conv_std_logic_vector(16150, 16),
24491 => conv_std_logic_vector(16245, 16),
24492 => conv_std_logic_vector(16340, 16),
24493 => conv_std_logic_vector(16435, 16),
24494 => conv_std_logic_vector(16530, 16),
24495 => conv_std_logic_vector(16625, 16),
24496 => conv_std_logic_vector(16720, 16),
24497 => conv_std_logic_vector(16815, 16),
24498 => conv_std_logic_vector(16910, 16),
24499 => conv_std_logic_vector(17005, 16),
24500 => conv_std_logic_vector(17100, 16),
24501 => conv_std_logic_vector(17195, 16),
24502 => conv_std_logic_vector(17290, 16),
24503 => conv_std_logic_vector(17385, 16),
24504 => conv_std_logic_vector(17480, 16),
24505 => conv_std_logic_vector(17575, 16),
24506 => conv_std_logic_vector(17670, 16),
24507 => conv_std_logic_vector(17765, 16),
24508 => conv_std_logic_vector(17860, 16),
24509 => conv_std_logic_vector(17955, 16),
24510 => conv_std_logic_vector(18050, 16),
24511 => conv_std_logic_vector(18145, 16),
24512 => conv_std_logic_vector(18240, 16),
24513 => conv_std_logic_vector(18335, 16),
24514 => conv_std_logic_vector(18430, 16),
24515 => conv_std_logic_vector(18525, 16),
24516 => conv_std_logic_vector(18620, 16),
24517 => conv_std_logic_vector(18715, 16),
24518 => conv_std_logic_vector(18810, 16),
24519 => conv_std_logic_vector(18905, 16),
24520 => conv_std_logic_vector(19000, 16),
24521 => conv_std_logic_vector(19095, 16),
24522 => conv_std_logic_vector(19190, 16),
24523 => conv_std_logic_vector(19285, 16),
24524 => conv_std_logic_vector(19380, 16),
24525 => conv_std_logic_vector(19475, 16),
24526 => conv_std_logic_vector(19570, 16),
24527 => conv_std_logic_vector(19665, 16),
24528 => conv_std_logic_vector(19760, 16),
24529 => conv_std_logic_vector(19855, 16),
24530 => conv_std_logic_vector(19950, 16),
24531 => conv_std_logic_vector(20045, 16),
24532 => conv_std_logic_vector(20140, 16),
24533 => conv_std_logic_vector(20235, 16),
24534 => conv_std_logic_vector(20330, 16),
24535 => conv_std_logic_vector(20425, 16),
24536 => conv_std_logic_vector(20520, 16),
24537 => conv_std_logic_vector(20615, 16),
24538 => conv_std_logic_vector(20710, 16),
24539 => conv_std_logic_vector(20805, 16),
24540 => conv_std_logic_vector(20900, 16),
24541 => conv_std_logic_vector(20995, 16),
24542 => conv_std_logic_vector(21090, 16),
24543 => conv_std_logic_vector(21185, 16),
24544 => conv_std_logic_vector(21280, 16),
24545 => conv_std_logic_vector(21375, 16),
24546 => conv_std_logic_vector(21470, 16),
24547 => conv_std_logic_vector(21565, 16),
24548 => conv_std_logic_vector(21660, 16),
24549 => conv_std_logic_vector(21755, 16),
24550 => conv_std_logic_vector(21850, 16),
24551 => conv_std_logic_vector(21945, 16),
24552 => conv_std_logic_vector(22040, 16),
24553 => conv_std_logic_vector(22135, 16),
24554 => conv_std_logic_vector(22230, 16),
24555 => conv_std_logic_vector(22325, 16),
24556 => conv_std_logic_vector(22420, 16),
24557 => conv_std_logic_vector(22515, 16),
24558 => conv_std_logic_vector(22610, 16),
24559 => conv_std_logic_vector(22705, 16),
24560 => conv_std_logic_vector(22800, 16),
24561 => conv_std_logic_vector(22895, 16),
24562 => conv_std_logic_vector(22990, 16),
24563 => conv_std_logic_vector(23085, 16),
24564 => conv_std_logic_vector(23180, 16),
24565 => conv_std_logic_vector(23275, 16),
24566 => conv_std_logic_vector(23370, 16),
24567 => conv_std_logic_vector(23465, 16),
24568 => conv_std_logic_vector(23560, 16),
24569 => conv_std_logic_vector(23655, 16),
24570 => conv_std_logic_vector(23750, 16),
24571 => conv_std_logic_vector(23845, 16),
24572 => conv_std_logic_vector(23940, 16),
24573 => conv_std_logic_vector(24035, 16),
24574 => conv_std_logic_vector(24130, 16),
24575 => conv_std_logic_vector(24225, 16),
24576 => conv_std_logic_vector(0, 16),
24577 => conv_std_logic_vector(96, 16),
24578 => conv_std_logic_vector(192, 16),
24579 => conv_std_logic_vector(288, 16),
24580 => conv_std_logic_vector(384, 16),
24581 => conv_std_logic_vector(480, 16),
24582 => conv_std_logic_vector(576, 16),
24583 => conv_std_logic_vector(672, 16),
24584 => conv_std_logic_vector(768, 16),
24585 => conv_std_logic_vector(864, 16),
24586 => conv_std_logic_vector(960, 16),
24587 => conv_std_logic_vector(1056, 16),
24588 => conv_std_logic_vector(1152, 16),
24589 => conv_std_logic_vector(1248, 16),
24590 => conv_std_logic_vector(1344, 16),
24591 => conv_std_logic_vector(1440, 16),
24592 => conv_std_logic_vector(1536, 16),
24593 => conv_std_logic_vector(1632, 16),
24594 => conv_std_logic_vector(1728, 16),
24595 => conv_std_logic_vector(1824, 16),
24596 => conv_std_logic_vector(1920, 16),
24597 => conv_std_logic_vector(2016, 16),
24598 => conv_std_logic_vector(2112, 16),
24599 => conv_std_logic_vector(2208, 16),
24600 => conv_std_logic_vector(2304, 16),
24601 => conv_std_logic_vector(2400, 16),
24602 => conv_std_logic_vector(2496, 16),
24603 => conv_std_logic_vector(2592, 16),
24604 => conv_std_logic_vector(2688, 16),
24605 => conv_std_logic_vector(2784, 16),
24606 => conv_std_logic_vector(2880, 16),
24607 => conv_std_logic_vector(2976, 16),
24608 => conv_std_logic_vector(3072, 16),
24609 => conv_std_logic_vector(3168, 16),
24610 => conv_std_logic_vector(3264, 16),
24611 => conv_std_logic_vector(3360, 16),
24612 => conv_std_logic_vector(3456, 16),
24613 => conv_std_logic_vector(3552, 16),
24614 => conv_std_logic_vector(3648, 16),
24615 => conv_std_logic_vector(3744, 16),
24616 => conv_std_logic_vector(3840, 16),
24617 => conv_std_logic_vector(3936, 16),
24618 => conv_std_logic_vector(4032, 16),
24619 => conv_std_logic_vector(4128, 16),
24620 => conv_std_logic_vector(4224, 16),
24621 => conv_std_logic_vector(4320, 16),
24622 => conv_std_logic_vector(4416, 16),
24623 => conv_std_logic_vector(4512, 16),
24624 => conv_std_logic_vector(4608, 16),
24625 => conv_std_logic_vector(4704, 16),
24626 => conv_std_logic_vector(4800, 16),
24627 => conv_std_logic_vector(4896, 16),
24628 => conv_std_logic_vector(4992, 16),
24629 => conv_std_logic_vector(5088, 16),
24630 => conv_std_logic_vector(5184, 16),
24631 => conv_std_logic_vector(5280, 16),
24632 => conv_std_logic_vector(5376, 16),
24633 => conv_std_logic_vector(5472, 16),
24634 => conv_std_logic_vector(5568, 16),
24635 => conv_std_logic_vector(5664, 16),
24636 => conv_std_logic_vector(5760, 16),
24637 => conv_std_logic_vector(5856, 16),
24638 => conv_std_logic_vector(5952, 16),
24639 => conv_std_logic_vector(6048, 16),
24640 => conv_std_logic_vector(6144, 16),
24641 => conv_std_logic_vector(6240, 16),
24642 => conv_std_logic_vector(6336, 16),
24643 => conv_std_logic_vector(6432, 16),
24644 => conv_std_logic_vector(6528, 16),
24645 => conv_std_logic_vector(6624, 16),
24646 => conv_std_logic_vector(6720, 16),
24647 => conv_std_logic_vector(6816, 16),
24648 => conv_std_logic_vector(6912, 16),
24649 => conv_std_logic_vector(7008, 16),
24650 => conv_std_logic_vector(7104, 16),
24651 => conv_std_logic_vector(7200, 16),
24652 => conv_std_logic_vector(7296, 16),
24653 => conv_std_logic_vector(7392, 16),
24654 => conv_std_logic_vector(7488, 16),
24655 => conv_std_logic_vector(7584, 16),
24656 => conv_std_logic_vector(7680, 16),
24657 => conv_std_logic_vector(7776, 16),
24658 => conv_std_logic_vector(7872, 16),
24659 => conv_std_logic_vector(7968, 16),
24660 => conv_std_logic_vector(8064, 16),
24661 => conv_std_logic_vector(8160, 16),
24662 => conv_std_logic_vector(8256, 16),
24663 => conv_std_logic_vector(8352, 16),
24664 => conv_std_logic_vector(8448, 16),
24665 => conv_std_logic_vector(8544, 16),
24666 => conv_std_logic_vector(8640, 16),
24667 => conv_std_logic_vector(8736, 16),
24668 => conv_std_logic_vector(8832, 16),
24669 => conv_std_logic_vector(8928, 16),
24670 => conv_std_logic_vector(9024, 16),
24671 => conv_std_logic_vector(9120, 16),
24672 => conv_std_logic_vector(9216, 16),
24673 => conv_std_logic_vector(9312, 16),
24674 => conv_std_logic_vector(9408, 16),
24675 => conv_std_logic_vector(9504, 16),
24676 => conv_std_logic_vector(9600, 16),
24677 => conv_std_logic_vector(9696, 16),
24678 => conv_std_logic_vector(9792, 16),
24679 => conv_std_logic_vector(9888, 16),
24680 => conv_std_logic_vector(9984, 16),
24681 => conv_std_logic_vector(10080, 16),
24682 => conv_std_logic_vector(10176, 16),
24683 => conv_std_logic_vector(10272, 16),
24684 => conv_std_logic_vector(10368, 16),
24685 => conv_std_logic_vector(10464, 16),
24686 => conv_std_logic_vector(10560, 16),
24687 => conv_std_logic_vector(10656, 16),
24688 => conv_std_logic_vector(10752, 16),
24689 => conv_std_logic_vector(10848, 16),
24690 => conv_std_logic_vector(10944, 16),
24691 => conv_std_logic_vector(11040, 16),
24692 => conv_std_logic_vector(11136, 16),
24693 => conv_std_logic_vector(11232, 16),
24694 => conv_std_logic_vector(11328, 16),
24695 => conv_std_logic_vector(11424, 16),
24696 => conv_std_logic_vector(11520, 16),
24697 => conv_std_logic_vector(11616, 16),
24698 => conv_std_logic_vector(11712, 16),
24699 => conv_std_logic_vector(11808, 16),
24700 => conv_std_logic_vector(11904, 16),
24701 => conv_std_logic_vector(12000, 16),
24702 => conv_std_logic_vector(12096, 16),
24703 => conv_std_logic_vector(12192, 16),
24704 => conv_std_logic_vector(12288, 16),
24705 => conv_std_logic_vector(12384, 16),
24706 => conv_std_logic_vector(12480, 16),
24707 => conv_std_logic_vector(12576, 16),
24708 => conv_std_logic_vector(12672, 16),
24709 => conv_std_logic_vector(12768, 16),
24710 => conv_std_logic_vector(12864, 16),
24711 => conv_std_logic_vector(12960, 16),
24712 => conv_std_logic_vector(13056, 16),
24713 => conv_std_logic_vector(13152, 16),
24714 => conv_std_logic_vector(13248, 16),
24715 => conv_std_logic_vector(13344, 16),
24716 => conv_std_logic_vector(13440, 16),
24717 => conv_std_logic_vector(13536, 16),
24718 => conv_std_logic_vector(13632, 16),
24719 => conv_std_logic_vector(13728, 16),
24720 => conv_std_logic_vector(13824, 16),
24721 => conv_std_logic_vector(13920, 16),
24722 => conv_std_logic_vector(14016, 16),
24723 => conv_std_logic_vector(14112, 16),
24724 => conv_std_logic_vector(14208, 16),
24725 => conv_std_logic_vector(14304, 16),
24726 => conv_std_logic_vector(14400, 16),
24727 => conv_std_logic_vector(14496, 16),
24728 => conv_std_logic_vector(14592, 16),
24729 => conv_std_logic_vector(14688, 16),
24730 => conv_std_logic_vector(14784, 16),
24731 => conv_std_logic_vector(14880, 16),
24732 => conv_std_logic_vector(14976, 16),
24733 => conv_std_logic_vector(15072, 16),
24734 => conv_std_logic_vector(15168, 16),
24735 => conv_std_logic_vector(15264, 16),
24736 => conv_std_logic_vector(15360, 16),
24737 => conv_std_logic_vector(15456, 16),
24738 => conv_std_logic_vector(15552, 16),
24739 => conv_std_logic_vector(15648, 16),
24740 => conv_std_logic_vector(15744, 16),
24741 => conv_std_logic_vector(15840, 16),
24742 => conv_std_logic_vector(15936, 16),
24743 => conv_std_logic_vector(16032, 16),
24744 => conv_std_logic_vector(16128, 16),
24745 => conv_std_logic_vector(16224, 16),
24746 => conv_std_logic_vector(16320, 16),
24747 => conv_std_logic_vector(16416, 16),
24748 => conv_std_logic_vector(16512, 16),
24749 => conv_std_logic_vector(16608, 16),
24750 => conv_std_logic_vector(16704, 16),
24751 => conv_std_logic_vector(16800, 16),
24752 => conv_std_logic_vector(16896, 16),
24753 => conv_std_logic_vector(16992, 16),
24754 => conv_std_logic_vector(17088, 16),
24755 => conv_std_logic_vector(17184, 16),
24756 => conv_std_logic_vector(17280, 16),
24757 => conv_std_logic_vector(17376, 16),
24758 => conv_std_logic_vector(17472, 16),
24759 => conv_std_logic_vector(17568, 16),
24760 => conv_std_logic_vector(17664, 16),
24761 => conv_std_logic_vector(17760, 16),
24762 => conv_std_logic_vector(17856, 16),
24763 => conv_std_logic_vector(17952, 16),
24764 => conv_std_logic_vector(18048, 16),
24765 => conv_std_logic_vector(18144, 16),
24766 => conv_std_logic_vector(18240, 16),
24767 => conv_std_logic_vector(18336, 16),
24768 => conv_std_logic_vector(18432, 16),
24769 => conv_std_logic_vector(18528, 16),
24770 => conv_std_logic_vector(18624, 16),
24771 => conv_std_logic_vector(18720, 16),
24772 => conv_std_logic_vector(18816, 16),
24773 => conv_std_logic_vector(18912, 16),
24774 => conv_std_logic_vector(19008, 16),
24775 => conv_std_logic_vector(19104, 16),
24776 => conv_std_logic_vector(19200, 16),
24777 => conv_std_logic_vector(19296, 16),
24778 => conv_std_logic_vector(19392, 16),
24779 => conv_std_logic_vector(19488, 16),
24780 => conv_std_logic_vector(19584, 16),
24781 => conv_std_logic_vector(19680, 16),
24782 => conv_std_logic_vector(19776, 16),
24783 => conv_std_logic_vector(19872, 16),
24784 => conv_std_logic_vector(19968, 16),
24785 => conv_std_logic_vector(20064, 16),
24786 => conv_std_logic_vector(20160, 16),
24787 => conv_std_logic_vector(20256, 16),
24788 => conv_std_logic_vector(20352, 16),
24789 => conv_std_logic_vector(20448, 16),
24790 => conv_std_logic_vector(20544, 16),
24791 => conv_std_logic_vector(20640, 16),
24792 => conv_std_logic_vector(20736, 16),
24793 => conv_std_logic_vector(20832, 16),
24794 => conv_std_logic_vector(20928, 16),
24795 => conv_std_logic_vector(21024, 16),
24796 => conv_std_logic_vector(21120, 16),
24797 => conv_std_logic_vector(21216, 16),
24798 => conv_std_logic_vector(21312, 16),
24799 => conv_std_logic_vector(21408, 16),
24800 => conv_std_logic_vector(21504, 16),
24801 => conv_std_logic_vector(21600, 16),
24802 => conv_std_logic_vector(21696, 16),
24803 => conv_std_logic_vector(21792, 16),
24804 => conv_std_logic_vector(21888, 16),
24805 => conv_std_logic_vector(21984, 16),
24806 => conv_std_logic_vector(22080, 16),
24807 => conv_std_logic_vector(22176, 16),
24808 => conv_std_logic_vector(22272, 16),
24809 => conv_std_logic_vector(22368, 16),
24810 => conv_std_logic_vector(22464, 16),
24811 => conv_std_logic_vector(22560, 16),
24812 => conv_std_logic_vector(22656, 16),
24813 => conv_std_logic_vector(22752, 16),
24814 => conv_std_logic_vector(22848, 16),
24815 => conv_std_logic_vector(22944, 16),
24816 => conv_std_logic_vector(23040, 16),
24817 => conv_std_logic_vector(23136, 16),
24818 => conv_std_logic_vector(23232, 16),
24819 => conv_std_logic_vector(23328, 16),
24820 => conv_std_logic_vector(23424, 16),
24821 => conv_std_logic_vector(23520, 16),
24822 => conv_std_logic_vector(23616, 16),
24823 => conv_std_logic_vector(23712, 16),
24824 => conv_std_logic_vector(23808, 16),
24825 => conv_std_logic_vector(23904, 16),
24826 => conv_std_logic_vector(24000, 16),
24827 => conv_std_logic_vector(24096, 16),
24828 => conv_std_logic_vector(24192, 16),
24829 => conv_std_logic_vector(24288, 16),
24830 => conv_std_logic_vector(24384, 16),
24831 => conv_std_logic_vector(24480, 16),
24832 => conv_std_logic_vector(0, 16),
24833 => conv_std_logic_vector(97, 16),
24834 => conv_std_logic_vector(194, 16),
24835 => conv_std_logic_vector(291, 16),
24836 => conv_std_logic_vector(388, 16),
24837 => conv_std_logic_vector(485, 16),
24838 => conv_std_logic_vector(582, 16),
24839 => conv_std_logic_vector(679, 16),
24840 => conv_std_logic_vector(776, 16),
24841 => conv_std_logic_vector(873, 16),
24842 => conv_std_logic_vector(970, 16),
24843 => conv_std_logic_vector(1067, 16),
24844 => conv_std_logic_vector(1164, 16),
24845 => conv_std_logic_vector(1261, 16),
24846 => conv_std_logic_vector(1358, 16),
24847 => conv_std_logic_vector(1455, 16),
24848 => conv_std_logic_vector(1552, 16),
24849 => conv_std_logic_vector(1649, 16),
24850 => conv_std_logic_vector(1746, 16),
24851 => conv_std_logic_vector(1843, 16),
24852 => conv_std_logic_vector(1940, 16),
24853 => conv_std_logic_vector(2037, 16),
24854 => conv_std_logic_vector(2134, 16),
24855 => conv_std_logic_vector(2231, 16),
24856 => conv_std_logic_vector(2328, 16),
24857 => conv_std_logic_vector(2425, 16),
24858 => conv_std_logic_vector(2522, 16),
24859 => conv_std_logic_vector(2619, 16),
24860 => conv_std_logic_vector(2716, 16),
24861 => conv_std_logic_vector(2813, 16),
24862 => conv_std_logic_vector(2910, 16),
24863 => conv_std_logic_vector(3007, 16),
24864 => conv_std_logic_vector(3104, 16),
24865 => conv_std_logic_vector(3201, 16),
24866 => conv_std_logic_vector(3298, 16),
24867 => conv_std_logic_vector(3395, 16),
24868 => conv_std_logic_vector(3492, 16),
24869 => conv_std_logic_vector(3589, 16),
24870 => conv_std_logic_vector(3686, 16),
24871 => conv_std_logic_vector(3783, 16),
24872 => conv_std_logic_vector(3880, 16),
24873 => conv_std_logic_vector(3977, 16),
24874 => conv_std_logic_vector(4074, 16),
24875 => conv_std_logic_vector(4171, 16),
24876 => conv_std_logic_vector(4268, 16),
24877 => conv_std_logic_vector(4365, 16),
24878 => conv_std_logic_vector(4462, 16),
24879 => conv_std_logic_vector(4559, 16),
24880 => conv_std_logic_vector(4656, 16),
24881 => conv_std_logic_vector(4753, 16),
24882 => conv_std_logic_vector(4850, 16),
24883 => conv_std_logic_vector(4947, 16),
24884 => conv_std_logic_vector(5044, 16),
24885 => conv_std_logic_vector(5141, 16),
24886 => conv_std_logic_vector(5238, 16),
24887 => conv_std_logic_vector(5335, 16),
24888 => conv_std_logic_vector(5432, 16),
24889 => conv_std_logic_vector(5529, 16),
24890 => conv_std_logic_vector(5626, 16),
24891 => conv_std_logic_vector(5723, 16),
24892 => conv_std_logic_vector(5820, 16),
24893 => conv_std_logic_vector(5917, 16),
24894 => conv_std_logic_vector(6014, 16),
24895 => conv_std_logic_vector(6111, 16),
24896 => conv_std_logic_vector(6208, 16),
24897 => conv_std_logic_vector(6305, 16),
24898 => conv_std_logic_vector(6402, 16),
24899 => conv_std_logic_vector(6499, 16),
24900 => conv_std_logic_vector(6596, 16),
24901 => conv_std_logic_vector(6693, 16),
24902 => conv_std_logic_vector(6790, 16),
24903 => conv_std_logic_vector(6887, 16),
24904 => conv_std_logic_vector(6984, 16),
24905 => conv_std_logic_vector(7081, 16),
24906 => conv_std_logic_vector(7178, 16),
24907 => conv_std_logic_vector(7275, 16),
24908 => conv_std_logic_vector(7372, 16),
24909 => conv_std_logic_vector(7469, 16),
24910 => conv_std_logic_vector(7566, 16),
24911 => conv_std_logic_vector(7663, 16),
24912 => conv_std_logic_vector(7760, 16),
24913 => conv_std_logic_vector(7857, 16),
24914 => conv_std_logic_vector(7954, 16),
24915 => conv_std_logic_vector(8051, 16),
24916 => conv_std_logic_vector(8148, 16),
24917 => conv_std_logic_vector(8245, 16),
24918 => conv_std_logic_vector(8342, 16),
24919 => conv_std_logic_vector(8439, 16),
24920 => conv_std_logic_vector(8536, 16),
24921 => conv_std_logic_vector(8633, 16),
24922 => conv_std_logic_vector(8730, 16),
24923 => conv_std_logic_vector(8827, 16),
24924 => conv_std_logic_vector(8924, 16),
24925 => conv_std_logic_vector(9021, 16),
24926 => conv_std_logic_vector(9118, 16),
24927 => conv_std_logic_vector(9215, 16),
24928 => conv_std_logic_vector(9312, 16),
24929 => conv_std_logic_vector(9409, 16),
24930 => conv_std_logic_vector(9506, 16),
24931 => conv_std_logic_vector(9603, 16),
24932 => conv_std_logic_vector(9700, 16),
24933 => conv_std_logic_vector(9797, 16),
24934 => conv_std_logic_vector(9894, 16),
24935 => conv_std_logic_vector(9991, 16),
24936 => conv_std_logic_vector(10088, 16),
24937 => conv_std_logic_vector(10185, 16),
24938 => conv_std_logic_vector(10282, 16),
24939 => conv_std_logic_vector(10379, 16),
24940 => conv_std_logic_vector(10476, 16),
24941 => conv_std_logic_vector(10573, 16),
24942 => conv_std_logic_vector(10670, 16),
24943 => conv_std_logic_vector(10767, 16),
24944 => conv_std_logic_vector(10864, 16),
24945 => conv_std_logic_vector(10961, 16),
24946 => conv_std_logic_vector(11058, 16),
24947 => conv_std_logic_vector(11155, 16),
24948 => conv_std_logic_vector(11252, 16),
24949 => conv_std_logic_vector(11349, 16),
24950 => conv_std_logic_vector(11446, 16),
24951 => conv_std_logic_vector(11543, 16),
24952 => conv_std_logic_vector(11640, 16),
24953 => conv_std_logic_vector(11737, 16),
24954 => conv_std_logic_vector(11834, 16),
24955 => conv_std_logic_vector(11931, 16),
24956 => conv_std_logic_vector(12028, 16),
24957 => conv_std_logic_vector(12125, 16),
24958 => conv_std_logic_vector(12222, 16),
24959 => conv_std_logic_vector(12319, 16),
24960 => conv_std_logic_vector(12416, 16),
24961 => conv_std_logic_vector(12513, 16),
24962 => conv_std_logic_vector(12610, 16),
24963 => conv_std_logic_vector(12707, 16),
24964 => conv_std_logic_vector(12804, 16),
24965 => conv_std_logic_vector(12901, 16),
24966 => conv_std_logic_vector(12998, 16),
24967 => conv_std_logic_vector(13095, 16),
24968 => conv_std_logic_vector(13192, 16),
24969 => conv_std_logic_vector(13289, 16),
24970 => conv_std_logic_vector(13386, 16),
24971 => conv_std_logic_vector(13483, 16),
24972 => conv_std_logic_vector(13580, 16),
24973 => conv_std_logic_vector(13677, 16),
24974 => conv_std_logic_vector(13774, 16),
24975 => conv_std_logic_vector(13871, 16),
24976 => conv_std_logic_vector(13968, 16),
24977 => conv_std_logic_vector(14065, 16),
24978 => conv_std_logic_vector(14162, 16),
24979 => conv_std_logic_vector(14259, 16),
24980 => conv_std_logic_vector(14356, 16),
24981 => conv_std_logic_vector(14453, 16),
24982 => conv_std_logic_vector(14550, 16),
24983 => conv_std_logic_vector(14647, 16),
24984 => conv_std_logic_vector(14744, 16),
24985 => conv_std_logic_vector(14841, 16),
24986 => conv_std_logic_vector(14938, 16),
24987 => conv_std_logic_vector(15035, 16),
24988 => conv_std_logic_vector(15132, 16),
24989 => conv_std_logic_vector(15229, 16),
24990 => conv_std_logic_vector(15326, 16),
24991 => conv_std_logic_vector(15423, 16),
24992 => conv_std_logic_vector(15520, 16),
24993 => conv_std_logic_vector(15617, 16),
24994 => conv_std_logic_vector(15714, 16),
24995 => conv_std_logic_vector(15811, 16),
24996 => conv_std_logic_vector(15908, 16),
24997 => conv_std_logic_vector(16005, 16),
24998 => conv_std_logic_vector(16102, 16),
24999 => conv_std_logic_vector(16199, 16),
25000 => conv_std_logic_vector(16296, 16),
25001 => conv_std_logic_vector(16393, 16),
25002 => conv_std_logic_vector(16490, 16),
25003 => conv_std_logic_vector(16587, 16),
25004 => conv_std_logic_vector(16684, 16),
25005 => conv_std_logic_vector(16781, 16),
25006 => conv_std_logic_vector(16878, 16),
25007 => conv_std_logic_vector(16975, 16),
25008 => conv_std_logic_vector(17072, 16),
25009 => conv_std_logic_vector(17169, 16),
25010 => conv_std_logic_vector(17266, 16),
25011 => conv_std_logic_vector(17363, 16),
25012 => conv_std_logic_vector(17460, 16),
25013 => conv_std_logic_vector(17557, 16),
25014 => conv_std_logic_vector(17654, 16),
25015 => conv_std_logic_vector(17751, 16),
25016 => conv_std_logic_vector(17848, 16),
25017 => conv_std_logic_vector(17945, 16),
25018 => conv_std_logic_vector(18042, 16),
25019 => conv_std_logic_vector(18139, 16),
25020 => conv_std_logic_vector(18236, 16),
25021 => conv_std_logic_vector(18333, 16),
25022 => conv_std_logic_vector(18430, 16),
25023 => conv_std_logic_vector(18527, 16),
25024 => conv_std_logic_vector(18624, 16),
25025 => conv_std_logic_vector(18721, 16),
25026 => conv_std_logic_vector(18818, 16),
25027 => conv_std_logic_vector(18915, 16),
25028 => conv_std_logic_vector(19012, 16),
25029 => conv_std_logic_vector(19109, 16),
25030 => conv_std_logic_vector(19206, 16),
25031 => conv_std_logic_vector(19303, 16),
25032 => conv_std_logic_vector(19400, 16),
25033 => conv_std_logic_vector(19497, 16),
25034 => conv_std_logic_vector(19594, 16),
25035 => conv_std_logic_vector(19691, 16),
25036 => conv_std_logic_vector(19788, 16),
25037 => conv_std_logic_vector(19885, 16),
25038 => conv_std_logic_vector(19982, 16),
25039 => conv_std_logic_vector(20079, 16),
25040 => conv_std_logic_vector(20176, 16),
25041 => conv_std_logic_vector(20273, 16),
25042 => conv_std_logic_vector(20370, 16),
25043 => conv_std_logic_vector(20467, 16),
25044 => conv_std_logic_vector(20564, 16),
25045 => conv_std_logic_vector(20661, 16),
25046 => conv_std_logic_vector(20758, 16),
25047 => conv_std_logic_vector(20855, 16),
25048 => conv_std_logic_vector(20952, 16),
25049 => conv_std_logic_vector(21049, 16),
25050 => conv_std_logic_vector(21146, 16),
25051 => conv_std_logic_vector(21243, 16),
25052 => conv_std_logic_vector(21340, 16),
25053 => conv_std_logic_vector(21437, 16),
25054 => conv_std_logic_vector(21534, 16),
25055 => conv_std_logic_vector(21631, 16),
25056 => conv_std_logic_vector(21728, 16),
25057 => conv_std_logic_vector(21825, 16),
25058 => conv_std_logic_vector(21922, 16),
25059 => conv_std_logic_vector(22019, 16),
25060 => conv_std_logic_vector(22116, 16),
25061 => conv_std_logic_vector(22213, 16),
25062 => conv_std_logic_vector(22310, 16),
25063 => conv_std_logic_vector(22407, 16),
25064 => conv_std_logic_vector(22504, 16),
25065 => conv_std_logic_vector(22601, 16),
25066 => conv_std_logic_vector(22698, 16),
25067 => conv_std_logic_vector(22795, 16),
25068 => conv_std_logic_vector(22892, 16),
25069 => conv_std_logic_vector(22989, 16),
25070 => conv_std_logic_vector(23086, 16),
25071 => conv_std_logic_vector(23183, 16),
25072 => conv_std_logic_vector(23280, 16),
25073 => conv_std_logic_vector(23377, 16),
25074 => conv_std_logic_vector(23474, 16),
25075 => conv_std_logic_vector(23571, 16),
25076 => conv_std_logic_vector(23668, 16),
25077 => conv_std_logic_vector(23765, 16),
25078 => conv_std_logic_vector(23862, 16),
25079 => conv_std_logic_vector(23959, 16),
25080 => conv_std_logic_vector(24056, 16),
25081 => conv_std_logic_vector(24153, 16),
25082 => conv_std_logic_vector(24250, 16),
25083 => conv_std_logic_vector(24347, 16),
25084 => conv_std_logic_vector(24444, 16),
25085 => conv_std_logic_vector(24541, 16),
25086 => conv_std_logic_vector(24638, 16),
25087 => conv_std_logic_vector(24735, 16),
25088 => conv_std_logic_vector(0, 16),
25089 => conv_std_logic_vector(98, 16),
25090 => conv_std_logic_vector(196, 16),
25091 => conv_std_logic_vector(294, 16),
25092 => conv_std_logic_vector(392, 16),
25093 => conv_std_logic_vector(490, 16),
25094 => conv_std_logic_vector(588, 16),
25095 => conv_std_logic_vector(686, 16),
25096 => conv_std_logic_vector(784, 16),
25097 => conv_std_logic_vector(882, 16),
25098 => conv_std_logic_vector(980, 16),
25099 => conv_std_logic_vector(1078, 16),
25100 => conv_std_logic_vector(1176, 16),
25101 => conv_std_logic_vector(1274, 16),
25102 => conv_std_logic_vector(1372, 16),
25103 => conv_std_logic_vector(1470, 16),
25104 => conv_std_logic_vector(1568, 16),
25105 => conv_std_logic_vector(1666, 16),
25106 => conv_std_logic_vector(1764, 16),
25107 => conv_std_logic_vector(1862, 16),
25108 => conv_std_logic_vector(1960, 16),
25109 => conv_std_logic_vector(2058, 16),
25110 => conv_std_logic_vector(2156, 16),
25111 => conv_std_logic_vector(2254, 16),
25112 => conv_std_logic_vector(2352, 16),
25113 => conv_std_logic_vector(2450, 16),
25114 => conv_std_logic_vector(2548, 16),
25115 => conv_std_logic_vector(2646, 16),
25116 => conv_std_logic_vector(2744, 16),
25117 => conv_std_logic_vector(2842, 16),
25118 => conv_std_logic_vector(2940, 16),
25119 => conv_std_logic_vector(3038, 16),
25120 => conv_std_logic_vector(3136, 16),
25121 => conv_std_logic_vector(3234, 16),
25122 => conv_std_logic_vector(3332, 16),
25123 => conv_std_logic_vector(3430, 16),
25124 => conv_std_logic_vector(3528, 16),
25125 => conv_std_logic_vector(3626, 16),
25126 => conv_std_logic_vector(3724, 16),
25127 => conv_std_logic_vector(3822, 16),
25128 => conv_std_logic_vector(3920, 16),
25129 => conv_std_logic_vector(4018, 16),
25130 => conv_std_logic_vector(4116, 16),
25131 => conv_std_logic_vector(4214, 16),
25132 => conv_std_logic_vector(4312, 16),
25133 => conv_std_logic_vector(4410, 16),
25134 => conv_std_logic_vector(4508, 16),
25135 => conv_std_logic_vector(4606, 16),
25136 => conv_std_logic_vector(4704, 16),
25137 => conv_std_logic_vector(4802, 16),
25138 => conv_std_logic_vector(4900, 16),
25139 => conv_std_logic_vector(4998, 16),
25140 => conv_std_logic_vector(5096, 16),
25141 => conv_std_logic_vector(5194, 16),
25142 => conv_std_logic_vector(5292, 16),
25143 => conv_std_logic_vector(5390, 16),
25144 => conv_std_logic_vector(5488, 16),
25145 => conv_std_logic_vector(5586, 16),
25146 => conv_std_logic_vector(5684, 16),
25147 => conv_std_logic_vector(5782, 16),
25148 => conv_std_logic_vector(5880, 16),
25149 => conv_std_logic_vector(5978, 16),
25150 => conv_std_logic_vector(6076, 16),
25151 => conv_std_logic_vector(6174, 16),
25152 => conv_std_logic_vector(6272, 16),
25153 => conv_std_logic_vector(6370, 16),
25154 => conv_std_logic_vector(6468, 16),
25155 => conv_std_logic_vector(6566, 16),
25156 => conv_std_logic_vector(6664, 16),
25157 => conv_std_logic_vector(6762, 16),
25158 => conv_std_logic_vector(6860, 16),
25159 => conv_std_logic_vector(6958, 16),
25160 => conv_std_logic_vector(7056, 16),
25161 => conv_std_logic_vector(7154, 16),
25162 => conv_std_logic_vector(7252, 16),
25163 => conv_std_logic_vector(7350, 16),
25164 => conv_std_logic_vector(7448, 16),
25165 => conv_std_logic_vector(7546, 16),
25166 => conv_std_logic_vector(7644, 16),
25167 => conv_std_logic_vector(7742, 16),
25168 => conv_std_logic_vector(7840, 16),
25169 => conv_std_logic_vector(7938, 16),
25170 => conv_std_logic_vector(8036, 16),
25171 => conv_std_logic_vector(8134, 16),
25172 => conv_std_logic_vector(8232, 16),
25173 => conv_std_logic_vector(8330, 16),
25174 => conv_std_logic_vector(8428, 16),
25175 => conv_std_logic_vector(8526, 16),
25176 => conv_std_logic_vector(8624, 16),
25177 => conv_std_logic_vector(8722, 16),
25178 => conv_std_logic_vector(8820, 16),
25179 => conv_std_logic_vector(8918, 16),
25180 => conv_std_logic_vector(9016, 16),
25181 => conv_std_logic_vector(9114, 16),
25182 => conv_std_logic_vector(9212, 16),
25183 => conv_std_logic_vector(9310, 16),
25184 => conv_std_logic_vector(9408, 16),
25185 => conv_std_logic_vector(9506, 16),
25186 => conv_std_logic_vector(9604, 16),
25187 => conv_std_logic_vector(9702, 16),
25188 => conv_std_logic_vector(9800, 16),
25189 => conv_std_logic_vector(9898, 16),
25190 => conv_std_logic_vector(9996, 16),
25191 => conv_std_logic_vector(10094, 16),
25192 => conv_std_logic_vector(10192, 16),
25193 => conv_std_logic_vector(10290, 16),
25194 => conv_std_logic_vector(10388, 16),
25195 => conv_std_logic_vector(10486, 16),
25196 => conv_std_logic_vector(10584, 16),
25197 => conv_std_logic_vector(10682, 16),
25198 => conv_std_logic_vector(10780, 16),
25199 => conv_std_logic_vector(10878, 16),
25200 => conv_std_logic_vector(10976, 16),
25201 => conv_std_logic_vector(11074, 16),
25202 => conv_std_logic_vector(11172, 16),
25203 => conv_std_logic_vector(11270, 16),
25204 => conv_std_logic_vector(11368, 16),
25205 => conv_std_logic_vector(11466, 16),
25206 => conv_std_logic_vector(11564, 16),
25207 => conv_std_logic_vector(11662, 16),
25208 => conv_std_logic_vector(11760, 16),
25209 => conv_std_logic_vector(11858, 16),
25210 => conv_std_logic_vector(11956, 16),
25211 => conv_std_logic_vector(12054, 16),
25212 => conv_std_logic_vector(12152, 16),
25213 => conv_std_logic_vector(12250, 16),
25214 => conv_std_logic_vector(12348, 16),
25215 => conv_std_logic_vector(12446, 16),
25216 => conv_std_logic_vector(12544, 16),
25217 => conv_std_logic_vector(12642, 16),
25218 => conv_std_logic_vector(12740, 16),
25219 => conv_std_logic_vector(12838, 16),
25220 => conv_std_logic_vector(12936, 16),
25221 => conv_std_logic_vector(13034, 16),
25222 => conv_std_logic_vector(13132, 16),
25223 => conv_std_logic_vector(13230, 16),
25224 => conv_std_logic_vector(13328, 16),
25225 => conv_std_logic_vector(13426, 16),
25226 => conv_std_logic_vector(13524, 16),
25227 => conv_std_logic_vector(13622, 16),
25228 => conv_std_logic_vector(13720, 16),
25229 => conv_std_logic_vector(13818, 16),
25230 => conv_std_logic_vector(13916, 16),
25231 => conv_std_logic_vector(14014, 16),
25232 => conv_std_logic_vector(14112, 16),
25233 => conv_std_logic_vector(14210, 16),
25234 => conv_std_logic_vector(14308, 16),
25235 => conv_std_logic_vector(14406, 16),
25236 => conv_std_logic_vector(14504, 16),
25237 => conv_std_logic_vector(14602, 16),
25238 => conv_std_logic_vector(14700, 16),
25239 => conv_std_logic_vector(14798, 16),
25240 => conv_std_logic_vector(14896, 16),
25241 => conv_std_logic_vector(14994, 16),
25242 => conv_std_logic_vector(15092, 16),
25243 => conv_std_logic_vector(15190, 16),
25244 => conv_std_logic_vector(15288, 16),
25245 => conv_std_logic_vector(15386, 16),
25246 => conv_std_logic_vector(15484, 16),
25247 => conv_std_logic_vector(15582, 16),
25248 => conv_std_logic_vector(15680, 16),
25249 => conv_std_logic_vector(15778, 16),
25250 => conv_std_logic_vector(15876, 16),
25251 => conv_std_logic_vector(15974, 16),
25252 => conv_std_logic_vector(16072, 16),
25253 => conv_std_logic_vector(16170, 16),
25254 => conv_std_logic_vector(16268, 16),
25255 => conv_std_logic_vector(16366, 16),
25256 => conv_std_logic_vector(16464, 16),
25257 => conv_std_logic_vector(16562, 16),
25258 => conv_std_logic_vector(16660, 16),
25259 => conv_std_logic_vector(16758, 16),
25260 => conv_std_logic_vector(16856, 16),
25261 => conv_std_logic_vector(16954, 16),
25262 => conv_std_logic_vector(17052, 16),
25263 => conv_std_logic_vector(17150, 16),
25264 => conv_std_logic_vector(17248, 16),
25265 => conv_std_logic_vector(17346, 16),
25266 => conv_std_logic_vector(17444, 16),
25267 => conv_std_logic_vector(17542, 16),
25268 => conv_std_logic_vector(17640, 16),
25269 => conv_std_logic_vector(17738, 16),
25270 => conv_std_logic_vector(17836, 16),
25271 => conv_std_logic_vector(17934, 16),
25272 => conv_std_logic_vector(18032, 16),
25273 => conv_std_logic_vector(18130, 16),
25274 => conv_std_logic_vector(18228, 16),
25275 => conv_std_logic_vector(18326, 16),
25276 => conv_std_logic_vector(18424, 16),
25277 => conv_std_logic_vector(18522, 16),
25278 => conv_std_logic_vector(18620, 16),
25279 => conv_std_logic_vector(18718, 16),
25280 => conv_std_logic_vector(18816, 16),
25281 => conv_std_logic_vector(18914, 16),
25282 => conv_std_logic_vector(19012, 16),
25283 => conv_std_logic_vector(19110, 16),
25284 => conv_std_logic_vector(19208, 16),
25285 => conv_std_logic_vector(19306, 16),
25286 => conv_std_logic_vector(19404, 16),
25287 => conv_std_logic_vector(19502, 16),
25288 => conv_std_logic_vector(19600, 16),
25289 => conv_std_logic_vector(19698, 16),
25290 => conv_std_logic_vector(19796, 16),
25291 => conv_std_logic_vector(19894, 16),
25292 => conv_std_logic_vector(19992, 16),
25293 => conv_std_logic_vector(20090, 16),
25294 => conv_std_logic_vector(20188, 16),
25295 => conv_std_logic_vector(20286, 16),
25296 => conv_std_logic_vector(20384, 16),
25297 => conv_std_logic_vector(20482, 16),
25298 => conv_std_logic_vector(20580, 16),
25299 => conv_std_logic_vector(20678, 16),
25300 => conv_std_logic_vector(20776, 16),
25301 => conv_std_logic_vector(20874, 16),
25302 => conv_std_logic_vector(20972, 16),
25303 => conv_std_logic_vector(21070, 16),
25304 => conv_std_logic_vector(21168, 16),
25305 => conv_std_logic_vector(21266, 16),
25306 => conv_std_logic_vector(21364, 16),
25307 => conv_std_logic_vector(21462, 16),
25308 => conv_std_logic_vector(21560, 16),
25309 => conv_std_logic_vector(21658, 16),
25310 => conv_std_logic_vector(21756, 16),
25311 => conv_std_logic_vector(21854, 16),
25312 => conv_std_logic_vector(21952, 16),
25313 => conv_std_logic_vector(22050, 16),
25314 => conv_std_logic_vector(22148, 16),
25315 => conv_std_logic_vector(22246, 16),
25316 => conv_std_logic_vector(22344, 16),
25317 => conv_std_logic_vector(22442, 16),
25318 => conv_std_logic_vector(22540, 16),
25319 => conv_std_logic_vector(22638, 16),
25320 => conv_std_logic_vector(22736, 16),
25321 => conv_std_logic_vector(22834, 16),
25322 => conv_std_logic_vector(22932, 16),
25323 => conv_std_logic_vector(23030, 16),
25324 => conv_std_logic_vector(23128, 16),
25325 => conv_std_logic_vector(23226, 16),
25326 => conv_std_logic_vector(23324, 16),
25327 => conv_std_logic_vector(23422, 16),
25328 => conv_std_logic_vector(23520, 16),
25329 => conv_std_logic_vector(23618, 16),
25330 => conv_std_logic_vector(23716, 16),
25331 => conv_std_logic_vector(23814, 16),
25332 => conv_std_logic_vector(23912, 16),
25333 => conv_std_logic_vector(24010, 16),
25334 => conv_std_logic_vector(24108, 16),
25335 => conv_std_logic_vector(24206, 16),
25336 => conv_std_logic_vector(24304, 16),
25337 => conv_std_logic_vector(24402, 16),
25338 => conv_std_logic_vector(24500, 16),
25339 => conv_std_logic_vector(24598, 16),
25340 => conv_std_logic_vector(24696, 16),
25341 => conv_std_logic_vector(24794, 16),
25342 => conv_std_logic_vector(24892, 16),
25343 => conv_std_logic_vector(24990, 16),
25344 => conv_std_logic_vector(0, 16),
25345 => conv_std_logic_vector(99, 16),
25346 => conv_std_logic_vector(198, 16),
25347 => conv_std_logic_vector(297, 16),
25348 => conv_std_logic_vector(396, 16),
25349 => conv_std_logic_vector(495, 16),
25350 => conv_std_logic_vector(594, 16),
25351 => conv_std_logic_vector(693, 16),
25352 => conv_std_logic_vector(792, 16),
25353 => conv_std_logic_vector(891, 16),
25354 => conv_std_logic_vector(990, 16),
25355 => conv_std_logic_vector(1089, 16),
25356 => conv_std_logic_vector(1188, 16),
25357 => conv_std_logic_vector(1287, 16),
25358 => conv_std_logic_vector(1386, 16),
25359 => conv_std_logic_vector(1485, 16),
25360 => conv_std_logic_vector(1584, 16),
25361 => conv_std_logic_vector(1683, 16),
25362 => conv_std_logic_vector(1782, 16),
25363 => conv_std_logic_vector(1881, 16),
25364 => conv_std_logic_vector(1980, 16),
25365 => conv_std_logic_vector(2079, 16),
25366 => conv_std_logic_vector(2178, 16),
25367 => conv_std_logic_vector(2277, 16),
25368 => conv_std_logic_vector(2376, 16),
25369 => conv_std_logic_vector(2475, 16),
25370 => conv_std_logic_vector(2574, 16),
25371 => conv_std_logic_vector(2673, 16),
25372 => conv_std_logic_vector(2772, 16),
25373 => conv_std_logic_vector(2871, 16),
25374 => conv_std_logic_vector(2970, 16),
25375 => conv_std_logic_vector(3069, 16),
25376 => conv_std_logic_vector(3168, 16),
25377 => conv_std_logic_vector(3267, 16),
25378 => conv_std_logic_vector(3366, 16),
25379 => conv_std_logic_vector(3465, 16),
25380 => conv_std_logic_vector(3564, 16),
25381 => conv_std_logic_vector(3663, 16),
25382 => conv_std_logic_vector(3762, 16),
25383 => conv_std_logic_vector(3861, 16),
25384 => conv_std_logic_vector(3960, 16),
25385 => conv_std_logic_vector(4059, 16),
25386 => conv_std_logic_vector(4158, 16),
25387 => conv_std_logic_vector(4257, 16),
25388 => conv_std_logic_vector(4356, 16),
25389 => conv_std_logic_vector(4455, 16),
25390 => conv_std_logic_vector(4554, 16),
25391 => conv_std_logic_vector(4653, 16),
25392 => conv_std_logic_vector(4752, 16),
25393 => conv_std_logic_vector(4851, 16),
25394 => conv_std_logic_vector(4950, 16),
25395 => conv_std_logic_vector(5049, 16),
25396 => conv_std_logic_vector(5148, 16),
25397 => conv_std_logic_vector(5247, 16),
25398 => conv_std_logic_vector(5346, 16),
25399 => conv_std_logic_vector(5445, 16),
25400 => conv_std_logic_vector(5544, 16),
25401 => conv_std_logic_vector(5643, 16),
25402 => conv_std_logic_vector(5742, 16),
25403 => conv_std_logic_vector(5841, 16),
25404 => conv_std_logic_vector(5940, 16),
25405 => conv_std_logic_vector(6039, 16),
25406 => conv_std_logic_vector(6138, 16),
25407 => conv_std_logic_vector(6237, 16),
25408 => conv_std_logic_vector(6336, 16),
25409 => conv_std_logic_vector(6435, 16),
25410 => conv_std_logic_vector(6534, 16),
25411 => conv_std_logic_vector(6633, 16),
25412 => conv_std_logic_vector(6732, 16),
25413 => conv_std_logic_vector(6831, 16),
25414 => conv_std_logic_vector(6930, 16),
25415 => conv_std_logic_vector(7029, 16),
25416 => conv_std_logic_vector(7128, 16),
25417 => conv_std_logic_vector(7227, 16),
25418 => conv_std_logic_vector(7326, 16),
25419 => conv_std_logic_vector(7425, 16),
25420 => conv_std_logic_vector(7524, 16),
25421 => conv_std_logic_vector(7623, 16),
25422 => conv_std_logic_vector(7722, 16),
25423 => conv_std_logic_vector(7821, 16),
25424 => conv_std_logic_vector(7920, 16),
25425 => conv_std_logic_vector(8019, 16),
25426 => conv_std_logic_vector(8118, 16),
25427 => conv_std_logic_vector(8217, 16),
25428 => conv_std_logic_vector(8316, 16),
25429 => conv_std_logic_vector(8415, 16),
25430 => conv_std_logic_vector(8514, 16),
25431 => conv_std_logic_vector(8613, 16),
25432 => conv_std_logic_vector(8712, 16),
25433 => conv_std_logic_vector(8811, 16),
25434 => conv_std_logic_vector(8910, 16),
25435 => conv_std_logic_vector(9009, 16),
25436 => conv_std_logic_vector(9108, 16),
25437 => conv_std_logic_vector(9207, 16),
25438 => conv_std_logic_vector(9306, 16),
25439 => conv_std_logic_vector(9405, 16),
25440 => conv_std_logic_vector(9504, 16),
25441 => conv_std_logic_vector(9603, 16),
25442 => conv_std_logic_vector(9702, 16),
25443 => conv_std_logic_vector(9801, 16),
25444 => conv_std_logic_vector(9900, 16),
25445 => conv_std_logic_vector(9999, 16),
25446 => conv_std_logic_vector(10098, 16),
25447 => conv_std_logic_vector(10197, 16),
25448 => conv_std_logic_vector(10296, 16),
25449 => conv_std_logic_vector(10395, 16),
25450 => conv_std_logic_vector(10494, 16),
25451 => conv_std_logic_vector(10593, 16),
25452 => conv_std_logic_vector(10692, 16),
25453 => conv_std_logic_vector(10791, 16),
25454 => conv_std_logic_vector(10890, 16),
25455 => conv_std_logic_vector(10989, 16),
25456 => conv_std_logic_vector(11088, 16),
25457 => conv_std_logic_vector(11187, 16),
25458 => conv_std_logic_vector(11286, 16),
25459 => conv_std_logic_vector(11385, 16),
25460 => conv_std_logic_vector(11484, 16),
25461 => conv_std_logic_vector(11583, 16),
25462 => conv_std_logic_vector(11682, 16),
25463 => conv_std_logic_vector(11781, 16),
25464 => conv_std_logic_vector(11880, 16),
25465 => conv_std_logic_vector(11979, 16),
25466 => conv_std_logic_vector(12078, 16),
25467 => conv_std_logic_vector(12177, 16),
25468 => conv_std_logic_vector(12276, 16),
25469 => conv_std_logic_vector(12375, 16),
25470 => conv_std_logic_vector(12474, 16),
25471 => conv_std_logic_vector(12573, 16),
25472 => conv_std_logic_vector(12672, 16),
25473 => conv_std_logic_vector(12771, 16),
25474 => conv_std_logic_vector(12870, 16),
25475 => conv_std_logic_vector(12969, 16),
25476 => conv_std_logic_vector(13068, 16),
25477 => conv_std_logic_vector(13167, 16),
25478 => conv_std_logic_vector(13266, 16),
25479 => conv_std_logic_vector(13365, 16),
25480 => conv_std_logic_vector(13464, 16),
25481 => conv_std_logic_vector(13563, 16),
25482 => conv_std_logic_vector(13662, 16),
25483 => conv_std_logic_vector(13761, 16),
25484 => conv_std_logic_vector(13860, 16),
25485 => conv_std_logic_vector(13959, 16),
25486 => conv_std_logic_vector(14058, 16),
25487 => conv_std_logic_vector(14157, 16),
25488 => conv_std_logic_vector(14256, 16),
25489 => conv_std_logic_vector(14355, 16),
25490 => conv_std_logic_vector(14454, 16),
25491 => conv_std_logic_vector(14553, 16),
25492 => conv_std_logic_vector(14652, 16),
25493 => conv_std_logic_vector(14751, 16),
25494 => conv_std_logic_vector(14850, 16),
25495 => conv_std_logic_vector(14949, 16),
25496 => conv_std_logic_vector(15048, 16),
25497 => conv_std_logic_vector(15147, 16),
25498 => conv_std_logic_vector(15246, 16),
25499 => conv_std_logic_vector(15345, 16),
25500 => conv_std_logic_vector(15444, 16),
25501 => conv_std_logic_vector(15543, 16),
25502 => conv_std_logic_vector(15642, 16),
25503 => conv_std_logic_vector(15741, 16),
25504 => conv_std_logic_vector(15840, 16),
25505 => conv_std_logic_vector(15939, 16),
25506 => conv_std_logic_vector(16038, 16),
25507 => conv_std_logic_vector(16137, 16),
25508 => conv_std_logic_vector(16236, 16),
25509 => conv_std_logic_vector(16335, 16),
25510 => conv_std_logic_vector(16434, 16),
25511 => conv_std_logic_vector(16533, 16),
25512 => conv_std_logic_vector(16632, 16),
25513 => conv_std_logic_vector(16731, 16),
25514 => conv_std_logic_vector(16830, 16),
25515 => conv_std_logic_vector(16929, 16),
25516 => conv_std_logic_vector(17028, 16),
25517 => conv_std_logic_vector(17127, 16),
25518 => conv_std_logic_vector(17226, 16),
25519 => conv_std_logic_vector(17325, 16),
25520 => conv_std_logic_vector(17424, 16),
25521 => conv_std_logic_vector(17523, 16),
25522 => conv_std_logic_vector(17622, 16),
25523 => conv_std_logic_vector(17721, 16),
25524 => conv_std_logic_vector(17820, 16),
25525 => conv_std_logic_vector(17919, 16),
25526 => conv_std_logic_vector(18018, 16),
25527 => conv_std_logic_vector(18117, 16),
25528 => conv_std_logic_vector(18216, 16),
25529 => conv_std_logic_vector(18315, 16),
25530 => conv_std_logic_vector(18414, 16),
25531 => conv_std_logic_vector(18513, 16),
25532 => conv_std_logic_vector(18612, 16),
25533 => conv_std_logic_vector(18711, 16),
25534 => conv_std_logic_vector(18810, 16),
25535 => conv_std_logic_vector(18909, 16),
25536 => conv_std_logic_vector(19008, 16),
25537 => conv_std_logic_vector(19107, 16),
25538 => conv_std_logic_vector(19206, 16),
25539 => conv_std_logic_vector(19305, 16),
25540 => conv_std_logic_vector(19404, 16),
25541 => conv_std_logic_vector(19503, 16),
25542 => conv_std_logic_vector(19602, 16),
25543 => conv_std_logic_vector(19701, 16),
25544 => conv_std_logic_vector(19800, 16),
25545 => conv_std_logic_vector(19899, 16),
25546 => conv_std_logic_vector(19998, 16),
25547 => conv_std_logic_vector(20097, 16),
25548 => conv_std_logic_vector(20196, 16),
25549 => conv_std_logic_vector(20295, 16),
25550 => conv_std_logic_vector(20394, 16),
25551 => conv_std_logic_vector(20493, 16),
25552 => conv_std_logic_vector(20592, 16),
25553 => conv_std_logic_vector(20691, 16),
25554 => conv_std_logic_vector(20790, 16),
25555 => conv_std_logic_vector(20889, 16),
25556 => conv_std_logic_vector(20988, 16),
25557 => conv_std_logic_vector(21087, 16),
25558 => conv_std_logic_vector(21186, 16),
25559 => conv_std_logic_vector(21285, 16),
25560 => conv_std_logic_vector(21384, 16),
25561 => conv_std_logic_vector(21483, 16),
25562 => conv_std_logic_vector(21582, 16),
25563 => conv_std_logic_vector(21681, 16),
25564 => conv_std_logic_vector(21780, 16),
25565 => conv_std_logic_vector(21879, 16),
25566 => conv_std_logic_vector(21978, 16),
25567 => conv_std_logic_vector(22077, 16),
25568 => conv_std_logic_vector(22176, 16),
25569 => conv_std_logic_vector(22275, 16),
25570 => conv_std_logic_vector(22374, 16),
25571 => conv_std_logic_vector(22473, 16),
25572 => conv_std_logic_vector(22572, 16),
25573 => conv_std_logic_vector(22671, 16),
25574 => conv_std_logic_vector(22770, 16),
25575 => conv_std_logic_vector(22869, 16),
25576 => conv_std_logic_vector(22968, 16),
25577 => conv_std_logic_vector(23067, 16),
25578 => conv_std_logic_vector(23166, 16),
25579 => conv_std_logic_vector(23265, 16),
25580 => conv_std_logic_vector(23364, 16),
25581 => conv_std_logic_vector(23463, 16),
25582 => conv_std_logic_vector(23562, 16),
25583 => conv_std_logic_vector(23661, 16),
25584 => conv_std_logic_vector(23760, 16),
25585 => conv_std_logic_vector(23859, 16),
25586 => conv_std_logic_vector(23958, 16),
25587 => conv_std_logic_vector(24057, 16),
25588 => conv_std_logic_vector(24156, 16),
25589 => conv_std_logic_vector(24255, 16),
25590 => conv_std_logic_vector(24354, 16),
25591 => conv_std_logic_vector(24453, 16),
25592 => conv_std_logic_vector(24552, 16),
25593 => conv_std_logic_vector(24651, 16),
25594 => conv_std_logic_vector(24750, 16),
25595 => conv_std_logic_vector(24849, 16),
25596 => conv_std_logic_vector(24948, 16),
25597 => conv_std_logic_vector(25047, 16),
25598 => conv_std_logic_vector(25146, 16),
25599 => conv_std_logic_vector(25245, 16),
25600 => conv_std_logic_vector(0, 16),
25601 => conv_std_logic_vector(100, 16),
25602 => conv_std_logic_vector(200, 16),
25603 => conv_std_logic_vector(300, 16),
25604 => conv_std_logic_vector(400, 16),
25605 => conv_std_logic_vector(500, 16),
25606 => conv_std_logic_vector(600, 16),
25607 => conv_std_logic_vector(700, 16),
25608 => conv_std_logic_vector(800, 16),
25609 => conv_std_logic_vector(900, 16),
25610 => conv_std_logic_vector(1000, 16),
25611 => conv_std_logic_vector(1100, 16),
25612 => conv_std_logic_vector(1200, 16),
25613 => conv_std_logic_vector(1300, 16),
25614 => conv_std_logic_vector(1400, 16),
25615 => conv_std_logic_vector(1500, 16),
25616 => conv_std_logic_vector(1600, 16),
25617 => conv_std_logic_vector(1700, 16),
25618 => conv_std_logic_vector(1800, 16),
25619 => conv_std_logic_vector(1900, 16),
25620 => conv_std_logic_vector(2000, 16),
25621 => conv_std_logic_vector(2100, 16),
25622 => conv_std_logic_vector(2200, 16),
25623 => conv_std_logic_vector(2300, 16),
25624 => conv_std_logic_vector(2400, 16),
25625 => conv_std_logic_vector(2500, 16),
25626 => conv_std_logic_vector(2600, 16),
25627 => conv_std_logic_vector(2700, 16),
25628 => conv_std_logic_vector(2800, 16),
25629 => conv_std_logic_vector(2900, 16),
25630 => conv_std_logic_vector(3000, 16),
25631 => conv_std_logic_vector(3100, 16),
25632 => conv_std_logic_vector(3200, 16),
25633 => conv_std_logic_vector(3300, 16),
25634 => conv_std_logic_vector(3400, 16),
25635 => conv_std_logic_vector(3500, 16),
25636 => conv_std_logic_vector(3600, 16),
25637 => conv_std_logic_vector(3700, 16),
25638 => conv_std_logic_vector(3800, 16),
25639 => conv_std_logic_vector(3900, 16),
25640 => conv_std_logic_vector(4000, 16),
25641 => conv_std_logic_vector(4100, 16),
25642 => conv_std_logic_vector(4200, 16),
25643 => conv_std_logic_vector(4300, 16),
25644 => conv_std_logic_vector(4400, 16),
25645 => conv_std_logic_vector(4500, 16),
25646 => conv_std_logic_vector(4600, 16),
25647 => conv_std_logic_vector(4700, 16),
25648 => conv_std_logic_vector(4800, 16),
25649 => conv_std_logic_vector(4900, 16),
25650 => conv_std_logic_vector(5000, 16),
25651 => conv_std_logic_vector(5100, 16),
25652 => conv_std_logic_vector(5200, 16),
25653 => conv_std_logic_vector(5300, 16),
25654 => conv_std_logic_vector(5400, 16),
25655 => conv_std_logic_vector(5500, 16),
25656 => conv_std_logic_vector(5600, 16),
25657 => conv_std_logic_vector(5700, 16),
25658 => conv_std_logic_vector(5800, 16),
25659 => conv_std_logic_vector(5900, 16),
25660 => conv_std_logic_vector(6000, 16),
25661 => conv_std_logic_vector(6100, 16),
25662 => conv_std_logic_vector(6200, 16),
25663 => conv_std_logic_vector(6300, 16),
25664 => conv_std_logic_vector(6400, 16),
25665 => conv_std_logic_vector(6500, 16),
25666 => conv_std_logic_vector(6600, 16),
25667 => conv_std_logic_vector(6700, 16),
25668 => conv_std_logic_vector(6800, 16),
25669 => conv_std_logic_vector(6900, 16),
25670 => conv_std_logic_vector(7000, 16),
25671 => conv_std_logic_vector(7100, 16),
25672 => conv_std_logic_vector(7200, 16),
25673 => conv_std_logic_vector(7300, 16),
25674 => conv_std_logic_vector(7400, 16),
25675 => conv_std_logic_vector(7500, 16),
25676 => conv_std_logic_vector(7600, 16),
25677 => conv_std_logic_vector(7700, 16),
25678 => conv_std_logic_vector(7800, 16),
25679 => conv_std_logic_vector(7900, 16),
25680 => conv_std_logic_vector(8000, 16),
25681 => conv_std_logic_vector(8100, 16),
25682 => conv_std_logic_vector(8200, 16),
25683 => conv_std_logic_vector(8300, 16),
25684 => conv_std_logic_vector(8400, 16),
25685 => conv_std_logic_vector(8500, 16),
25686 => conv_std_logic_vector(8600, 16),
25687 => conv_std_logic_vector(8700, 16),
25688 => conv_std_logic_vector(8800, 16),
25689 => conv_std_logic_vector(8900, 16),
25690 => conv_std_logic_vector(9000, 16),
25691 => conv_std_logic_vector(9100, 16),
25692 => conv_std_logic_vector(9200, 16),
25693 => conv_std_logic_vector(9300, 16),
25694 => conv_std_logic_vector(9400, 16),
25695 => conv_std_logic_vector(9500, 16),
25696 => conv_std_logic_vector(9600, 16),
25697 => conv_std_logic_vector(9700, 16),
25698 => conv_std_logic_vector(9800, 16),
25699 => conv_std_logic_vector(9900, 16),
25700 => conv_std_logic_vector(10000, 16),
25701 => conv_std_logic_vector(10100, 16),
25702 => conv_std_logic_vector(10200, 16),
25703 => conv_std_logic_vector(10300, 16),
25704 => conv_std_logic_vector(10400, 16),
25705 => conv_std_logic_vector(10500, 16),
25706 => conv_std_logic_vector(10600, 16),
25707 => conv_std_logic_vector(10700, 16),
25708 => conv_std_logic_vector(10800, 16),
25709 => conv_std_logic_vector(10900, 16),
25710 => conv_std_logic_vector(11000, 16),
25711 => conv_std_logic_vector(11100, 16),
25712 => conv_std_logic_vector(11200, 16),
25713 => conv_std_logic_vector(11300, 16),
25714 => conv_std_logic_vector(11400, 16),
25715 => conv_std_logic_vector(11500, 16),
25716 => conv_std_logic_vector(11600, 16),
25717 => conv_std_logic_vector(11700, 16),
25718 => conv_std_logic_vector(11800, 16),
25719 => conv_std_logic_vector(11900, 16),
25720 => conv_std_logic_vector(12000, 16),
25721 => conv_std_logic_vector(12100, 16),
25722 => conv_std_logic_vector(12200, 16),
25723 => conv_std_logic_vector(12300, 16),
25724 => conv_std_logic_vector(12400, 16),
25725 => conv_std_logic_vector(12500, 16),
25726 => conv_std_logic_vector(12600, 16),
25727 => conv_std_logic_vector(12700, 16),
25728 => conv_std_logic_vector(12800, 16),
25729 => conv_std_logic_vector(12900, 16),
25730 => conv_std_logic_vector(13000, 16),
25731 => conv_std_logic_vector(13100, 16),
25732 => conv_std_logic_vector(13200, 16),
25733 => conv_std_logic_vector(13300, 16),
25734 => conv_std_logic_vector(13400, 16),
25735 => conv_std_logic_vector(13500, 16),
25736 => conv_std_logic_vector(13600, 16),
25737 => conv_std_logic_vector(13700, 16),
25738 => conv_std_logic_vector(13800, 16),
25739 => conv_std_logic_vector(13900, 16),
25740 => conv_std_logic_vector(14000, 16),
25741 => conv_std_logic_vector(14100, 16),
25742 => conv_std_logic_vector(14200, 16),
25743 => conv_std_logic_vector(14300, 16),
25744 => conv_std_logic_vector(14400, 16),
25745 => conv_std_logic_vector(14500, 16),
25746 => conv_std_logic_vector(14600, 16),
25747 => conv_std_logic_vector(14700, 16),
25748 => conv_std_logic_vector(14800, 16),
25749 => conv_std_logic_vector(14900, 16),
25750 => conv_std_logic_vector(15000, 16),
25751 => conv_std_logic_vector(15100, 16),
25752 => conv_std_logic_vector(15200, 16),
25753 => conv_std_logic_vector(15300, 16),
25754 => conv_std_logic_vector(15400, 16),
25755 => conv_std_logic_vector(15500, 16),
25756 => conv_std_logic_vector(15600, 16),
25757 => conv_std_logic_vector(15700, 16),
25758 => conv_std_logic_vector(15800, 16),
25759 => conv_std_logic_vector(15900, 16),
25760 => conv_std_logic_vector(16000, 16),
25761 => conv_std_logic_vector(16100, 16),
25762 => conv_std_logic_vector(16200, 16),
25763 => conv_std_logic_vector(16300, 16),
25764 => conv_std_logic_vector(16400, 16),
25765 => conv_std_logic_vector(16500, 16),
25766 => conv_std_logic_vector(16600, 16),
25767 => conv_std_logic_vector(16700, 16),
25768 => conv_std_logic_vector(16800, 16),
25769 => conv_std_logic_vector(16900, 16),
25770 => conv_std_logic_vector(17000, 16),
25771 => conv_std_logic_vector(17100, 16),
25772 => conv_std_logic_vector(17200, 16),
25773 => conv_std_logic_vector(17300, 16),
25774 => conv_std_logic_vector(17400, 16),
25775 => conv_std_logic_vector(17500, 16),
25776 => conv_std_logic_vector(17600, 16),
25777 => conv_std_logic_vector(17700, 16),
25778 => conv_std_logic_vector(17800, 16),
25779 => conv_std_logic_vector(17900, 16),
25780 => conv_std_logic_vector(18000, 16),
25781 => conv_std_logic_vector(18100, 16),
25782 => conv_std_logic_vector(18200, 16),
25783 => conv_std_logic_vector(18300, 16),
25784 => conv_std_logic_vector(18400, 16),
25785 => conv_std_logic_vector(18500, 16),
25786 => conv_std_logic_vector(18600, 16),
25787 => conv_std_logic_vector(18700, 16),
25788 => conv_std_logic_vector(18800, 16),
25789 => conv_std_logic_vector(18900, 16),
25790 => conv_std_logic_vector(19000, 16),
25791 => conv_std_logic_vector(19100, 16),
25792 => conv_std_logic_vector(19200, 16),
25793 => conv_std_logic_vector(19300, 16),
25794 => conv_std_logic_vector(19400, 16),
25795 => conv_std_logic_vector(19500, 16),
25796 => conv_std_logic_vector(19600, 16),
25797 => conv_std_logic_vector(19700, 16),
25798 => conv_std_logic_vector(19800, 16),
25799 => conv_std_logic_vector(19900, 16),
25800 => conv_std_logic_vector(20000, 16),
25801 => conv_std_logic_vector(20100, 16),
25802 => conv_std_logic_vector(20200, 16),
25803 => conv_std_logic_vector(20300, 16),
25804 => conv_std_logic_vector(20400, 16),
25805 => conv_std_logic_vector(20500, 16),
25806 => conv_std_logic_vector(20600, 16),
25807 => conv_std_logic_vector(20700, 16),
25808 => conv_std_logic_vector(20800, 16),
25809 => conv_std_logic_vector(20900, 16),
25810 => conv_std_logic_vector(21000, 16),
25811 => conv_std_logic_vector(21100, 16),
25812 => conv_std_logic_vector(21200, 16),
25813 => conv_std_logic_vector(21300, 16),
25814 => conv_std_logic_vector(21400, 16),
25815 => conv_std_logic_vector(21500, 16),
25816 => conv_std_logic_vector(21600, 16),
25817 => conv_std_logic_vector(21700, 16),
25818 => conv_std_logic_vector(21800, 16),
25819 => conv_std_logic_vector(21900, 16),
25820 => conv_std_logic_vector(22000, 16),
25821 => conv_std_logic_vector(22100, 16),
25822 => conv_std_logic_vector(22200, 16),
25823 => conv_std_logic_vector(22300, 16),
25824 => conv_std_logic_vector(22400, 16),
25825 => conv_std_logic_vector(22500, 16),
25826 => conv_std_logic_vector(22600, 16),
25827 => conv_std_logic_vector(22700, 16),
25828 => conv_std_logic_vector(22800, 16),
25829 => conv_std_logic_vector(22900, 16),
25830 => conv_std_logic_vector(23000, 16),
25831 => conv_std_logic_vector(23100, 16),
25832 => conv_std_logic_vector(23200, 16),
25833 => conv_std_logic_vector(23300, 16),
25834 => conv_std_logic_vector(23400, 16),
25835 => conv_std_logic_vector(23500, 16),
25836 => conv_std_logic_vector(23600, 16),
25837 => conv_std_logic_vector(23700, 16),
25838 => conv_std_logic_vector(23800, 16),
25839 => conv_std_logic_vector(23900, 16),
25840 => conv_std_logic_vector(24000, 16),
25841 => conv_std_logic_vector(24100, 16),
25842 => conv_std_logic_vector(24200, 16),
25843 => conv_std_logic_vector(24300, 16),
25844 => conv_std_logic_vector(24400, 16),
25845 => conv_std_logic_vector(24500, 16),
25846 => conv_std_logic_vector(24600, 16),
25847 => conv_std_logic_vector(24700, 16),
25848 => conv_std_logic_vector(24800, 16),
25849 => conv_std_logic_vector(24900, 16),
25850 => conv_std_logic_vector(25000, 16),
25851 => conv_std_logic_vector(25100, 16),
25852 => conv_std_logic_vector(25200, 16),
25853 => conv_std_logic_vector(25300, 16),
25854 => conv_std_logic_vector(25400, 16),
25855 => conv_std_logic_vector(25500, 16),
25856 => conv_std_logic_vector(0, 16),
25857 => conv_std_logic_vector(101, 16),
25858 => conv_std_logic_vector(202, 16),
25859 => conv_std_logic_vector(303, 16),
25860 => conv_std_logic_vector(404, 16),
25861 => conv_std_logic_vector(505, 16),
25862 => conv_std_logic_vector(606, 16),
25863 => conv_std_logic_vector(707, 16),
25864 => conv_std_logic_vector(808, 16),
25865 => conv_std_logic_vector(909, 16),
25866 => conv_std_logic_vector(1010, 16),
25867 => conv_std_logic_vector(1111, 16),
25868 => conv_std_logic_vector(1212, 16),
25869 => conv_std_logic_vector(1313, 16),
25870 => conv_std_logic_vector(1414, 16),
25871 => conv_std_logic_vector(1515, 16),
25872 => conv_std_logic_vector(1616, 16),
25873 => conv_std_logic_vector(1717, 16),
25874 => conv_std_logic_vector(1818, 16),
25875 => conv_std_logic_vector(1919, 16),
25876 => conv_std_logic_vector(2020, 16),
25877 => conv_std_logic_vector(2121, 16),
25878 => conv_std_logic_vector(2222, 16),
25879 => conv_std_logic_vector(2323, 16),
25880 => conv_std_logic_vector(2424, 16),
25881 => conv_std_logic_vector(2525, 16),
25882 => conv_std_logic_vector(2626, 16),
25883 => conv_std_logic_vector(2727, 16),
25884 => conv_std_logic_vector(2828, 16),
25885 => conv_std_logic_vector(2929, 16),
25886 => conv_std_logic_vector(3030, 16),
25887 => conv_std_logic_vector(3131, 16),
25888 => conv_std_logic_vector(3232, 16),
25889 => conv_std_logic_vector(3333, 16),
25890 => conv_std_logic_vector(3434, 16),
25891 => conv_std_logic_vector(3535, 16),
25892 => conv_std_logic_vector(3636, 16),
25893 => conv_std_logic_vector(3737, 16),
25894 => conv_std_logic_vector(3838, 16),
25895 => conv_std_logic_vector(3939, 16),
25896 => conv_std_logic_vector(4040, 16),
25897 => conv_std_logic_vector(4141, 16),
25898 => conv_std_logic_vector(4242, 16),
25899 => conv_std_logic_vector(4343, 16),
25900 => conv_std_logic_vector(4444, 16),
25901 => conv_std_logic_vector(4545, 16),
25902 => conv_std_logic_vector(4646, 16),
25903 => conv_std_logic_vector(4747, 16),
25904 => conv_std_logic_vector(4848, 16),
25905 => conv_std_logic_vector(4949, 16),
25906 => conv_std_logic_vector(5050, 16),
25907 => conv_std_logic_vector(5151, 16),
25908 => conv_std_logic_vector(5252, 16),
25909 => conv_std_logic_vector(5353, 16),
25910 => conv_std_logic_vector(5454, 16),
25911 => conv_std_logic_vector(5555, 16),
25912 => conv_std_logic_vector(5656, 16),
25913 => conv_std_logic_vector(5757, 16),
25914 => conv_std_logic_vector(5858, 16),
25915 => conv_std_logic_vector(5959, 16),
25916 => conv_std_logic_vector(6060, 16),
25917 => conv_std_logic_vector(6161, 16),
25918 => conv_std_logic_vector(6262, 16),
25919 => conv_std_logic_vector(6363, 16),
25920 => conv_std_logic_vector(6464, 16),
25921 => conv_std_logic_vector(6565, 16),
25922 => conv_std_logic_vector(6666, 16),
25923 => conv_std_logic_vector(6767, 16),
25924 => conv_std_logic_vector(6868, 16),
25925 => conv_std_logic_vector(6969, 16),
25926 => conv_std_logic_vector(7070, 16),
25927 => conv_std_logic_vector(7171, 16),
25928 => conv_std_logic_vector(7272, 16),
25929 => conv_std_logic_vector(7373, 16),
25930 => conv_std_logic_vector(7474, 16),
25931 => conv_std_logic_vector(7575, 16),
25932 => conv_std_logic_vector(7676, 16),
25933 => conv_std_logic_vector(7777, 16),
25934 => conv_std_logic_vector(7878, 16),
25935 => conv_std_logic_vector(7979, 16),
25936 => conv_std_logic_vector(8080, 16),
25937 => conv_std_logic_vector(8181, 16),
25938 => conv_std_logic_vector(8282, 16),
25939 => conv_std_logic_vector(8383, 16),
25940 => conv_std_logic_vector(8484, 16),
25941 => conv_std_logic_vector(8585, 16),
25942 => conv_std_logic_vector(8686, 16),
25943 => conv_std_logic_vector(8787, 16),
25944 => conv_std_logic_vector(8888, 16),
25945 => conv_std_logic_vector(8989, 16),
25946 => conv_std_logic_vector(9090, 16),
25947 => conv_std_logic_vector(9191, 16),
25948 => conv_std_logic_vector(9292, 16),
25949 => conv_std_logic_vector(9393, 16),
25950 => conv_std_logic_vector(9494, 16),
25951 => conv_std_logic_vector(9595, 16),
25952 => conv_std_logic_vector(9696, 16),
25953 => conv_std_logic_vector(9797, 16),
25954 => conv_std_logic_vector(9898, 16),
25955 => conv_std_logic_vector(9999, 16),
25956 => conv_std_logic_vector(10100, 16),
25957 => conv_std_logic_vector(10201, 16),
25958 => conv_std_logic_vector(10302, 16),
25959 => conv_std_logic_vector(10403, 16),
25960 => conv_std_logic_vector(10504, 16),
25961 => conv_std_logic_vector(10605, 16),
25962 => conv_std_logic_vector(10706, 16),
25963 => conv_std_logic_vector(10807, 16),
25964 => conv_std_logic_vector(10908, 16),
25965 => conv_std_logic_vector(11009, 16),
25966 => conv_std_logic_vector(11110, 16),
25967 => conv_std_logic_vector(11211, 16),
25968 => conv_std_logic_vector(11312, 16),
25969 => conv_std_logic_vector(11413, 16),
25970 => conv_std_logic_vector(11514, 16),
25971 => conv_std_logic_vector(11615, 16),
25972 => conv_std_logic_vector(11716, 16),
25973 => conv_std_logic_vector(11817, 16),
25974 => conv_std_logic_vector(11918, 16),
25975 => conv_std_logic_vector(12019, 16),
25976 => conv_std_logic_vector(12120, 16),
25977 => conv_std_logic_vector(12221, 16),
25978 => conv_std_logic_vector(12322, 16),
25979 => conv_std_logic_vector(12423, 16),
25980 => conv_std_logic_vector(12524, 16),
25981 => conv_std_logic_vector(12625, 16),
25982 => conv_std_logic_vector(12726, 16),
25983 => conv_std_logic_vector(12827, 16),
25984 => conv_std_logic_vector(12928, 16),
25985 => conv_std_logic_vector(13029, 16),
25986 => conv_std_logic_vector(13130, 16),
25987 => conv_std_logic_vector(13231, 16),
25988 => conv_std_logic_vector(13332, 16),
25989 => conv_std_logic_vector(13433, 16),
25990 => conv_std_logic_vector(13534, 16),
25991 => conv_std_logic_vector(13635, 16),
25992 => conv_std_logic_vector(13736, 16),
25993 => conv_std_logic_vector(13837, 16),
25994 => conv_std_logic_vector(13938, 16),
25995 => conv_std_logic_vector(14039, 16),
25996 => conv_std_logic_vector(14140, 16),
25997 => conv_std_logic_vector(14241, 16),
25998 => conv_std_logic_vector(14342, 16),
25999 => conv_std_logic_vector(14443, 16),
26000 => conv_std_logic_vector(14544, 16),
26001 => conv_std_logic_vector(14645, 16),
26002 => conv_std_logic_vector(14746, 16),
26003 => conv_std_logic_vector(14847, 16),
26004 => conv_std_logic_vector(14948, 16),
26005 => conv_std_logic_vector(15049, 16),
26006 => conv_std_logic_vector(15150, 16),
26007 => conv_std_logic_vector(15251, 16),
26008 => conv_std_logic_vector(15352, 16),
26009 => conv_std_logic_vector(15453, 16),
26010 => conv_std_logic_vector(15554, 16),
26011 => conv_std_logic_vector(15655, 16),
26012 => conv_std_logic_vector(15756, 16),
26013 => conv_std_logic_vector(15857, 16),
26014 => conv_std_logic_vector(15958, 16),
26015 => conv_std_logic_vector(16059, 16),
26016 => conv_std_logic_vector(16160, 16),
26017 => conv_std_logic_vector(16261, 16),
26018 => conv_std_logic_vector(16362, 16),
26019 => conv_std_logic_vector(16463, 16),
26020 => conv_std_logic_vector(16564, 16),
26021 => conv_std_logic_vector(16665, 16),
26022 => conv_std_logic_vector(16766, 16),
26023 => conv_std_logic_vector(16867, 16),
26024 => conv_std_logic_vector(16968, 16),
26025 => conv_std_logic_vector(17069, 16),
26026 => conv_std_logic_vector(17170, 16),
26027 => conv_std_logic_vector(17271, 16),
26028 => conv_std_logic_vector(17372, 16),
26029 => conv_std_logic_vector(17473, 16),
26030 => conv_std_logic_vector(17574, 16),
26031 => conv_std_logic_vector(17675, 16),
26032 => conv_std_logic_vector(17776, 16),
26033 => conv_std_logic_vector(17877, 16),
26034 => conv_std_logic_vector(17978, 16),
26035 => conv_std_logic_vector(18079, 16),
26036 => conv_std_logic_vector(18180, 16),
26037 => conv_std_logic_vector(18281, 16),
26038 => conv_std_logic_vector(18382, 16),
26039 => conv_std_logic_vector(18483, 16),
26040 => conv_std_logic_vector(18584, 16),
26041 => conv_std_logic_vector(18685, 16),
26042 => conv_std_logic_vector(18786, 16),
26043 => conv_std_logic_vector(18887, 16),
26044 => conv_std_logic_vector(18988, 16),
26045 => conv_std_logic_vector(19089, 16),
26046 => conv_std_logic_vector(19190, 16),
26047 => conv_std_logic_vector(19291, 16),
26048 => conv_std_logic_vector(19392, 16),
26049 => conv_std_logic_vector(19493, 16),
26050 => conv_std_logic_vector(19594, 16),
26051 => conv_std_logic_vector(19695, 16),
26052 => conv_std_logic_vector(19796, 16),
26053 => conv_std_logic_vector(19897, 16),
26054 => conv_std_logic_vector(19998, 16),
26055 => conv_std_logic_vector(20099, 16),
26056 => conv_std_logic_vector(20200, 16),
26057 => conv_std_logic_vector(20301, 16),
26058 => conv_std_logic_vector(20402, 16),
26059 => conv_std_logic_vector(20503, 16),
26060 => conv_std_logic_vector(20604, 16),
26061 => conv_std_logic_vector(20705, 16),
26062 => conv_std_logic_vector(20806, 16),
26063 => conv_std_logic_vector(20907, 16),
26064 => conv_std_logic_vector(21008, 16),
26065 => conv_std_logic_vector(21109, 16),
26066 => conv_std_logic_vector(21210, 16),
26067 => conv_std_logic_vector(21311, 16),
26068 => conv_std_logic_vector(21412, 16),
26069 => conv_std_logic_vector(21513, 16),
26070 => conv_std_logic_vector(21614, 16),
26071 => conv_std_logic_vector(21715, 16),
26072 => conv_std_logic_vector(21816, 16),
26073 => conv_std_logic_vector(21917, 16),
26074 => conv_std_logic_vector(22018, 16),
26075 => conv_std_logic_vector(22119, 16),
26076 => conv_std_logic_vector(22220, 16),
26077 => conv_std_logic_vector(22321, 16),
26078 => conv_std_logic_vector(22422, 16),
26079 => conv_std_logic_vector(22523, 16),
26080 => conv_std_logic_vector(22624, 16),
26081 => conv_std_logic_vector(22725, 16),
26082 => conv_std_logic_vector(22826, 16),
26083 => conv_std_logic_vector(22927, 16),
26084 => conv_std_logic_vector(23028, 16),
26085 => conv_std_logic_vector(23129, 16),
26086 => conv_std_logic_vector(23230, 16),
26087 => conv_std_logic_vector(23331, 16),
26088 => conv_std_logic_vector(23432, 16),
26089 => conv_std_logic_vector(23533, 16),
26090 => conv_std_logic_vector(23634, 16),
26091 => conv_std_logic_vector(23735, 16),
26092 => conv_std_logic_vector(23836, 16),
26093 => conv_std_logic_vector(23937, 16),
26094 => conv_std_logic_vector(24038, 16),
26095 => conv_std_logic_vector(24139, 16),
26096 => conv_std_logic_vector(24240, 16),
26097 => conv_std_logic_vector(24341, 16),
26098 => conv_std_logic_vector(24442, 16),
26099 => conv_std_logic_vector(24543, 16),
26100 => conv_std_logic_vector(24644, 16),
26101 => conv_std_logic_vector(24745, 16),
26102 => conv_std_logic_vector(24846, 16),
26103 => conv_std_logic_vector(24947, 16),
26104 => conv_std_logic_vector(25048, 16),
26105 => conv_std_logic_vector(25149, 16),
26106 => conv_std_logic_vector(25250, 16),
26107 => conv_std_logic_vector(25351, 16),
26108 => conv_std_logic_vector(25452, 16),
26109 => conv_std_logic_vector(25553, 16),
26110 => conv_std_logic_vector(25654, 16),
26111 => conv_std_logic_vector(25755, 16),
26112 => conv_std_logic_vector(0, 16),
26113 => conv_std_logic_vector(102, 16),
26114 => conv_std_logic_vector(204, 16),
26115 => conv_std_logic_vector(306, 16),
26116 => conv_std_logic_vector(408, 16),
26117 => conv_std_logic_vector(510, 16),
26118 => conv_std_logic_vector(612, 16),
26119 => conv_std_logic_vector(714, 16),
26120 => conv_std_logic_vector(816, 16),
26121 => conv_std_logic_vector(918, 16),
26122 => conv_std_logic_vector(1020, 16),
26123 => conv_std_logic_vector(1122, 16),
26124 => conv_std_logic_vector(1224, 16),
26125 => conv_std_logic_vector(1326, 16),
26126 => conv_std_logic_vector(1428, 16),
26127 => conv_std_logic_vector(1530, 16),
26128 => conv_std_logic_vector(1632, 16),
26129 => conv_std_logic_vector(1734, 16),
26130 => conv_std_logic_vector(1836, 16),
26131 => conv_std_logic_vector(1938, 16),
26132 => conv_std_logic_vector(2040, 16),
26133 => conv_std_logic_vector(2142, 16),
26134 => conv_std_logic_vector(2244, 16),
26135 => conv_std_logic_vector(2346, 16),
26136 => conv_std_logic_vector(2448, 16),
26137 => conv_std_logic_vector(2550, 16),
26138 => conv_std_logic_vector(2652, 16),
26139 => conv_std_logic_vector(2754, 16),
26140 => conv_std_logic_vector(2856, 16),
26141 => conv_std_logic_vector(2958, 16),
26142 => conv_std_logic_vector(3060, 16),
26143 => conv_std_logic_vector(3162, 16),
26144 => conv_std_logic_vector(3264, 16),
26145 => conv_std_logic_vector(3366, 16),
26146 => conv_std_logic_vector(3468, 16),
26147 => conv_std_logic_vector(3570, 16),
26148 => conv_std_logic_vector(3672, 16),
26149 => conv_std_logic_vector(3774, 16),
26150 => conv_std_logic_vector(3876, 16),
26151 => conv_std_logic_vector(3978, 16),
26152 => conv_std_logic_vector(4080, 16),
26153 => conv_std_logic_vector(4182, 16),
26154 => conv_std_logic_vector(4284, 16),
26155 => conv_std_logic_vector(4386, 16),
26156 => conv_std_logic_vector(4488, 16),
26157 => conv_std_logic_vector(4590, 16),
26158 => conv_std_logic_vector(4692, 16),
26159 => conv_std_logic_vector(4794, 16),
26160 => conv_std_logic_vector(4896, 16),
26161 => conv_std_logic_vector(4998, 16),
26162 => conv_std_logic_vector(5100, 16),
26163 => conv_std_logic_vector(5202, 16),
26164 => conv_std_logic_vector(5304, 16),
26165 => conv_std_logic_vector(5406, 16),
26166 => conv_std_logic_vector(5508, 16),
26167 => conv_std_logic_vector(5610, 16),
26168 => conv_std_logic_vector(5712, 16),
26169 => conv_std_logic_vector(5814, 16),
26170 => conv_std_logic_vector(5916, 16),
26171 => conv_std_logic_vector(6018, 16),
26172 => conv_std_logic_vector(6120, 16),
26173 => conv_std_logic_vector(6222, 16),
26174 => conv_std_logic_vector(6324, 16),
26175 => conv_std_logic_vector(6426, 16),
26176 => conv_std_logic_vector(6528, 16),
26177 => conv_std_logic_vector(6630, 16),
26178 => conv_std_logic_vector(6732, 16),
26179 => conv_std_logic_vector(6834, 16),
26180 => conv_std_logic_vector(6936, 16),
26181 => conv_std_logic_vector(7038, 16),
26182 => conv_std_logic_vector(7140, 16),
26183 => conv_std_logic_vector(7242, 16),
26184 => conv_std_logic_vector(7344, 16),
26185 => conv_std_logic_vector(7446, 16),
26186 => conv_std_logic_vector(7548, 16),
26187 => conv_std_logic_vector(7650, 16),
26188 => conv_std_logic_vector(7752, 16),
26189 => conv_std_logic_vector(7854, 16),
26190 => conv_std_logic_vector(7956, 16),
26191 => conv_std_logic_vector(8058, 16),
26192 => conv_std_logic_vector(8160, 16),
26193 => conv_std_logic_vector(8262, 16),
26194 => conv_std_logic_vector(8364, 16),
26195 => conv_std_logic_vector(8466, 16),
26196 => conv_std_logic_vector(8568, 16),
26197 => conv_std_logic_vector(8670, 16),
26198 => conv_std_logic_vector(8772, 16),
26199 => conv_std_logic_vector(8874, 16),
26200 => conv_std_logic_vector(8976, 16),
26201 => conv_std_logic_vector(9078, 16),
26202 => conv_std_logic_vector(9180, 16),
26203 => conv_std_logic_vector(9282, 16),
26204 => conv_std_logic_vector(9384, 16),
26205 => conv_std_logic_vector(9486, 16),
26206 => conv_std_logic_vector(9588, 16),
26207 => conv_std_logic_vector(9690, 16),
26208 => conv_std_logic_vector(9792, 16),
26209 => conv_std_logic_vector(9894, 16),
26210 => conv_std_logic_vector(9996, 16),
26211 => conv_std_logic_vector(10098, 16),
26212 => conv_std_logic_vector(10200, 16),
26213 => conv_std_logic_vector(10302, 16),
26214 => conv_std_logic_vector(10404, 16),
26215 => conv_std_logic_vector(10506, 16),
26216 => conv_std_logic_vector(10608, 16),
26217 => conv_std_logic_vector(10710, 16),
26218 => conv_std_logic_vector(10812, 16),
26219 => conv_std_logic_vector(10914, 16),
26220 => conv_std_logic_vector(11016, 16),
26221 => conv_std_logic_vector(11118, 16),
26222 => conv_std_logic_vector(11220, 16),
26223 => conv_std_logic_vector(11322, 16),
26224 => conv_std_logic_vector(11424, 16),
26225 => conv_std_logic_vector(11526, 16),
26226 => conv_std_logic_vector(11628, 16),
26227 => conv_std_logic_vector(11730, 16),
26228 => conv_std_logic_vector(11832, 16),
26229 => conv_std_logic_vector(11934, 16),
26230 => conv_std_logic_vector(12036, 16),
26231 => conv_std_logic_vector(12138, 16),
26232 => conv_std_logic_vector(12240, 16),
26233 => conv_std_logic_vector(12342, 16),
26234 => conv_std_logic_vector(12444, 16),
26235 => conv_std_logic_vector(12546, 16),
26236 => conv_std_logic_vector(12648, 16),
26237 => conv_std_logic_vector(12750, 16),
26238 => conv_std_logic_vector(12852, 16),
26239 => conv_std_logic_vector(12954, 16),
26240 => conv_std_logic_vector(13056, 16),
26241 => conv_std_logic_vector(13158, 16),
26242 => conv_std_logic_vector(13260, 16),
26243 => conv_std_logic_vector(13362, 16),
26244 => conv_std_logic_vector(13464, 16),
26245 => conv_std_logic_vector(13566, 16),
26246 => conv_std_logic_vector(13668, 16),
26247 => conv_std_logic_vector(13770, 16),
26248 => conv_std_logic_vector(13872, 16),
26249 => conv_std_logic_vector(13974, 16),
26250 => conv_std_logic_vector(14076, 16),
26251 => conv_std_logic_vector(14178, 16),
26252 => conv_std_logic_vector(14280, 16),
26253 => conv_std_logic_vector(14382, 16),
26254 => conv_std_logic_vector(14484, 16),
26255 => conv_std_logic_vector(14586, 16),
26256 => conv_std_logic_vector(14688, 16),
26257 => conv_std_logic_vector(14790, 16),
26258 => conv_std_logic_vector(14892, 16),
26259 => conv_std_logic_vector(14994, 16),
26260 => conv_std_logic_vector(15096, 16),
26261 => conv_std_logic_vector(15198, 16),
26262 => conv_std_logic_vector(15300, 16),
26263 => conv_std_logic_vector(15402, 16),
26264 => conv_std_logic_vector(15504, 16),
26265 => conv_std_logic_vector(15606, 16),
26266 => conv_std_logic_vector(15708, 16),
26267 => conv_std_logic_vector(15810, 16),
26268 => conv_std_logic_vector(15912, 16),
26269 => conv_std_logic_vector(16014, 16),
26270 => conv_std_logic_vector(16116, 16),
26271 => conv_std_logic_vector(16218, 16),
26272 => conv_std_logic_vector(16320, 16),
26273 => conv_std_logic_vector(16422, 16),
26274 => conv_std_logic_vector(16524, 16),
26275 => conv_std_logic_vector(16626, 16),
26276 => conv_std_logic_vector(16728, 16),
26277 => conv_std_logic_vector(16830, 16),
26278 => conv_std_logic_vector(16932, 16),
26279 => conv_std_logic_vector(17034, 16),
26280 => conv_std_logic_vector(17136, 16),
26281 => conv_std_logic_vector(17238, 16),
26282 => conv_std_logic_vector(17340, 16),
26283 => conv_std_logic_vector(17442, 16),
26284 => conv_std_logic_vector(17544, 16),
26285 => conv_std_logic_vector(17646, 16),
26286 => conv_std_logic_vector(17748, 16),
26287 => conv_std_logic_vector(17850, 16),
26288 => conv_std_logic_vector(17952, 16),
26289 => conv_std_logic_vector(18054, 16),
26290 => conv_std_logic_vector(18156, 16),
26291 => conv_std_logic_vector(18258, 16),
26292 => conv_std_logic_vector(18360, 16),
26293 => conv_std_logic_vector(18462, 16),
26294 => conv_std_logic_vector(18564, 16),
26295 => conv_std_logic_vector(18666, 16),
26296 => conv_std_logic_vector(18768, 16),
26297 => conv_std_logic_vector(18870, 16),
26298 => conv_std_logic_vector(18972, 16),
26299 => conv_std_logic_vector(19074, 16),
26300 => conv_std_logic_vector(19176, 16),
26301 => conv_std_logic_vector(19278, 16),
26302 => conv_std_logic_vector(19380, 16),
26303 => conv_std_logic_vector(19482, 16),
26304 => conv_std_logic_vector(19584, 16),
26305 => conv_std_logic_vector(19686, 16),
26306 => conv_std_logic_vector(19788, 16),
26307 => conv_std_logic_vector(19890, 16),
26308 => conv_std_logic_vector(19992, 16),
26309 => conv_std_logic_vector(20094, 16),
26310 => conv_std_logic_vector(20196, 16),
26311 => conv_std_logic_vector(20298, 16),
26312 => conv_std_logic_vector(20400, 16),
26313 => conv_std_logic_vector(20502, 16),
26314 => conv_std_logic_vector(20604, 16),
26315 => conv_std_logic_vector(20706, 16),
26316 => conv_std_logic_vector(20808, 16),
26317 => conv_std_logic_vector(20910, 16),
26318 => conv_std_logic_vector(21012, 16),
26319 => conv_std_logic_vector(21114, 16),
26320 => conv_std_logic_vector(21216, 16),
26321 => conv_std_logic_vector(21318, 16),
26322 => conv_std_logic_vector(21420, 16),
26323 => conv_std_logic_vector(21522, 16),
26324 => conv_std_logic_vector(21624, 16),
26325 => conv_std_logic_vector(21726, 16),
26326 => conv_std_logic_vector(21828, 16),
26327 => conv_std_logic_vector(21930, 16),
26328 => conv_std_logic_vector(22032, 16),
26329 => conv_std_logic_vector(22134, 16),
26330 => conv_std_logic_vector(22236, 16),
26331 => conv_std_logic_vector(22338, 16),
26332 => conv_std_logic_vector(22440, 16),
26333 => conv_std_logic_vector(22542, 16),
26334 => conv_std_logic_vector(22644, 16),
26335 => conv_std_logic_vector(22746, 16),
26336 => conv_std_logic_vector(22848, 16),
26337 => conv_std_logic_vector(22950, 16),
26338 => conv_std_logic_vector(23052, 16),
26339 => conv_std_logic_vector(23154, 16),
26340 => conv_std_logic_vector(23256, 16),
26341 => conv_std_logic_vector(23358, 16),
26342 => conv_std_logic_vector(23460, 16),
26343 => conv_std_logic_vector(23562, 16),
26344 => conv_std_logic_vector(23664, 16),
26345 => conv_std_logic_vector(23766, 16),
26346 => conv_std_logic_vector(23868, 16),
26347 => conv_std_logic_vector(23970, 16),
26348 => conv_std_logic_vector(24072, 16),
26349 => conv_std_logic_vector(24174, 16),
26350 => conv_std_logic_vector(24276, 16),
26351 => conv_std_logic_vector(24378, 16),
26352 => conv_std_logic_vector(24480, 16),
26353 => conv_std_logic_vector(24582, 16),
26354 => conv_std_logic_vector(24684, 16),
26355 => conv_std_logic_vector(24786, 16),
26356 => conv_std_logic_vector(24888, 16),
26357 => conv_std_logic_vector(24990, 16),
26358 => conv_std_logic_vector(25092, 16),
26359 => conv_std_logic_vector(25194, 16),
26360 => conv_std_logic_vector(25296, 16),
26361 => conv_std_logic_vector(25398, 16),
26362 => conv_std_logic_vector(25500, 16),
26363 => conv_std_logic_vector(25602, 16),
26364 => conv_std_logic_vector(25704, 16),
26365 => conv_std_logic_vector(25806, 16),
26366 => conv_std_logic_vector(25908, 16),
26367 => conv_std_logic_vector(26010, 16),
26368 => conv_std_logic_vector(0, 16),
26369 => conv_std_logic_vector(103, 16),
26370 => conv_std_logic_vector(206, 16),
26371 => conv_std_logic_vector(309, 16),
26372 => conv_std_logic_vector(412, 16),
26373 => conv_std_logic_vector(515, 16),
26374 => conv_std_logic_vector(618, 16),
26375 => conv_std_logic_vector(721, 16),
26376 => conv_std_logic_vector(824, 16),
26377 => conv_std_logic_vector(927, 16),
26378 => conv_std_logic_vector(1030, 16),
26379 => conv_std_logic_vector(1133, 16),
26380 => conv_std_logic_vector(1236, 16),
26381 => conv_std_logic_vector(1339, 16),
26382 => conv_std_logic_vector(1442, 16),
26383 => conv_std_logic_vector(1545, 16),
26384 => conv_std_logic_vector(1648, 16),
26385 => conv_std_logic_vector(1751, 16),
26386 => conv_std_logic_vector(1854, 16),
26387 => conv_std_logic_vector(1957, 16),
26388 => conv_std_logic_vector(2060, 16),
26389 => conv_std_logic_vector(2163, 16),
26390 => conv_std_logic_vector(2266, 16),
26391 => conv_std_logic_vector(2369, 16),
26392 => conv_std_logic_vector(2472, 16),
26393 => conv_std_logic_vector(2575, 16),
26394 => conv_std_logic_vector(2678, 16),
26395 => conv_std_logic_vector(2781, 16),
26396 => conv_std_logic_vector(2884, 16),
26397 => conv_std_logic_vector(2987, 16),
26398 => conv_std_logic_vector(3090, 16),
26399 => conv_std_logic_vector(3193, 16),
26400 => conv_std_logic_vector(3296, 16),
26401 => conv_std_logic_vector(3399, 16),
26402 => conv_std_logic_vector(3502, 16),
26403 => conv_std_logic_vector(3605, 16),
26404 => conv_std_logic_vector(3708, 16),
26405 => conv_std_logic_vector(3811, 16),
26406 => conv_std_logic_vector(3914, 16),
26407 => conv_std_logic_vector(4017, 16),
26408 => conv_std_logic_vector(4120, 16),
26409 => conv_std_logic_vector(4223, 16),
26410 => conv_std_logic_vector(4326, 16),
26411 => conv_std_logic_vector(4429, 16),
26412 => conv_std_logic_vector(4532, 16),
26413 => conv_std_logic_vector(4635, 16),
26414 => conv_std_logic_vector(4738, 16),
26415 => conv_std_logic_vector(4841, 16),
26416 => conv_std_logic_vector(4944, 16),
26417 => conv_std_logic_vector(5047, 16),
26418 => conv_std_logic_vector(5150, 16),
26419 => conv_std_logic_vector(5253, 16),
26420 => conv_std_logic_vector(5356, 16),
26421 => conv_std_logic_vector(5459, 16),
26422 => conv_std_logic_vector(5562, 16),
26423 => conv_std_logic_vector(5665, 16),
26424 => conv_std_logic_vector(5768, 16),
26425 => conv_std_logic_vector(5871, 16),
26426 => conv_std_logic_vector(5974, 16),
26427 => conv_std_logic_vector(6077, 16),
26428 => conv_std_logic_vector(6180, 16),
26429 => conv_std_logic_vector(6283, 16),
26430 => conv_std_logic_vector(6386, 16),
26431 => conv_std_logic_vector(6489, 16),
26432 => conv_std_logic_vector(6592, 16),
26433 => conv_std_logic_vector(6695, 16),
26434 => conv_std_logic_vector(6798, 16),
26435 => conv_std_logic_vector(6901, 16),
26436 => conv_std_logic_vector(7004, 16),
26437 => conv_std_logic_vector(7107, 16),
26438 => conv_std_logic_vector(7210, 16),
26439 => conv_std_logic_vector(7313, 16),
26440 => conv_std_logic_vector(7416, 16),
26441 => conv_std_logic_vector(7519, 16),
26442 => conv_std_logic_vector(7622, 16),
26443 => conv_std_logic_vector(7725, 16),
26444 => conv_std_logic_vector(7828, 16),
26445 => conv_std_logic_vector(7931, 16),
26446 => conv_std_logic_vector(8034, 16),
26447 => conv_std_logic_vector(8137, 16),
26448 => conv_std_logic_vector(8240, 16),
26449 => conv_std_logic_vector(8343, 16),
26450 => conv_std_logic_vector(8446, 16),
26451 => conv_std_logic_vector(8549, 16),
26452 => conv_std_logic_vector(8652, 16),
26453 => conv_std_logic_vector(8755, 16),
26454 => conv_std_logic_vector(8858, 16),
26455 => conv_std_logic_vector(8961, 16),
26456 => conv_std_logic_vector(9064, 16),
26457 => conv_std_logic_vector(9167, 16),
26458 => conv_std_logic_vector(9270, 16),
26459 => conv_std_logic_vector(9373, 16),
26460 => conv_std_logic_vector(9476, 16),
26461 => conv_std_logic_vector(9579, 16),
26462 => conv_std_logic_vector(9682, 16),
26463 => conv_std_logic_vector(9785, 16),
26464 => conv_std_logic_vector(9888, 16),
26465 => conv_std_logic_vector(9991, 16),
26466 => conv_std_logic_vector(10094, 16),
26467 => conv_std_logic_vector(10197, 16),
26468 => conv_std_logic_vector(10300, 16),
26469 => conv_std_logic_vector(10403, 16),
26470 => conv_std_logic_vector(10506, 16),
26471 => conv_std_logic_vector(10609, 16),
26472 => conv_std_logic_vector(10712, 16),
26473 => conv_std_logic_vector(10815, 16),
26474 => conv_std_logic_vector(10918, 16),
26475 => conv_std_logic_vector(11021, 16),
26476 => conv_std_logic_vector(11124, 16),
26477 => conv_std_logic_vector(11227, 16),
26478 => conv_std_logic_vector(11330, 16),
26479 => conv_std_logic_vector(11433, 16),
26480 => conv_std_logic_vector(11536, 16),
26481 => conv_std_logic_vector(11639, 16),
26482 => conv_std_logic_vector(11742, 16),
26483 => conv_std_logic_vector(11845, 16),
26484 => conv_std_logic_vector(11948, 16),
26485 => conv_std_logic_vector(12051, 16),
26486 => conv_std_logic_vector(12154, 16),
26487 => conv_std_logic_vector(12257, 16),
26488 => conv_std_logic_vector(12360, 16),
26489 => conv_std_logic_vector(12463, 16),
26490 => conv_std_logic_vector(12566, 16),
26491 => conv_std_logic_vector(12669, 16),
26492 => conv_std_logic_vector(12772, 16),
26493 => conv_std_logic_vector(12875, 16),
26494 => conv_std_logic_vector(12978, 16),
26495 => conv_std_logic_vector(13081, 16),
26496 => conv_std_logic_vector(13184, 16),
26497 => conv_std_logic_vector(13287, 16),
26498 => conv_std_logic_vector(13390, 16),
26499 => conv_std_logic_vector(13493, 16),
26500 => conv_std_logic_vector(13596, 16),
26501 => conv_std_logic_vector(13699, 16),
26502 => conv_std_logic_vector(13802, 16),
26503 => conv_std_logic_vector(13905, 16),
26504 => conv_std_logic_vector(14008, 16),
26505 => conv_std_logic_vector(14111, 16),
26506 => conv_std_logic_vector(14214, 16),
26507 => conv_std_logic_vector(14317, 16),
26508 => conv_std_logic_vector(14420, 16),
26509 => conv_std_logic_vector(14523, 16),
26510 => conv_std_logic_vector(14626, 16),
26511 => conv_std_logic_vector(14729, 16),
26512 => conv_std_logic_vector(14832, 16),
26513 => conv_std_logic_vector(14935, 16),
26514 => conv_std_logic_vector(15038, 16),
26515 => conv_std_logic_vector(15141, 16),
26516 => conv_std_logic_vector(15244, 16),
26517 => conv_std_logic_vector(15347, 16),
26518 => conv_std_logic_vector(15450, 16),
26519 => conv_std_logic_vector(15553, 16),
26520 => conv_std_logic_vector(15656, 16),
26521 => conv_std_logic_vector(15759, 16),
26522 => conv_std_logic_vector(15862, 16),
26523 => conv_std_logic_vector(15965, 16),
26524 => conv_std_logic_vector(16068, 16),
26525 => conv_std_logic_vector(16171, 16),
26526 => conv_std_logic_vector(16274, 16),
26527 => conv_std_logic_vector(16377, 16),
26528 => conv_std_logic_vector(16480, 16),
26529 => conv_std_logic_vector(16583, 16),
26530 => conv_std_logic_vector(16686, 16),
26531 => conv_std_logic_vector(16789, 16),
26532 => conv_std_logic_vector(16892, 16),
26533 => conv_std_logic_vector(16995, 16),
26534 => conv_std_logic_vector(17098, 16),
26535 => conv_std_logic_vector(17201, 16),
26536 => conv_std_logic_vector(17304, 16),
26537 => conv_std_logic_vector(17407, 16),
26538 => conv_std_logic_vector(17510, 16),
26539 => conv_std_logic_vector(17613, 16),
26540 => conv_std_logic_vector(17716, 16),
26541 => conv_std_logic_vector(17819, 16),
26542 => conv_std_logic_vector(17922, 16),
26543 => conv_std_logic_vector(18025, 16),
26544 => conv_std_logic_vector(18128, 16),
26545 => conv_std_logic_vector(18231, 16),
26546 => conv_std_logic_vector(18334, 16),
26547 => conv_std_logic_vector(18437, 16),
26548 => conv_std_logic_vector(18540, 16),
26549 => conv_std_logic_vector(18643, 16),
26550 => conv_std_logic_vector(18746, 16),
26551 => conv_std_logic_vector(18849, 16),
26552 => conv_std_logic_vector(18952, 16),
26553 => conv_std_logic_vector(19055, 16),
26554 => conv_std_logic_vector(19158, 16),
26555 => conv_std_logic_vector(19261, 16),
26556 => conv_std_logic_vector(19364, 16),
26557 => conv_std_logic_vector(19467, 16),
26558 => conv_std_logic_vector(19570, 16),
26559 => conv_std_logic_vector(19673, 16),
26560 => conv_std_logic_vector(19776, 16),
26561 => conv_std_logic_vector(19879, 16),
26562 => conv_std_logic_vector(19982, 16),
26563 => conv_std_logic_vector(20085, 16),
26564 => conv_std_logic_vector(20188, 16),
26565 => conv_std_logic_vector(20291, 16),
26566 => conv_std_logic_vector(20394, 16),
26567 => conv_std_logic_vector(20497, 16),
26568 => conv_std_logic_vector(20600, 16),
26569 => conv_std_logic_vector(20703, 16),
26570 => conv_std_logic_vector(20806, 16),
26571 => conv_std_logic_vector(20909, 16),
26572 => conv_std_logic_vector(21012, 16),
26573 => conv_std_logic_vector(21115, 16),
26574 => conv_std_logic_vector(21218, 16),
26575 => conv_std_logic_vector(21321, 16),
26576 => conv_std_logic_vector(21424, 16),
26577 => conv_std_logic_vector(21527, 16),
26578 => conv_std_logic_vector(21630, 16),
26579 => conv_std_logic_vector(21733, 16),
26580 => conv_std_logic_vector(21836, 16),
26581 => conv_std_logic_vector(21939, 16),
26582 => conv_std_logic_vector(22042, 16),
26583 => conv_std_logic_vector(22145, 16),
26584 => conv_std_logic_vector(22248, 16),
26585 => conv_std_logic_vector(22351, 16),
26586 => conv_std_logic_vector(22454, 16),
26587 => conv_std_logic_vector(22557, 16),
26588 => conv_std_logic_vector(22660, 16),
26589 => conv_std_logic_vector(22763, 16),
26590 => conv_std_logic_vector(22866, 16),
26591 => conv_std_logic_vector(22969, 16),
26592 => conv_std_logic_vector(23072, 16),
26593 => conv_std_logic_vector(23175, 16),
26594 => conv_std_logic_vector(23278, 16),
26595 => conv_std_logic_vector(23381, 16),
26596 => conv_std_logic_vector(23484, 16),
26597 => conv_std_logic_vector(23587, 16),
26598 => conv_std_logic_vector(23690, 16),
26599 => conv_std_logic_vector(23793, 16),
26600 => conv_std_logic_vector(23896, 16),
26601 => conv_std_logic_vector(23999, 16),
26602 => conv_std_logic_vector(24102, 16),
26603 => conv_std_logic_vector(24205, 16),
26604 => conv_std_logic_vector(24308, 16),
26605 => conv_std_logic_vector(24411, 16),
26606 => conv_std_logic_vector(24514, 16),
26607 => conv_std_logic_vector(24617, 16),
26608 => conv_std_logic_vector(24720, 16),
26609 => conv_std_logic_vector(24823, 16),
26610 => conv_std_logic_vector(24926, 16),
26611 => conv_std_logic_vector(25029, 16),
26612 => conv_std_logic_vector(25132, 16),
26613 => conv_std_logic_vector(25235, 16),
26614 => conv_std_logic_vector(25338, 16),
26615 => conv_std_logic_vector(25441, 16),
26616 => conv_std_logic_vector(25544, 16),
26617 => conv_std_logic_vector(25647, 16),
26618 => conv_std_logic_vector(25750, 16),
26619 => conv_std_logic_vector(25853, 16),
26620 => conv_std_logic_vector(25956, 16),
26621 => conv_std_logic_vector(26059, 16),
26622 => conv_std_logic_vector(26162, 16),
26623 => conv_std_logic_vector(26265, 16),
26624 => conv_std_logic_vector(0, 16),
26625 => conv_std_logic_vector(104, 16),
26626 => conv_std_logic_vector(208, 16),
26627 => conv_std_logic_vector(312, 16),
26628 => conv_std_logic_vector(416, 16),
26629 => conv_std_logic_vector(520, 16),
26630 => conv_std_logic_vector(624, 16),
26631 => conv_std_logic_vector(728, 16),
26632 => conv_std_logic_vector(832, 16),
26633 => conv_std_logic_vector(936, 16),
26634 => conv_std_logic_vector(1040, 16),
26635 => conv_std_logic_vector(1144, 16),
26636 => conv_std_logic_vector(1248, 16),
26637 => conv_std_logic_vector(1352, 16),
26638 => conv_std_logic_vector(1456, 16),
26639 => conv_std_logic_vector(1560, 16),
26640 => conv_std_logic_vector(1664, 16),
26641 => conv_std_logic_vector(1768, 16),
26642 => conv_std_logic_vector(1872, 16),
26643 => conv_std_logic_vector(1976, 16),
26644 => conv_std_logic_vector(2080, 16),
26645 => conv_std_logic_vector(2184, 16),
26646 => conv_std_logic_vector(2288, 16),
26647 => conv_std_logic_vector(2392, 16),
26648 => conv_std_logic_vector(2496, 16),
26649 => conv_std_logic_vector(2600, 16),
26650 => conv_std_logic_vector(2704, 16),
26651 => conv_std_logic_vector(2808, 16),
26652 => conv_std_logic_vector(2912, 16),
26653 => conv_std_logic_vector(3016, 16),
26654 => conv_std_logic_vector(3120, 16),
26655 => conv_std_logic_vector(3224, 16),
26656 => conv_std_logic_vector(3328, 16),
26657 => conv_std_logic_vector(3432, 16),
26658 => conv_std_logic_vector(3536, 16),
26659 => conv_std_logic_vector(3640, 16),
26660 => conv_std_logic_vector(3744, 16),
26661 => conv_std_logic_vector(3848, 16),
26662 => conv_std_logic_vector(3952, 16),
26663 => conv_std_logic_vector(4056, 16),
26664 => conv_std_logic_vector(4160, 16),
26665 => conv_std_logic_vector(4264, 16),
26666 => conv_std_logic_vector(4368, 16),
26667 => conv_std_logic_vector(4472, 16),
26668 => conv_std_logic_vector(4576, 16),
26669 => conv_std_logic_vector(4680, 16),
26670 => conv_std_logic_vector(4784, 16),
26671 => conv_std_logic_vector(4888, 16),
26672 => conv_std_logic_vector(4992, 16),
26673 => conv_std_logic_vector(5096, 16),
26674 => conv_std_logic_vector(5200, 16),
26675 => conv_std_logic_vector(5304, 16),
26676 => conv_std_logic_vector(5408, 16),
26677 => conv_std_logic_vector(5512, 16),
26678 => conv_std_logic_vector(5616, 16),
26679 => conv_std_logic_vector(5720, 16),
26680 => conv_std_logic_vector(5824, 16),
26681 => conv_std_logic_vector(5928, 16),
26682 => conv_std_logic_vector(6032, 16),
26683 => conv_std_logic_vector(6136, 16),
26684 => conv_std_logic_vector(6240, 16),
26685 => conv_std_logic_vector(6344, 16),
26686 => conv_std_logic_vector(6448, 16),
26687 => conv_std_logic_vector(6552, 16),
26688 => conv_std_logic_vector(6656, 16),
26689 => conv_std_logic_vector(6760, 16),
26690 => conv_std_logic_vector(6864, 16),
26691 => conv_std_logic_vector(6968, 16),
26692 => conv_std_logic_vector(7072, 16),
26693 => conv_std_logic_vector(7176, 16),
26694 => conv_std_logic_vector(7280, 16),
26695 => conv_std_logic_vector(7384, 16),
26696 => conv_std_logic_vector(7488, 16),
26697 => conv_std_logic_vector(7592, 16),
26698 => conv_std_logic_vector(7696, 16),
26699 => conv_std_logic_vector(7800, 16),
26700 => conv_std_logic_vector(7904, 16),
26701 => conv_std_logic_vector(8008, 16),
26702 => conv_std_logic_vector(8112, 16),
26703 => conv_std_logic_vector(8216, 16),
26704 => conv_std_logic_vector(8320, 16),
26705 => conv_std_logic_vector(8424, 16),
26706 => conv_std_logic_vector(8528, 16),
26707 => conv_std_logic_vector(8632, 16),
26708 => conv_std_logic_vector(8736, 16),
26709 => conv_std_logic_vector(8840, 16),
26710 => conv_std_logic_vector(8944, 16),
26711 => conv_std_logic_vector(9048, 16),
26712 => conv_std_logic_vector(9152, 16),
26713 => conv_std_logic_vector(9256, 16),
26714 => conv_std_logic_vector(9360, 16),
26715 => conv_std_logic_vector(9464, 16),
26716 => conv_std_logic_vector(9568, 16),
26717 => conv_std_logic_vector(9672, 16),
26718 => conv_std_logic_vector(9776, 16),
26719 => conv_std_logic_vector(9880, 16),
26720 => conv_std_logic_vector(9984, 16),
26721 => conv_std_logic_vector(10088, 16),
26722 => conv_std_logic_vector(10192, 16),
26723 => conv_std_logic_vector(10296, 16),
26724 => conv_std_logic_vector(10400, 16),
26725 => conv_std_logic_vector(10504, 16),
26726 => conv_std_logic_vector(10608, 16),
26727 => conv_std_logic_vector(10712, 16),
26728 => conv_std_logic_vector(10816, 16),
26729 => conv_std_logic_vector(10920, 16),
26730 => conv_std_logic_vector(11024, 16),
26731 => conv_std_logic_vector(11128, 16),
26732 => conv_std_logic_vector(11232, 16),
26733 => conv_std_logic_vector(11336, 16),
26734 => conv_std_logic_vector(11440, 16),
26735 => conv_std_logic_vector(11544, 16),
26736 => conv_std_logic_vector(11648, 16),
26737 => conv_std_logic_vector(11752, 16),
26738 => conv_std_logic_vector(11856, 16),
26739 => conv_std_logic_vector(11960, 16),
26740 => conv_std_logic_vector(12064, 16),
26741 => conv_std_logic_vector(12168, 16),
26742 => conv_std_logic_vector(12272, 16),
26743 => conv_std_logic_vector(12376, 16),
26744 => conv_std_logic_vector(12480, 16),
26745 => conv_std_logic_vector(12584, 16),
26746 => conv_std_logic_vector(12688, 16),
26747 => conv_std_logic_vector(12792, 16),
26748 => conv_std_logic_vector(12896, 16),
26749 => conv_std_logic_vector(13000, 16),
26750 => conv_std_logic_vector(13104, 16),
26751 => conv_std_logic_vector(13208, 16),
26752 => conv_std_logic_vector(13312, 16),
26753 => conv_std_logic_vector(13416, 16),
26754 => conv_std_logic_vector(13520, 16),
26755 => conv_std_logic_vector(13624, 16),
26756 => conv_std_logic_vector(13728, 16),
26757 => conv_std_logic_vector(13832, 16),
26758 => conv_std_logic_vector(13936, 16),
26759 => conv_std_logic_vector(14040, 16),
26760 => conv_std_logic_vector(14144, 16),
26761 => conv_std_logic_vector(14248, 16),
26762 => conv_std_logic_vector(14352, 16),
26763 => conv_std_logic_vector(14456, 16),
26764 => conv_std_logic_vector(14560, 16),
26765 => conv_std_logic_vector(14664, 16),
26766 => conv_std_logic_vector(14768, 16),
26767 => conv_std_logic_vector(14872, 16),
26768 => conv_std_logic_vector(14976, 16),
26769 => conv_std_logic_vector(15080, 16),
26770 => conv_std_logic_vector(15184, 16),
26771 => conv_std_logic_vector(15288, 16),
26772 => conv_std_logic_vector(15392, 16),
26773 => conv_std_logic_vector(15496, 16),
26774 => conv_std_logic_vector(15600, 16),
26775 => conv_std_logic_vector(15704, 16),
26776 => conv_std_logic_vector(15808, 16),
26777 => conv_std_logic_vector(15912, 16),
26778 => conv_std_logic_vector(16016, 16),
26779 => conv_std_logic_vector(16120, 16),
26780 => conv_std_logic_vector(16224, 16),
26781 => conv_std_logic_vector(16328, 16),
26782 => conv_std_logic_vector(16432, 16),
26783 => conv_std_logic_vector(16536, 16),
26784 => conv_std_logic_vector(16640, 16),
26785 => conv_std_logic_vector(16744, 16),
26786 => conv_std_logic_vector(16848, 16),
26787 => conv_std_logic_vector(16952, 16),
26788 => conv_std_logic_vector(17056, 16),
26789 => conv_std_logic_vector(17160, 16),
26790 => conv_std_logic_vector(17264, 16),
26791 => conv_std_logic_vector(17368, 16),
26792 => conv_std_logic_vector(17472, 16),
26793 => conv_std_logic_vector(17576, 16),
26794 => conv_std_logic_vector(17680, 16),
26795 => conv_std_logic_vector(17784, 16),
26796 => conv_std_logic_vector(17888, 16),
26797 => conv_std_logic_vector(17992, 16),
26798 => conv_std_logic_vector(18096, 16),
26799 => conv_std_logic_vector(18200, 16),
26800 => conv_std_logic_vector(18304, 16),
26801 => conv_std_logic_vector(18408, 16),
26802 => conv_std_logic_vector(18512, 16),
26803 => conv_std_logic_vector(18616, 16),
26804 => conv_std_logic_vector(18720, 16),
26805 => conv_std_logic_vector(18824, 16),
26806 => conv_std_logic_vector(18928, 16),
26807 => conv_std_logic_vector(19032, 16),
26808 => conv_std_logic_vector(19136, 16),
26809 => conv_std_logic_vector(19240, 16),
26810 => conv_std_logic_vector(19344, 16),
26811 => conv_std_logic_vector(19448, 16),
26812 => conv_std_logic_vector(19552, 16),
26813 => conv_std_logic_vector(19656, 16),
26814 => conv_std_logic_vector(19760, 16),
26815 => conv_std_logic_vector(19864, 16),
26816 => conv_std_logic_vector(19968, 16),
26817 => conv_std_logic_vector(20072, 16),
26818 => conv_std_logic_vector(20176, 16),
26819 => conv_std_logic_vector(20280, 16),
26820 => conv_std_logic_vector(20384, 16),
26821 => conv_std_logic_vector(20488, 16),
26822 => conv_std_logic_vector(20592, 16),
26823 => conv_std_logic_vector(20696, 16),
26824 => conv_std_logic_vector(20800, 16),
26825 => conv_std_logic_vector(20904, 16),
26826 => conv_std_logic_vector(21008, 16),
26827 => conv_std_logic_vector(21112, 16),
26828 => conv_std_logic_vector(21216, 16),
26829 => conv_std_logic_vector(21320, 16),
26830 => conv_std_logic_vector(21424, 16),
26831 => conv_std_logic_vector(21528, 16),
26832 => conv_std_logic_vector(21632, 16),
26833 => conv_std_logic_vector(21736, 16),
26834 => conv_std_logic_vector(21840, 16),
26835 => conv_std_logic_vector(21944, 16),
26836 => conv_std_logic_vector(22048, 16),
26837 => conv_std_logic_vector(22152, 16),
26838 => conv_std_logic_vector(22256, 16),
26839 => conv_std_logic_vector(22360, 16),
26840 => conv_std_logic_vector(22464, 16),
26841 => conv_std_logic_vector(22568, 16),
26842 => conv_std_logic_vector(22672, 16),
26843 => conv_std_logic_vector(22776, 16),
26844 => conv_std_logic_vector(22880, 16),
26845 => conv_std_logic_vector(22984, 16),
26846 => conv_std_logic_vector(23088, 16),
26847 => conv_std_logic_vector(23192, 16),
26848 => conv_std_logic_vector(23296, 16),
26849 => conv_std_logic_vector(23400, 16),
26850 => conv_std_logic_vector(23504, 16),
26851 => conv_std_logic_vector(23608, 16),
26852 => conv_std_logic_vector(23712, 16),
26853 => conv_std_logic_vector(23816, 16),
26854 => conv_std_logic_vector(23920, 16),
26855 => conv_std_logic_vector(24024, 16),
26856 => conv_std_logic_vector(24128, 16),
26857 => conv_std_logic_vector(24232, 16),
26858 => conv_std_logic_vector(24336, 16),
26859 => conv_std_logic_vector(24440, 16),
26860 => conv_std_logic_vector(24544, 16),
26861 => conv_std_logic_vector(24648, 16),
26862 => conv_std_logic_vector(24752, 16),
26863 => conv_std_logic_vector(24856, 16),
26864 => conv_std_logic_vector(24960, 16),
26865 => conv_std_logic_vector(25064, 16),
26866 => conv_std_logic_vector(25168, 16),
26867 => conv_std_logic_vector(25272, 16),
26868 => conv_std_logic_vector(25376, 16),
26869 => conv_std_logic_vector(25480, 16),
26870 => conv_std_logic_vector(25584, 16),
26871 => conv_std_logic_vector(25688, 16),
26872 => conv_std_logic_vector(25792, 16),
26873 => conv_std_logic_vector(25896, 16),
26874 => conv_std_logic_vector(26000, 16),
26875 => conv_std_logic_vector(26104, 16),
26876 => conv_std_logic_vector(26208, 16),
26877 => conv_std_logic_vector(26312, 16),
26878 => conv_std_logic_vector(26416, 16),
26879 => conv_std_logic_vector(26520, 16),
26880 => conv_std_logic_vector(0, 16),
26881 => conv_std_logic_vector(105, 16),
26882 => conv_std_logic_vector(210, 16),
26883 => conv_std_logic_vector(315, 16),
26884 => conv_std_logic_vector(420, 16),
26885 => conv_std_logic_vector(525, 16),
26886 => conv_std_logic_vector(630, 16),
26887 => conv_std_logic_vector(735, 16),
26888 => conv_std_logic_vector(840, 16),
26889 => conv_std_logic_vector(945, 16),
26890 => conv_std_logic_vector(1050, 16),
26891 => conv_std_logic_vector(1155, 16),
26892 => conv_std_logic_vector(1260, 16),
26893 => conv_std_logic_vector(1365, 16),
26894 => conv_std_logic_vector(1470, 16),
26895 => conv_std_logic_vector(1575, 16),
26896 => conv_std_logic_vector(1680, 16),
26897 => conv_std_logic_vector(1785, 16),
26898 => conv_std_logic_vector(1890, 16),
26899 => conv_std_logic_vector(1995, 16),
26900 => conv_std_logic_vector(2100, 16),
26901 => conv_std_logic_vector(2205, 16),
26902 => conv_std_logic_vector(2310, 16),
26903 => conv_std_logic_vector(2415, 16),
26904 => conv_std_logic_vector(2520, 16),
26905 => conv_std_logic_vector(2625, 16),
26906 => conv_std_logic_vector(2730, 16),
26907 => conv_std_logic_vector(2835, 16),
26908 => conv_std_logic_vector(2940, 16),
26909 => conv_std_logic_vector(3045, 16),
26910 => conv_std_logic_vector(3150, 16),
26911 => conv_std_logic_vector(3255, 16),
26912 => conv_std_logic_vector(3360, 16),
26913 => conv_std_logic_vector(3465, 16),
26914 => conv_std_logic_vector(3570, 16),
26915 => conv_std_logic_vector(3675, 16),
26916 => conv_std_logic_vector(3780, 16),
26917 => conv_std_logic_vector(3885, 16),
26918 => conv_std_logic_vector(3990, 16),
26919 => conv_std_logic_vector(4095, 16),
26920 => conv_std_logic_vector(4200, 16),
26921 => conv_std_logic_vector(4305, 16),
26922 => conv_std_logic_vector(4410, 16),
26923 => conv_std_logic_vector(4515, 16),
26924 => conv_std_logic_vector(4620, 16),
26925 => conv_std_logic_vector(4725, 16),
26926 => conv_std_logic_vector(4830, 16),
26927 => conv_std_logic_vector(4935, 16),
26928 => conv_std_logic_vector(5040, 16),
26929 => conv_std_logic_vector(5145, 16),
26930 => conv_std_logic_vector(5250, 16),
26931 => conv_std_logic_vector(5355, 16),
26932 => conv_std_logic_vector(5460, 16),
26933 => conv_std_logic_vector(5565, 16),
26934 => conv_std_logic_vector(5670, 16),
26935 => conv_std_logic_vector(5775, 16),
26936 => conv_std_logic_vector(5880, 16),
26937 => conv_std_logic_vector(5985, 16),
26938 => conv_std_logic_vector(6090, 16),
26939 => conv_std_logic_vector(6195, 16),
26940 => conv_std_logic_vector(6300, 16),
26941 => conv_std_logic_vector(6405, 16),
26942 => conv_std_logic_vector(6510, 16),
26943 => conv_std_logic_vector(6615, 16),
26944 => conv_std_logic_vector(6720, 16),
26945 => conv_std_logic_vector(6825, 16),
26946 => conv_std_logic_vector(6930, 16),
26947 => conv_std_logic_vector(7035, 16),
26948 => conv_std_logic_vector(7140, 16),
26949 => conv_std_logic_vector(7245, 16),
26950 => conv_std_logic_vector(7350, 16),
26951 => conv_std_logic_vector(7455, 16),
26952 => conv_std_logic_vector(7560, 16),
26953 => conv_std_logic_vector(7665, 16),
26954 => conv_std_logic_vector(7770, 16),
26955 => conv_std_logic_vector(7875, 16),
26956 => conv_std_logic_vector(7980, 16),
26957 => conv_std_logic_vector(8085, 16),
26958 => conv_std_logic_vector(8190, 16),
26959 => conv_std_logic_vector(8295, 16),
26960 => conv_std_logic_vector(8400, 16),
26961 => conv_std_logic_vector(8505, 16),
26962 => conv_std_logic_vector(8610, 16),
26963 => conv_std_logic_vector(8715, 16),
26964 => conv_std_logic_vector(8820, 16),
26965 => conv_std_logic_vector(8925, 16),
26966 => conv_std_logic_vector(9030, 16),
26967 => conv_std_logic_vector(9135, 16),
26968 => conv_std_logic_vector(9240, 16),
26969 => conv_std_logic_vector(9345, 16),
26970 => conv_std_logic_vector(9450, 16),
26971 => conv_std_logic_vector(9555, 16),
26972 => conv_std_logic_vector(9660, 16),
26973 => conv_std_logic_vector(9765, 16),
26974 => conv_std_logic_vector(9870, 16),
26975 => conv_std_logic_vector(9975, 16),
26976 => conv_std_logic_vector(10080, 16),
26977 => conv_std_logic_vector(10185, 16),
26978 => conv_std_logic_vector(10290, 16),
26979 => conv_std_logic_vector(10395, 16),
26980 => conv_std_logic_vector(10500, 16),
26981 => conv_std_logic_vector(10605, 16),
26982 => conv_std_logic_vector(10710, 16),
26983 => conv_std_logic_vector(10815, 16),
26984 => conv_std_logic_vector(10920, 16),
26985 => conv_std_logic_vector(11025, 16),
26986 => conv_std_logic_vector(11130, 16),
26987 => conv_std_logic_vector(11235, 16),
26988 => conv_std_logic_vector(11340, 16),
26989 => conv_std_logic_vector(11445, 16),
26990 => conv_std_logic_vector(11550, 16),
26991 => conv_std_logic_vector(11655, 16),
26992 => conv_std_logic_vector(11760, 16),
26993 => conv_std_logic_vector(11865, 16),
26994 => conv_std_logic_vector(11970, 16),
26995 => conv_std_logic_vector(12075, 16),
26996 => conv_std_logic_vector(12180, 16),
26997 => conv_std_logic_vector(12285, 16),
26998 => conv_std_logic_vector(12390, 16),
26999 => conv_std_logic_vector(12495, 16),
27000 => conv_std_logic_vector(12600, 16),
27001 => conv_std_logic_vector(12705, 16),
27002 => conv_std_logic_vector(12810, 16),
27003 => conv_std_logic_vector(12915, 16),
27004 => conv_std_logic_vector(13020, 16),
27005 => conv_std_logic_vector(13125, 16),
27006 => conv_std_logic_vector(13230, 16),
27007 => conv_std_logic_vector(13335, 16),
27008 => conv_std_logic_vector(13440, 16),
27009 => conv_std_logic_vector(13545, 16),
27010 => conv_std_logic_vector(13650, 16),
27011 => conv_std_logic_vector(13755, 16),
27012 => conv_std_logic_vector(13860, 16),
27013 => conv_std_logic_vector(13965, 16),
27014 => conv_std_logic_vector(14070, 16),
27015 => conv_std_logic_vector(14175, 16),
27016 => conv_std_logic_vector(14280, 16),
27017 => conv_std_logic_vector(14385, 16),
27018 => conv_std_logic_vector(14490, 16),
27019 => conv_std_logic_vector(14595, 16),
27020 => conv_std_logic_vector(14700, 16),
27021 => conv_std_logic_vector(14805, 16),
27022 => conv_std_logic_vector(14910, 16),
27023 => conv_std_logic_vector(15015, 16),
27024 => conv_std_logic_vector(15120, 16),
27025 => conv_std_logic_vector(15225, 16),
27026 => conv_std_logic_vector(15330, 16),
27027 => conv_std_logic_vector(15435, 16),
27028 => conv_std_logic_vector(15540, 16),
27029 => conv_std_logic_vector(15645, 16),
27030 => conv_std_logic_vector(15750, 16),
27031 => conv_std_logic_vector(15855, 16),
27032 => conv_std_logic_vector(15960, 16),
27033 => conv_std_logic_vector(16065, 16),
27034 => conv_std_logic_vector(16170, 16),
27035 => conv_std_logic_vector(16275, 16),
27036 => conv_std_logic_vector(16380, 16),
27037 => conv_std_logic_vector(16485, 16),
27038 => conv_std_logic_vector(16590, 16),
27039 => conv_std_logic_vector(16695, 16),
27040 => conv_std_logic_vector(16800, 16),
27041 => conv_std_logic_vector(16905, 16),
27042 => conv_std_logic_vector(17010, 16),
27043 => conv_std_logic_vector(17115, 16),
27044 => conv_std_logic_vector(17220, 16),
27045 => conv_std_logic_vector(17325, 16),
27046 => conv_std_logic_vector(17430, 16),
27047 => conv_std_logic_vector(17535, 16),
27048 => conv_std_logic_vector(17640, 16),
27049 => conv_std_logic_vector(17745, 16),
27050 => conv_std_logic_vector(17850, 16),
27051 => conv_std_logic_vector(17955, 16),
27052 => conv_std_logic_vector(18060, 16),
27053 => conv_std_logic_vector(18165, 16),
27054 => conv_std_logic_vector(18270, 16),
27055 => conv_std_logic_vector(18375, 16),
27056 => conv_std_logic_vector(18480, 16),
27057 => conv_std_logic_vector(18585, 16),
27058 => conv_std_logic_vector(18690, 16),
27059 => conv_std_logic_vector(18795, 16),
27060 => conv_std_logic_vector(18900, 16),
27061 => conv_std_logic_vector(19005, 16),
27062 => conv_std_logic_vector(19110, 16),
27063 => conv_std_logic_vector(19215, 16),
27064 => conv_std_logic_vector(19320, 16),
27065 => conv_std_logic_vector(19425, 16),
27066 => conv_std_logic_vector(19530, 16),
27067 => conv_std_logic_vector(19635, 16),
27068 => conv_std_logic_vector(19740, 16),
27069 => conv_std_logic_vector(19845, 16),
27070 => conv_std_logic_vector(19950, 16),
27071 => conv_std_logic_vector(20055, 16),
27072 => conv_std_logic_vector(20160, 16),
27073 => conv_std_logic_vector(20265, 16),
27074 => conv_std_logic_vector(20370, 16),
27075 => conv_std_logic_vector(20475, 16),
27076 => conv_std_logic_vector(20580, 16),
27077 => conv_std_logic_vector(20685, 16),
27078 => conv_std_logic_vector(20790, 16),
27079 => conv_std_logic_vector(20895, 16),
27080 => conv_std_logic_vector(21000, 16),
27081 => conv_std_logic_vector(21105, 16),
27082 => conv_std_logic_vector(21210, 16),
27083 => conv_std_logic_vector(21315, 16),
27084 => conv_std_logic_vector(21420, 16),
27085 => conv_std_logic_vector(21525, 16),
27086 => conv_std_logic_vector(21630, 16),
27087 => conv_std_logic_vector(21735, 16),
27088 => conv_std_logic_vector(21840, 16),
27089 => conv_std_logic_vector(21945, 16),
27090 => conv_std_logic_vector(22050, 16),
27091 => conv_std_logic_vector(22155, 16),
27092 => conv_std_logic_vector(22260, 16),
27093 => conv_std_logic_vector(22365, 16),
27094 => conv_std_logic_vector(22470, 16),
27095 => conv_std_logic_vector(22575, 16),
27096 => conv_std_logic_vector(22680, 16),
27097 => conv_std_logic_vector(22785, 16),
27098 => conv_std_logic_vector(22890, 16),
27099 => conv_std_logic_vector(22995, 16),
27100 => conv_std_logic_vector(23100, 16),
27101 => conv_std_logic_vector(23205, 16),
27102 => conv_std_logic_vector(23310, 16),
27103 => conv_std_logic_vector(23415, 16),
27104 => conv_std_logic_vector(23520, 16),
27105 => conv_std_logic_vector(23625, 16),
27106 => conv_std_logic_vector(23730, 16),
27107 => conv_std_logic_vector(23835, 16),
27108 => conv_std_logic_vector(23940, 16),
27109 => conv_std_logic_vector(24045, 16),
27110 => conv_std_logic_vector(24150, 16),
27111 => conv_std_logic_vector(24255, 16),
27112 => conv_std_logic_vector(24360, 16),
27113 => conv_std_logic_vector(24465, 16),
27114 => conv_std_logic_vector(24570, 16),
27115 => conv_std_logic_vector(24675, 16),
27116 => conv_std_logic_vector(24780, 16),
27117 => conv_std_logic_vector(24885, 16),
27118 => conv_std_logic_vector(24990, 16),
27119 => conv_std_logic_vector(25095, 16),
27120 => conv_std_logic_vector(25200, 16),
27121 => conv_std_logic_vector(25305, 16),
27122 => conv_std_logic_vector(25410, 16),
27123 => conv_std_logic_vector(25515, 16),
27124 => conv_std_logic_vector(25620, 16),
27125 => conv_std_logic_vector(25725, 16),
27126 => conv_std_logic_vector(25830, 16),
27127 => conv_std_logic_vector(25935, 16),
27128 => conv_std_logic_vector(26040, 16),
27129 => conv_std_logic_vector(26145, 16),
27130 => conv_std_logic_vector(26250, 16),
27131 => conv_std_logic_vector(26355, 16),
27132 => conv_std_logic_vector(26460, 16),
27133 => conv_std_logic_vector(26565, 16),
27134 => conv_std_logic_vector(26670, 16),
27135 => conv_std_logic_vector(26775, 16),
27136 => conv_std_logic_vector(0, 16),
27137 => conv_std_logic_vector(106, 16),
27138 => conv_std_logic_vector(212, 16),
27139 => conv_std_logic_vector(318, 16),
27140 => conv_std_logic_vector(424, 16),
27141 => conv_std_logic_vector(530, 16),
27142 => conv_std_logic_vector(636, 16),
27143 => conv_std_logic_vector(742, 16),
27144 => conv_std_logic_vector(848, 16),
27145 => conv_std_logic_vector(954, 16),
27146 => conv_std_logic_vector(1060, 16),
27147 => conv_std_logic_vector(1166, 16),
27148 => conv_std_logic_vector(1272, 16),
27149 => conv_std_logic_vector(1378, 16),
27150 => conv_std_logic_vector(1484, 16),
27151 => conv_std_logic_vector(1590, 16),
27152 => conv_std_logic_vector(1696, 16),
27153 => conv_std_logic_vector(1802, 16),
27154 => conv_std_logic_vector(1908, 16),
27155 => conv_std_logic_vector(2014, 16),
27156 => conv_std_logic_vector(2120, 16),
27157 => conv_std_logic_vector(2226, 16),
27158 => conv_std_logic_vector(2332, 16),
27159 => conv_std_logic_vector(2438, 16),
27160 => conv_std_logic_vector(2544, 16),
27161 => conv_std_logic_vector(2650, 16),
27162 => conv_std_logic_vector(2756, 16),
27163 => conv_std_logic_vector(2862, 16),
27164 => conv_std_logic_vector(2968, 16),
27165 => conv_std_logic_vector(3074, 16),
27166 => conv_std_logic_vector(3180, 16),
27167 => conv_std_logic_vector(3286, 16),
27168 => conv_std_logic_vector(3392, 16),
27169 => conv_std_logic_vector(3498, 16),
27170 => conv_std_logic_vector(3604, 16),
27171 => conv_std_logic_vector(3710, 16),
27172 => conv_std_logic_vector(3816, 16),
27173 => conv_std_logic_vector(3922, 16),
27174 => conv_std_logic_vector(4028, 16),
27175 => conv_std_logic_vector(4134, 16),
27176 => conv_std_logic_vector(4240, 16),
27177 => conv_std_logic_vector(4346, 16),
27178 => conv_std_logic_vector(4452, 16),
27179 => conv_std_logic_vector(4558, 16),
27180 => conv_std_logic_vector(4664, 16),
27181 => conv_std_logic_vector(4770, 16),
27182 => conv_std_logic_vector(4876, 16),
27183 => conv_std_logic_vector(4982, 16),
27184 => conv_std_logic_vector(5088, 16),
27185 => conv_std_logic_vector(5194, 16),
27186 => conv_std_logic_vector(5300, 16),
27187 => conv_std_logic_vector(5406, 16),
27188 => conv_std_logic_vector(5512, 16),
27189 => conv_std_logic_vector(5618, 16),
27190 => conv_std_logic_vector(5724, 16),
27191 => conv_std_logic_vector(5830, 16),
27192 => conv_std_logic_vector(5936, 16),
27193 => conv_std_logic_vector(6042, 16),
27194 => conv_std_logic_vector(6148, 16),
27195 => conv_std_logic_vector(6254, 16),
27196 => conv_std_logic_vector(6360, 16),
27197 => conv_std_logic_vector(6466, 16),
27198 => conv_std_logic_vector(6572, 16),
27199 => conv_std_logic_vector(6678, 16),
27200 => conv_std_logic_vector(6784, 16),
27201 => conv_std_logic_vector(6890, 16),
27202 => conv_std_logic_vector(6996, 16),
27203 => conv_std_logic_vector(7102, 16),
27204 => conv_std_logic_vector(7208, 16),
27205 => conv_std_logic_vector(7314, 16),
27206 => conv_std_logic_vector(7420, 16),
27207 => conv_std_logic_vector(7526, 16),
27208 => conv_std_logic_vector(7632, 16),
27209 => conv_std_logic_vector(7738, 16),
27210 => conv_std_logic_vector(7844, 16),
27211 => conv_std_logic_vector(7950, 16),
27212 => conv_std_logic_vector(8056, 16),
27213 => conv_std_logic_vector(8162, 16),
27214 => conv_std_logic_vector(8268, 16),
27215 => conv_std_logic_vector(8374, 16),
27216 => conv_std_logic_vector(8480, 16),
27217 => conv_std_logic_vector(8586, 16),
27218 => conv_std_logic_vector(8692, 16),
27219 => conv_std_logic_vector(8798, 16),
27220 => conv_std_logic_vector(8904, 16),
27221 => conv_std_logic_vector(9010, 16),
27222 => conv_std_logic_vector(9116, 16),
27223 => conv_std_logic_vector(9222, 16),
27224 => conv_std_logic_vector(9328, 16),
27225 => conv_std_logic_vector(9434, 16),
27226 => conv_std_logic_vector(9540, 16),
27227 => conv_std_logic_vector(9646, 16),
27228 => conv_std_logic_vector(9752, 16),
27229 => conv_std_logic_vector(9858, 16),
27230 => conv_std_logic_vector(9964, 16),
27231 => conv_std_logic_vector(10070, 16),
27232 => conv_std_logic_vector(10176, 16),
27233 => conv_std_logic_vector(10282, 16),
27234 => conv_std_logic_vector(10388, 16),
27235 => conv_std_logic_vector(10494, 16),
27236 => conv_std_logic_vector(10600, 16),
27237 => conv_std_logic_vector(10706, 16),
27238 => conv_std_logic_vector(10812, 16),
27239 => conv_std_logic_vector(10918, 16),
27240 => conv_std_logic_vector(11024, 16),
27241 => conv_std_logic_vector(11130, 16),
27242 => conv_std_logic_vector(11236, 16),
27243 => conv_std_logic_vector(11342, 16),
27244 => conv_std_logic_vector(11448, 16),
27245 => conv_std_logic_vector(11554, 16),
27246 => conv_std_logic_vector(11660, 16),
27247 => conv_std_logic_vector(11766, 16),
27248 => conv_std_logic_vector(11872, 16),
27249 => conv_std_logic_vector(11978, 16),
27250 => conv_std_logic_vector(12084, 16),
27251 => conv_std_logic_vector(12190, 16),
27252 => conv_std_logic_vector(12296, 16),
27253 => conv_std_logic_vector(12402, 16),
27254 => conv_std_logic_vector(12508, 16),
27255 => conv_std_logic_vector(12614, 16),
27256 => conv_std_logic_vector(12720, 16),
27257 => conv_std_logic_vector(12826, 16),
27258 => conv_std_logic_vector(12932, 16),
27259 => conv_std_logic_vector(13038, 16),
27260 => conv_std_logic_vector(13144, 16),
27261 => conv_std_logic_vector(13250, 16),
27262 => conv_std_logic_vector(13356, 16),
27263 => conv_std_logic_vector(13462, 16),
27264 => conv_std_logic_vector(13568, 16),
27265 => conv_std_logic_vector(13674, 16),
27266 => conv_std_logic_vector(13780, 16),
27267 => conv_std_logic_vector(13886, 16),
27268 => conv_std_logic_vector(13992, 16),
27269 => conv_std_logic_vector(14098, 16),
27270 => conv_std_logic_vector(14204, 16),
27271 => conv_std_logic_vector(14310, 16),
27272 => conv_std_logic_vector(14416, 16),
27273 => conv_std_logic_vector(14522, 16),
27274 => conv_std_logic_vector(14628, 16),
27275 => conv_std_logic_vector(14734, 16),
27276 => conv_std_logic_vector(14840, 16),
27277 => conv_std_logic_vector(14946, 16),
27278 => conv_std_logic_vector(15052, 16),
27279 => conv_std_logic_vector(15158, 16),
27280 => conv_std_logic_vector(15264, 16),
27281 => conv_std_logic_vector(15370, 16),
27282 => conv_std_logic_vector(15476, 16),
27283 => conv_std_logic_vector(15582, 16),
27284 => conv_std_logic_vector(15688, 16),
27285 => conv_std_logic_vector(15794, 16),
27286 => conv_std_logic_vector(15900, 16),
27287 => conv_std_logic_vector(16006, 16),
27288 => conv_std_logic_vector(16112, 16),
27289 => conv_std_logic_vector(16218, 16),
27290 => conv_std_logic_vector(16324, 16),
27291 => conv_std_logic_vector(16430, 16),
27292 => conv_std_logic_vector(16536, 16),
27293 => conv_std_logic_vector(16642, 16),
27294 => conv_std_logic_vector(16748, 16),
27295 => conv_std_logic_vector(16854, 16),
27296 => conv_std_logic_vector(16960, 16),
27297 => conv_std_logic_vector(17066, 16),
27298 => conv_std_logic_vector(17172, 16),
27299 => conv_std_logic_vector(17278, 16),
27300 => conv_std_logic_vector(17384, 16),
27301 => conv_std_logic_vector(17490, 16),
27302 => conv_std_logic_vector(17596, 16),
27303 => conv_std_logic_vector(17702, 16),
27304 => conv_std_logic_vector(17808, 16),
27305 => conv_std_logic_vector(17914, 16),
27306 => conv_std_logic_vector(18020, 16),
27307 => conv_std_logic_vector(18126, 16),
27308 => conv_std_logic_vector(18232, 16),
27309 => conv_std_logic_vector(18338, 16),
27310 => conv_std_logic_vector(18444, 16),
27311 => conv_std_logic_vector(18550, 16),
27312 => conv_std_logic_vector(18656, 16),
27313 => conv_std_logic_vector(18762, 16),
27314 => conv_std_logic_vector(18868, 16),
27315 => conv_std_logic_vector(18974, 16),
27316 => conv_std_logic_vector(19080, 16),
27317 => conv_std_logic_vector(19186, 16),
27318 => conv_std_logic_vector(19292, 16),
27319 => conv_std_logic_vector(19398, 16),
27320 => conv_std_logic_vector(19504, 16),
27321 => conv_std_logic_vector(19610, 16),
27322 => conv_std_logic_vector(19716, 16),
27323 => conv_std_logic_vector(19822, 16),
27324 => conv_std_logic_vector(19928, 16),
27325 => conv_std_logic_vector(20034, 16),
27326 => conv_std_logic_vector(20140, 16),
27327 => conv_std_logic_vector(20246, 16),
27328 => conv_std_logic_vector(20352, 16),
27329 => conv_std_logic_vector(20458, 16),
27330 => conv_std_logic_vector(20564, 16),
27331 => conv_std_logic_vector(20670, 16),
27332 => conv_std_logic_vector(20776, 16),
27333 => conv_std_logic_vector(20882, 16),
27334 => conv_std_logic_vector(20988, 16),
27335 => conv_std_logic_vector(21094, 16),
27336 => conv_std_logic_vector(21200, 16),
27337 => conv_std_logic_vector(21306, 16),
27338 => conv_std_logic_vector(21412, 16),
27339 => conv_std_logic_vector(21518, 16),
27340 => conv_std_logic_vector(21624, 16),
27341 => conv_std_logic_vector(21730, 16),
27342 => conv_std_logic_vector(21836, 16),
27343 => conv_std_logic_vector(21942, 16),
27344 => conv_std_logic_vector(22048, 16),
27345 => conv_std_logic_vector(22154, 16),
27346 => conv_std_logic_vector(22260, 16),
27347 => conv_std_logic_vector(22366, 16),
27348 => conv_std_logic_vector(22472, 16),
27349 => conv_std_logic_vector(22578, 16),
27350 => conv_std_logic_vector(22684, 16),
27351 => conv_std_logic_vector(22790, 16),
27352 => conv_std_logic_vector(22896, 16),
27353 => conv_std_logic_vector(23002, 16),
27354 => conv_std_logic_vector(23108, 16),
27355 => conv_std_logic_vector(23214, 16),
27356 => conv_std_logic_vector(23320, 16),
27357 => conv_std_logic_vector(23426, 16),
27358 => conv_std_logic_vector(23532, 16),
27359 => conv_std_logic_vector(23638, 16),
27360 => conv_std_logic_vector(23744, 16),
27361 => conv_std_logic_vector(23850, 16),
27362 => conv_std_logic_vector(23956, 16),
27363 => conv_std_logic_vector(24062, 16),
27364 => conv_std_logic_vector(24168, 16),
27365 => conv_std_logic_vector(24274, 16),
27366 => conv_std_logic_vector(24380, 16),
27367 => conv_std_logic_vector(24486, 16),
27368 => conv_std_logic_vector(24592, 16),
27369 => conv_std_logic_vector(24698, 16),
27370 => conv_std_logic_vector(24804, 16),
27371 => conv_std_logic_vector(24910, 16),
27372 => conv_std_logic_vector(25016, 16),
27373 => conv_std_logic_vector(25122, 16),
27374 => conv_std_logic_vector(25228, 16),
27375 => conv_std_logic_vector(25334, 16),
27376 => conv_std_logic_vector(25440, 16),
27377 => conv_std_logic_vector(25546, 16),
27378 => conv_std_logic_vector(25652, 16),
27379 => conv_std_logic_vector(25758, 16),
27380 => conv_std_logic_vector(25864, 16),
27381 => conv_std_logic_vector(25970, 16),
27382 => conv_std_logic_vector(26076, 16),
27383 => conv_std_logic_vector(26182, 16),
27384 => conv_std_logic_vector(26288, 16),
27385 => conv_std_logic_vector(26394, 16),
27386 => conv_std_logic_vector(26500, 16),
27387 => conv_std_logic_vector(26606, 16),
27388 => conv_std_logic_vector(26712, 16),
27389 => conv_std_logic_vector(26818, 16),
27390 => conv_std_logic_vector(26924, 16),
27391 => conv_std_logic_vector(27030, 16),
27392 => conv_std_logic_vector(0, 16),
27393 => conv_std_logic_vector(107, 16),
27394 => conv_std_logic_vector(214, 16),
27395 => conv_std_logic_vector(321, 16),
27396 => conv_std_logic_vector(428, 16),
27397 => conv_std_logic_vector(535, 16),
27398 => conv_std_logic_vector(642, 16),
27399 => conv_std_logic_vector(749, 16),
27400 => conv_std_logic_vector(856, 16),
27401 => conv_std_logic_vector(963, 16),
27402 => conv_std_logic_vector(1070, 16),
27403 => conv_std_logic_vector(1177, 16),
27404 => conv_std_logic_vector(1284, 16),
27405 => conv_std_logic_vector(1391, 16),
27406 => conv_std_logic_vector(1498, 16),
27407 => conv_std_logic_vector(1605, 16),
27408 => conv_std_logic_vector(1712, 16),
27409 => conv_std_logic_vector(1819, 16),
27410 => conv_std_logic_vector(1926, 16),
27411 => conv_std_logic_vector(2033, 16),
27412 => conv_std_logic_vector(2140, 16),
27413 => conv_std_logic_vector(2247, 16),
27414 => conv_std_logic_vector(2354, 16),
27415 => conv_std_logic_vector(2461, 16),
27416 => conv_std_logic_vector(2568, 16),
27417 => conv_std_logic_vector(2675, 16),
27418 => conv_std_logic_vector(2782, 16),
27419 => conv_std_logic_vector(2889, 16),
27420 => conv_std_logic_vector(2996, 16),
27421 => conv_std_logic_vector(3103, 16),
27422 => conv_std_logic_vector(3210, 16),
27423 => conv_std_logic_vector(3317, 16),
27424 => conv_std_logic_vector(3424, 16),
27425 => conv_std_logic_vector(3531, 16),
27426 => conv_std_logic_vector(3638, 16),
27427 => conv_std_logic_vector(3745, 16),
27428 => conv_std_logic_vector(3852, 16),
27429 => conv_std_logic_vector(3959, 16),
27430 => conv_std_logic_vector(4066, 16),
27431 => conv_std_logic_vector(4173, 16),
27432 => conv_std_logic_vector(4280, 16),
27433 => conv_std_logic_vector(4387, 16),
27434 => conv_std_logic_vector(4494, 16),
27435 => conv_std_logic_vector(4601, 16),
27436 => conv_std_logic_vector(4708, 16),
27437 => conv_std_logic_vector(4815, 16),
27438 => conv_std_logic_vector(4922, 16),
27439 => conv_std_logic_vector(5029, 16),
27440 => conv_std_logic_vector(5136, 16),
27441 => conv_std_logic_vector(5243, 16),
27442 => conv_std_logic_vector(5350, 16),
27443 => conv_std_logic_vector(5457, 16),
27444 => conv_std_logic_vector(5564, 16),
27445 => conv_std_logic_vector(5671, 16),
27446 => conv_std_logic_vector(5778, 16),
27447 => conv_std_logic_vector(5885, 16),
27448 => conv_std_logic_vector(5992, 16),
27449 => conv_std_logic_vector(6099, 16),
27450 => conv_std_logic_vector(6206, 16),
27451 => conv_std_logic_vector(6313, 16),
27452 => conv_std_logic_vector(6420, 16),
27453 => conv_std_logic_vector(6527, 16),
27454 => conv_std_logic_vector(6634, 16),
27455 => conv_std_logic_vector(6741, 16),
27456 => conv_std_logic_vector(6848, 16),
27457 => conv_std_logic_vector(6955, 16),
27458 => conv_std_logic_vector(7062, 16),
27459 => conv_std_logic_vector(7169, 16),
27460 => conv_std_logic_vector(7276, 16),
27461 => conv_std_logic_vector(7383, 16),
27462 => conv_std_logic_vector(7490, 16),
27463 => conv_std_logic_vector(7597, 16),
27464 => conv_std_logic_vector(7704, 16),
27465 => conv_std_logic_vector(7811, 16),
27466 => conv_std_logic_vector(7918, 16),
27467 => conv_std_logic_vector(8025, 16),
27468 => conv_std_logic_vector(8132, 16),
27469 => conv_std_logic_vector(8239, 16),
27470 => conv_std_logic_vector(8346, 16),
27471 => conv_std_logic_vector(8453, 16),
27472 => conv_std_logic_vector(8560, 16),
27473 => conv_std_logic_vector(8667, 16),
27474 => conv_std_logic_vector(8774, 16),
27475 => conv_std_logic_vector(8881, 16),
27476 => conv_std_logic_vector(8988, 16),
27477 => conv_std_logic_vector(9095, 16),
27478 => conv_std_logic_vector(9202, 16),
27479 => conv_std_logic_vector(9309, 16),
27480 => conv_std_logic_vector(9416, 16),
27481 => conv_std_logic_vector(9523, 16),
27482 => conv_std_logic_vector(9630, 16),
27483 => conv_std_logic_vector(9737, 16),
27484 => conv_std_logic_vector(9844, 16),
27485 => conv_std_logic_vector(9951, 16),
27486 => conv_std_logic_vector(10058, 16),
27487 => conv_std_logic_vector(10165, 16),
27488 => conv_std_logic_vector(10272, 16),
27489 => conv_std_logic_vector(10379, 16),
27490 => conv_std_logic_vector(10486, 16),
27491 => conv_std_logic_vector(10593, 16),
27492 => conv_std_logic_vector(10700, 16),
27493 => conv_std_logic_vector(10807, 16),
27494 => conv_std_logic_vector(10914, 16),
27495 => conv_std_logic_vector(11021, 16),
27496 => conv_std_logic_vector(11128, 16),
27497 => conv_std_logic_vector(11235, 16),
27498 => conv_std_logic_vector(11342, 16),
27499 => conv_std_logic_vector(11449, 16),
27500 => conv_std_logic_vector(11556, 16),
27501 => conv_std_logic_vector(11663, 16),
27502 => conv_std_logic_vector(11770, 16),
27503 => conv_std_logic_vector(11877, 16),
27504 => conv_std_logic_vector(11984, 16),
27505 => conv_std_logic_vector(12091, 16),
27506 => conv_std_logic_vector(12198, 16),
27507 => conv_std_logic_vector(12305, 16),
27508 => conv_std_logic_vector(12412, 16),
27509 => conv_std_logic_vector(12519, 16),
27510 => conv_std_logic_vector(12626, 16),
27511 => conv_std_logic_vector(12733, 16),
27512 => conv_std_logic_vector(12840, 16),
27513 => conv_std_logic_vector(12947, 16),
27514 => conv_std_logic_vector(13054, 16),
27515 => conv_std_logic_vector(13161, 16),
27516 => conv_std_logic_vector(13268, 16),
27517 => conv_std_logic_vector(13375, 16),
27518 => conv_std_logic_vector(13482, 16),
27519 => conv_std_logic_vector(13589, 16),
27520 => conv_std_logic_vector(13696, 16),
27521 => conv_std_logic_vector(13803, 16),
27522 => conv_std_logic_vector(13910, 16),
27523 => conv_std_logic_vector(14017, 16),
27524 => conv_std_logic_vector(14124, 16),
27525 => conv_std_logic_vector(14231, 16),
27526 => conv_std_logic_vector(14338, 16),
27527 => conv_std_logic_vector(14445, 16),
27528 => conv_std_logic_vector(14552, 16),
27529 => conv_std_logic_vector(14659, 16),
27530 => conv_std_logic_vector(14766, 16),
27531 => conv_std_logic_vector(14873, 16),
27532 => conv_std_logic_vector(14980, 16),
27533 => conv_std_logic_vector(15087, 16),
27534 => conv_std_logic_vector(15194, 16),
27535 => conv_std_logic_vector(15301, 16),
27536 => conv_std_logic_vector(15408, 16),
27537 => conv_std_logic_vector(15515, 16),
27538 => conv_std_logic_vector(15622, 16),
27539 => conv_std_logic_vector(15729, 16),
27540 => conv_std_logic_vector(15836, 16),
27541 => conv_std_logic_vector(15943, 16),
27542 => conv_std_logic_vector(16050, 16),
27543 => conv_std_logic_vector(16157, 16),
27544 => conv_std_logic_vector(16264, 16),
27545 => conv_std_logic_vector(16371, 16),
27546 => conv_std_logic_vector(16478, 16),
27547 => conv_std_logic_vector(16585, 16),
27548 => conv_std_logic_vector(16692, 16),
27549 => conv_std_logic_vector(16799, 16),
27550 => conv_std_logic_vector(16906, 16),
27551 => conv_std_logic_vector(17013, 16),
27552 => conv_std_logic_vector(17120, 16),
27553 => conv_std_logic_vector(17227, 16),
27554 => conv_std_logic_vector(17334, 16),
27555 => conv_std_logic_vector(17441, 16),
27556 => conv_std_logic_vector(17548, 16),
27557 => conv_std_logic_vector(17655, 16),
27558 => conv_std_logic_vector(17762, 16),
27559 => conv_std_logic_vector(17869, 16),
27560 => conv_std_logic_vector(17976, 16),
27561 => conv_std_logic_vector(18083, 16),
27562 => conv_std_logic_vector(18190, 16),
27563 => conv_std_logic_vector(18297, 16),
27564 => conv_std_logic_vector(18404, 16),
27565 => conv_std_logic_vector(18511, 16),
27566 => conv_std_logic_vector(18618, 16),
27567 => conv_std_logic_vector(18725, 16),
27568 => conv_std_logic_vector(18832, 16),
27569 => conv_std_logic_vector(18939, 16),
27570 => conv_std_logic_vector(19046, 16),
27571 => conv_std_logic_vector(19153, 16),
27572 => conv_std_logic_vector(19260, 16),
27573 => conv_std_logic_vector(19367, 16),
27574 => conv_std_logic_vector(19474, 16),
27575 => conv_std_logic_vector(19581, 16),
27576 => conv_std_logic_vector(19688, 16),
27577 => conv_std_logic_vector(19795, 16),
27578 => conv_std_logic_vector(19902, 16),
27579 => conv_std_logic_vector(20009, 16),
27580 => conv_std_logic_vector(20116, 16),
27581 => conv_std_logic_vector(20223, 16),
27582 => conv_std_logic_vector(20330, 16),
27583 => conv_std_logic_vector(20437, 16),
27584 => conv_std_logic_vector(20544, 16),
27585 => conv_std_logic_vector(20651, 16),
27586 => conv_std_logic_vector(20758, 16),
27587 => conv_std_logic_vector(20865, 16),
27588 => conv_std_logic_vector(20972, 16),
27589 => conv_std_logic_vector(21079, 16),
27590 => conv_std_logic_vector(21186, 16),
27591 => conv_std_logic_vector(21293, 16),
27592 => conv_std_logic_vector(21400, 16),
27593 => conv_std_logic_vector(21507, 16),
27594 => conv_std_logic_vector(21614, 16),
27595 => conv_std_logic_vector(21721, 16),
27596 => conv_std_logic_vector(21828, 16),
27597 => conv_std_logic_vector(21935, 16),
27598 => conv_std_logic_vector(22042, 16),
27599 => conv_std_logic_vector(22149, 16),
27600 => conv_std_logic_vector(22256, 16),
27601 => conv_std_logic_vector(22363, 16),
27602 => conv_std_logic_vector(22470, 16),
27603 => conv_std_logic_vector(22577, 16),
27604 => conv_std_logic_vector(22684, 16),
27605 => conv_std_logic_vector(22791, 16),
27606 => conv_std_logic_vector(22898, 16),
27607 => conv_std_logic_vector(23005, 16),
27608 => conv_std_logic_vector(23112, 16),
27609 => conv_std_logic_vector(23219, 16),
27610 => conv_std_logic_vector(23326, 16),
27611 => conv_std_logic_vector(23433, 16),
27612 => conv_std_logic_vector(23540, 16),
27613 => conv_std_logic_vector(23647, 16),
27614 => conv_std_logic_vector(23754, 16),
27615 => conv_std_logic_vector(23861, 16),
27616 => conv_std_logic_vector(23968, 16),
27617 => conv_std_logic_vector(24075, 16),
27618 => conv_std_logic_vector(24182, 16),
27619 => conv_std_logic_vector(24289, 16),
27620 => conv_std_logic_vector(24396, 16),
27621 => conv_std_logic_vector(24503, 16),
27622 => conv_std_logic_vector(24610, 16),
27623 => conv_std_logic_vector(24717, 16),
27624 => conv_std_logic_vector(24824, 16),
27625 => conv_std_logic_vector(24931, 16),
27626 => conv_std_logic_vector(25038, 16),
27627 => conv_std_logic_vector(25145, 16),
27628 => conv_std_logic_vector(25252, 16),
27629 => conv_std_logic_vector(25359, 16),
27630 => conv_std_logic_vector(25466, 16),
27631 => conv_std_logic_vector(25573, 16),
27632 => conv_std_logic_vector(25680, 16),
27633 => conv_std_logic_vector(25787, 16),
27634 => conv_std_logic_vector(25894, 16),
27635 => conv_std_logic_vector(26001, 16),
27636 => conv_std_logic_vector(26108, 16),
27637 => conv_std_logic_vector(26215, 16),
27638 => conv_std_logic_vector(26322, 16),
27639 => conv_std_logic_vector(26429, 16),
27640 => conv_std_logic_vector(26536, 16),
27641 => conv_std_logic_vector(26643, 16),
27642 => conv_std_logic_vector(26750, 16),
27643 => conv_std_logic_vector(26857, 16),
27644 => conv_std_logic_vector(26964, 16),
27645 => conv_std_logic_vector(27071, 16),
27646 => conv_std_logic_vector(27178, 16),
27647 => conv_std_logic_vector(27285, 16),
27648 => conv_std_logic_vector(0, 16),
27649 => conv_std_logic_vector(108, 16),
27650 => conv_std_logic_vector(216, 16),
27651 => conv_std_logic_vector(324, 16),
27652 => conv_std_logic_vector(432, 16),
27653 => conv_std_logic_vector(540, 16),
27654 => conv_std_logic_vector(648, 16),
27655 => conv_std_logic_vector(756, 16),
27656 => conv_std_logic_vector(864, 16),
27657 => conv_std_logic_vector(972, 16),
27658 => conv_std_logic_vector(1080, 16),
27659 => conv_std_logic_vector(1188, 16),
27660 => conv_std_logic_vector(1296, 16),
27661 => conv_std_logic_vector(1404, 16),
27662 => conv_std_logic_vector(1512, 16),
27663 => conv_std_logic_vector(1620, 16),
27664 => conv_std_logic_vector(1728, 16),
27665 => conv_std_logic_vector(1836, 16),
27666 => conv_std_logic_vector(1944, 16),
27667 => conv_std_logic_vector(2052, 16),
27668 => conv_std_logic_vector(2160, 16),
27669 => conv_std_logic_vector(2268, 16),
27670 => conv_std_logic_vector(2376, 16),
27671 => conv_std_logic_vector(2484, 16),
27672 => conv_std_logic_vector(2592, 16),
27673 => conv_std_logic_vector(2700, 16),
27674 => conv_std_logic_vector(2808, 16),
27675 => conv_std_logic_vector(2916, 16),
27676 => conv_std_logic_vector(3024, 16),
27677 => conv_std_logic_vector(3132, 16),
27678 => conv_std_logic_vector(3240, 16),
27679 => conv_std_logic_vector(3348, 16),
27680 => conv_std_logic_vector(3456, 16),
27681 => conv_std_logic_vector(3564, 16),
27682 => conv_std_logic_vector(3672, 16),
27683 => conv_std_logic_vector(3780, 16),
27684 => conv_std_logic_vector(3888, 16),
27685 => conv_std_logic_vector(3996, 16),
27686 => conv_std_logic_vector(4104, 16),
27687 => conv_std_logic_vector(4212, 16),
27688 => conv_std_logic_vector(4320, 16),
27689 => conv_std_logic_vector(4428, 16),
27690 => conv_std_logic_vector(4536, 16),
27691 => conv_std_logic_vector(4644, 16),
27692 => conv_std_logic_vector(4752, 16),
27693 => conv_std_logic_vector(4860, 16),
27694 => conv_std_logic_vector(4968, 16),
27695 => conv_std_logic_vector(5076, 16),
27696 => conv_std_logic_vector(5184, 16),
27697 => conv_std_logic_vector(5292, 16),
27698 => conv_std_logic_vector(5400, 16),
27699 => conv_std_logic_vector(5508, 16),
27700 => conv_std_logic_vector(5616, 16),
27701 => conv_std_logic_vector(5724, 16),
27702 => conv_std_logic_vector(5832, 16),
27703 => conv_std_logic_vector(5940, 16),
27704 => conv_std_logic_vector(6048, 16),
27705 => conv_std_logic_vector(6156, 16),
27706 => conv_std_logic_vector(6264, 16),
27707 => conv_std_logic_vector(6372, 16),
27708 => conv_std_logic_vector(6480, 16),
27709 => conv_std_logic_vector(6588, 16),
27710 => conv_std_logic_vector(6696, 16),
27711 => conv_std_logic_vector(6804, 16),
27712 => conv_std_logic_vector(6912, 16),
27713 => conv_std_logic_vector(7020, 16),
27714 => conv_std_logic_vector(7128, 16),
27715 => conv_std_logic_vector(7236, 16),
27716 => conv_std_logic_vector(7344, 16),
27717 => conv_std_logic_vector(7452, 16),
27718 => conv_std_logic_vector(7560, 16),
27719 => conv_std_logic_vector(7668, 16),
27720 => conv_std_logic_vector(7776, 16),
27721 => conv_std_logic_vector(7884, 16),
27722 => conv_std_logic_vector(7992, 16),
27723 => conv_std_logic_vector(8100, 16),
27724 => conv_std_logic_vector(8208, 16),
27725 => conv_std_logic_vector(8316, 16),
27726 => conv_std_logic_vector(8424, 16),
27727 => conv_std_logic_vector(8532, 16),
27728 => conv_std_logic_vector(8640, 16),
27729 => conv_std_logic_vector(8748, 16),
27730 => conv_std_logic_vector(8856, 16),
27731 => conv_std_logic_vector(8964, 16),
27732 => conv_std_logic_vector(9072, 16),
27733 => conv_std_logic_vector(9180, 16),
27734 => conv_std_logic_vector(9288, 16),
27735 => conv_std_logic_vector(9396, 16),
27736 => conv_std_logic_vector(9504, 16),
27737 => conv_std_logic_vector(9612, 16),
27738 => conv_std_logic_vector(9720, 16),
27739 => conv_std_logic_vector(9828, 16),
27740 => conv_std_logic_vector(9936, 16),
27741 => conv_std_logic_vector(10044, 16),
27742 => conv_std_logic_vector(10152, 16),
27743 => conv_std_logic_vector(10260, 16),
27744 => conv_std_logic_vector(10368, 16),
27745 => conv_std_logic_vector(10476, 16),
27746 => conv_std_logic_vector(10584, 16),
27747 => conv_std_logic_vector(10692, 16),
27748 => conv_std_logic_vector(10800, 16),
27749 => conv_std_logic_vector(10908, 16),
27750 => conv_std_logic_vector(11016, 16),
27751 => conv_std_logic_vector(11124, 16),
27752 => conv_std_logic_vector(11232, 16),
27753 => conv_std_logic_vector(11340, 16),
27754 => conv_std_logic_vector(11448, 16),
27755 => conv_std_logic_vector(11556, 16),
27756 => conv_std_logic_vector(11664, 16),
27757 => conv_std_logic_vector(11772, 16),
27758 => conv_std_logic_vector(11880, 16),
27759 => conv_std_logic_vector(11988, 16),
27760 => conv_std_logic_vector(12096, 16),
27761 => conv_std_logic_vector(12204, 16),
27762 => conv_std_logic_vector(12312, 16),
27763 => conv_std_logic_vector(12420, 16),
27764 => conv_std_logic_vector(12528, 16),
27765 => conv_std_logic_vector(12636, 16),
27766 => conv_std_logic_vector(12744, 16),
27767 => conv_std_logic_vector(12852, 16),
27768 => conv_std_logic_vector(12960, 16),
27769 => conv_std_logic_vector(13068, 16),
27770 => conv_std_logic_vector(13176, 16),
27771 => conv_std_logic_vector(13284, 16),
27772 => conv_std_logic_vector(13392, 16),
27773 => conv_std_logic_vector(13500, 16),
27774 => conv_std_logic_vector(13608, 16),
27775 => conv_std_logic_vector(13716, 16),
27776 => conv_std_logic_vector(13824, 16),
27777 => conv_std_logic_vector(13932, 16),
27778 => conv_std_logic_vector(14040, 16),
27779 => conv_std_logic_vector(14148, 16),
27780 => conv_std_logic_vector(14256, 16),
27781 => conv_std_logic_vector(14364, 16),
27782 => conv_std_logic_vector(14472, 16),
27783 => conv_std_logic_vector(14580, 16),
27784 => conv_std_logic_vector(14688, 16),
27785 => conv_std_logic_vector(14796, 16),
27786 => conv_std_logic_vector(14904, 16),
27787 => conv_std_logic_vector(15012, 16),
27788 => conv_std_logic_vector(15120, 16),
27789 => conv_std_logic_vector(15228, 16),
27790 => conv_std_logic_vector(15336, 16),
27791 => conv_std_logic_vector(15444, 16),
27792 => conv_std_logic_vector(15552, 16),
27793 => conv_std_logic_vector(15660, 16),
27794 => conv_std_logic_vector(15768, 16),
27795 => conv_std_logic_vector(15876, 16),
27796 => conv_std_logic_vector(15984, 16),
27797 => conv_std_logic_vector(16092, 16),
27798 => conv_std_logic_vector(16200, 16),
27799 => conv_std_logic_vector(16308, 16),
27800 => conv_std_logic_vector(16416, 16),
27801 => conv_std_logic_vector(16524, 16),
27802 => conv_std_logic_vector(16632, 16),
27803 => conv_std_logic_vector(16740, 16),
27804 => conv_std_logic_vector(16848, 16),
27805 => conv_std_logic_vector(16956, 16),
27806 => conv_std_logic_vector(17064, 16),
27807 => conv_std_logic_vector(17172, 16),
27808 => conv_std_logic_vector(17280, 16),
27809 => conv_std_logic_vector(17388, 16),
27810 => conv_std_logic_vector(17496, 16),
27811 => conv_std_logic_vector(17604, 16),
27812 => conv_std_logic_vector(17712, 16),
27813 => conv_std_logic_vector(17820, 16),
27814 => conv_std_logic_vector(17928, 16),
27815 => conv_std_logic_vector(18036, 16),
27816 => conv_std_logic_vector(18144, 16),
27817 => conv_std_logic_vector(18252, 16),
27818 => conv_std_logic_vector(18360, 16),
27819 => conv_std_logic_vector(18468, 16),
27820 => conv_std_logic_vector(18576, 16),
27821 => conv_std_logic_vector(18684, 16),
27822 => conv_std_logic_vector(18792, 16),
27823 => conv_std_logic_vector(18900, 16),
27824 => conv_std_logic_vector(19008, 16),
27825 => conv_std_logic_vector(19116, 16),
27826 => conv_std_logic_vector(19224, 16),
27827 => conv_std_logic_vector(19332, 16),
27828 => conv_std_logic_vector(19440, 16),
27829 => conv_std_logic_vector(19548, 16),
27830 => conv_std_logic_vector(19656, 16),
27831 => conv_std_logic_vector(19764, 16),
27832 => conv_std_logic_vector(19872, 16),
27833 => conv_std_logic_vector(19980, 16),
27834 => conv_std_logic_vector(20088, 16),
27835 => conv_std_logic_vector(20196, 16),
27836 => conv_std_logic_vector(20304, 16),
27837 => conv_std_logic_vector(20412, 16),
27838 => conv_std_logic_vector(20520, 16),
27839 => conv_std_logic_vector(20628, 16),
27840 => conv_std_logic_vector(20736, 16),
27841 => conv_std_logic_vector(20844, 16),
27842 => conv_std_logic_vector(20952, 16),
27843 => conv_std_logic_vector(21060, 16),
27844 => conv_std_logic_vector(21168, 16),
27845 => conv_std_logic_vector(21276, 16),
27846 => conv_std_logic_vector(21384, 16),
27847 => conv_std_logic_vector(21492, 16),
27848 => conv_std_logic_vector(21600, 16),
27849 => conv_std_logic_vector(21708, 16),
27850 => conv_std_logic_vector(21816, 16),
27851 => conv_std_logic_vector(21924, 16),
27852 => conv_std_logic_vector(22032, 16),
27853 => conv_std_logic_vector(22140, 16),
27854 => conv_std_logic_vector(22248, 16),
27855 => conv_std_logic_vector(22356, 16),
27856 => conv_std_logic_vector(22464, 16),
27857 => conv_std_logic_vector(22572, 16),
27858 => conv_std_logic_vector(22680, 16),
27859 => conv_std_logic_vector(22788, 16),
27860 => conv_std_logic_vector(22896, 16),
27861 => conv_std_logic_vector(23004, 16),
27862 => conv_std_logic_vector(23112, 16),
27863 => conv_std_logic_vector(23220, 16),
27864 => conv_std_logic_vector(23328, 16),
27865 => conv_std_logic_vector(23436, 16),
27866 => conv_std_logic_vector(23544, 16),
27867 => conv_std_logic_vector(23652, 16),
27868 => conv_std_logic_vector(23760, 16),
27869 => conv_std_logic_vector(23868, 16),
27870 => conv_std_logic_vector(23976, 16),
27871 => conv_std_logic_vector(24084, 16),
27872 => conv_std_logic_vector(24192, 16),
27873 => conv_std_logic_vector(24300, 16),
27874 => conv_std_logic_vector(24408, 16),
27875 => conv_std_logic_vector(24516, 16),
27876 => conv_std_logic_vector(24624, 16),
27877 => conv_std_logic_vector(24732, 16),
27878 => conv_std_logic_vector(24840, 16),
27879 => conv_std_logic_vector(24948, 16),
27880 => conv_std_logic_vector(25056, 16),
27881 => conv_std_logic_vector(25164, 16),
27882 => conv_std_logic_vector(25272, 16),
27883 => conv_std_logic_vector(25380, 16),
27884 => conv_std_logic_vector(25488, 16),
27885 => conv_std_logic_vector(25596, 16),
27886 => conv_std_logic_vector(25704, 16),
27887 => conv_std_logic_vector(25812, 16),
27888 => conv_std_logic_vector(25920, 16),
27889 => conv_std_logic_vector(26028, 16),
27890 => conv_std_logic_vector(26136, 16),
27891 => conv_std_logic_vector(26244, 16),
27892 => conv_std_logic_vector(26352, 16),
27893 => conv_std_logic_vector(26460, 16),
27894 => conv_std_logic_vector(26568, 16),
27895 => conv_std_logic_vector(26676, 16),
27896 => conv_std_logic_vector(26784, 16),
27897 => conv_std_logic_vector(26892, 16),
27898 => conv_std_logic_vector(27000, 16),
27899 => conv_std_logic_vector(27108, 16),
27900 => conv_std_logic_vector(27216, 16),
27901 => conv_std_logic_vector(27324, 16),
27902 => conv_std_logic_vector(27432, 16),
27903 => conv_std_logic_vector(27540, 16),
27904 => conv_std_logic_vector(0, 16),
27905 => conv_std_logic_vector(109, 16),
27906 => conv_std_logic_vector(218, 16),
27907 => conv_std_logic_vector(327, 16),
27908 => conv_std_logic_vector(436, 16),
27909 => conv_std_logic_vector(545, 16),
27910 => conv_std_logic_vector(654, 16),
27911 => conv_std_logic_vector(763, 16),
27912 => conv_std_logic_vector(872, 16),
27913 => conv_std_logic_vector(981, 16),
27914 => conv_std_logic_vector(1090, 16),
27915 => conv_std_logic_vector(1199, 16),
27916 => conv_std_logic_vector(1308, 16),
27917 => conv_std_logic_vector(1417, 16),
27918 => conv_std_logic_vector(1526, 16),
27919 => conv_std_logic_vector(1635, 16),
27920 => conv_std_logic_vector(1744, 16),
27921 => conv_std_logic_vector(1853, 16),
27922 => conv_std_logic_vector(1962, 16),
27923 => conv_std_logic_vector(2071, 16),
27924 => conv_std_logic_vector(2180, 16),
27925 => conv_std_logic_vector(2289, 16),
27926 => conv_std_logic_vector(2398, 16),
27927 => conv_std_logic_vector(2507, 16),
27928 => conv_std_logic_vector(2616, 16),
27929 => conv_std_logic_vector(2725, 16),
27930 => conv_std_logic_vector(2834, 16),
27931 => conv_std_logic_vector(2943, 16),
27932 => conv_std_logic_vector(3052, 16),
27933 => conv_std_logic_vector(3161, 16),
27934 => conv_std_logic_vector(3270, 16),
27935 => conv_std_logic_vector(3379, 16),
27936 => conv_std_logic_vector(3488, 16),
27937 => conv_std_logic_vector(3597, 16),
27938 => conv_std_logic_vector(3706, 16),
27939 => conv_std_logic_vector(3815, 16),
27940 => conv_std_logic_vector(3924, 16),
27941 => conv_std_logic_vector(4033, 16),
27942 => conv_std_logic_vector(4142, 16),
27943 => conv_std_logic_vector(4251, 16),
27944 => conv_std_logic_vector(4360, 16),
27945 => conv_std_logic_vector(4469, 16),
27946 => conv_std_logic_vector(4578, 16),
27947 => conv_std_logic_vector(4687, 16),
27948 => conv_std_logic_vector(4796, 16),
27949 => conv_std_logic_vector(4905, 16),
27950 => conv_std_logic_vector(5014, 16),
27951 => conv_std_logic_vector(5123, 16),
27952 => conv_std_logic_vector(5232, 16),
27953 => conv_std_logic_vector(5341, 16),
27954 => conv_std_logic_vector(5450, 16),
27955 => conv_std_logic_vector(5559, 16),
27956 => conv_std_logic_vector(5668, 16),
27957 => conv_std_logic_vector(5777, 16),
27958 => conv_std_logic_vector(5886, 16),
27959 => conv_std_logic_vector(5995, 16),
27960 => conv_std_logic_vector(6104, 16),
27961 => conv_std_logic_vector(6213, 16),
27962 => conv_std_logic_vector(6322, 16),
27963 => conv_std_logic_vector(6431, 16),
27964 => conv_std_logic_vector(6540, 16),
27965 => conv_std_logic_vector(6649, 16),
27966 => conv_std_logic_vector(6758, 16),
27967 => conv_std_logic_vector(6867, 16),
27968 => conv_std_logic_vector(6976, 16),
27969 => conv_std_logic_vector(7085, 16),
27970 => conv_std_logic_vector(7194, 16),
27971 => conv_std_logic_vector(7303, 16),
27972 => conv_std_logic_vector(7412, 16),
27973 => conv_std_logic_vector(7521, 16),
27974 => conv_std_logic_vector(7630, 16),
27975 => conv_std_logic_vector(7739, 16),
27976 => conv_std_logic_vector(7848, 16),
27977 => conv_std_logic_vector(7957, 16),
27978 => conv_std_logic_vector(8066, 16),
27979 => conv_std_logic_vector(8175, 16),
27980 => conv_std_logic_vector(8284, 16),
27981 => conv_std_logic_vector(8393, 16),
27982 => conv_std_logic_vector(8502, 16),
27983 => conv_std_logic_vector(8611, 16),
27984 => conv_std_logic_vector(8720, 16),
27985 => conv_std_logic_vector(8829, 16),
27986 => conv_std_logic_vector(8938, 16),
27987 => conv_std_logic_vector(9047, 16),
27988 => conv_std_logic_vector(9156, 16),
27989 => conv_std_logic_vector(9265, 16),
27990 => conv_std_logic_vector(9374, 16),
27991 => conv_std_logic_vector(9483, 16),
27992 => conv_std_logic_vector(9592, 16),
27993 => conv_std_logic_vector(9701, 16),
27994 => conv_std_logic_vector(9810, 16),
27995 => conv_std_logic_vector(9919, 16),
27996 => conv_std_logic_vector(10028, 16),
27997 => conv_std_logic_vector(10137, 16),
27998 => conv_std_logic_vector(10246, 16),
27999 => conv_std_logic_vector(10355, 16),
28000 => conv_std_logic_vector(10464, 16),
28001 => conv_std_logic_vector(10573, 16),
28002 => conv_std_logic_vector(10682, 16),
28003 => conv_std_logic_vector(10791, 16),
28004 => conv_std_logic_vector(10900, 16),
28005 => conv_std_logic_vector(11009, 16),
28006 => conv_std_logic_vector(11118, 16),
28007 => conv_std_logic_vector(11227, 16),
28008 => conv_std_logic_vector(11336, 16),
28009 => conv_std_logic_vector(11445, 16),
28010 => conv_std_logic_vector(11554, 16),
28011 => conv_std_logic_vector(11663, 16),
28012 => conv_std_logic_vector(11772, 16),
28013 => conv_std_logic_vector(11881, 16),
28014 => conv_std_logic_vector(11990, 16),
28015 => conv_std_logic_vector(12099, 16),
28016 => conv_std_logic_vector(12208, 16),
28017 => conv_std_logic_vector(12317, 16),
28018 => conv_std_logic_vector(12426, 16),
28019 => conv_std_logic_vector(12535, 16),
28020 => conv_std_logic_vector(12644, 16),
28021 => conv_std_logic_vector(12753, 16),
28022 => conv_std_logic_vector(12862, 16),
28023 => conv_std_logic_vector(12971, 16),
28024 => conv_std_logic_vector(13080, 16),
28025 => conv_std_logic_vector(13189, 16),
28026 => conv_std_logic_vector(13298, 16),
28027 => conv_std_logic_vector(13407, 16),
28028 => conv_std_logic_vector(13516, 16),
28029 => conv_std_logic_vector(13625, 16),
28030 => conv_std_logic_vector(13734, 16),
28031 => conv_std_logic_vector(13843, 16),
28032 => conv_std_logic_vector(13952, 16),
28033 => conv_std_logic_vector(14061, 16),
28034 => conv_std_logic_vector(14170, 16),
28035 => conv_std_logic_vector(14279, 16),
28036 => conv_std_logic_vector(14388, 16),
28037 => conv_std_logic_vector(14497, 16),
28038 => conv_std_logic_vector(14606, 16),
28039 => conv_std_logic_vector(14715, 16),
28040 => conv_std_logic_vector(14824, 16),
28041 => conv_std_logic_vector(14933, 16),
28042 => conv_std_logic_vector(15042, 16),
28043 => conv_std_logic_vector(15151, 16),
28044 => conv_std_logic_vector(15260, 16),
28045 => conv_std_logic_vector(15369, 16),
28046 => conv_std_logic_vector(15478, 16),
28047 => conv_std_logic_vector(15587, 16),
28048 => conv_std_logic_vector(15696, 16),
28049 => conv_std_logic_vector(15805, 16),
28050 => conv_std_logic_vector(15914, 16),
28051 => conv_std_logic_vector(16023, 16),
28052 => conv_std_logic_vector(16132, 16),
28053 => conv_std_logic_vector(16241, 16),
28054 => conv_std_logic_vector(16350, 16),
28055 => conv_std_logic_vector(16459, 16),
28056 => conv_std_logic_vector(16568, 16),
28057 => conv_std_logic_vector(16677, 16),
28058 => conv_std_logic_vector(16786, 16),
28059 => conv_std_logic_vector(16895, 16),
28060 => conv_std_logic_vector(17004, 16),
28061 => conv_std_logic_vector(17113, 16),
28062 => conv_std_logic_vector(17222, 16),
28063 => conv_std_logic_vector(17331, 16),
28064 => conv_std_logic_vector(17440, 16),
28065 => conv_std_logic_vector(17549, 16),
28066 => conv_std_logic_vector(17658, 16),
28067 => conv_std_logic_vector(17767, 16),
28068 => conv_std_logic_vector(17876, 16),
28069 => conv_std_logic_vector(17985, 16),
28070 => conv_std_logic_vector(18094, 16),
28071 => conv_std_logic_vector(18203, 16),
28072 => conv_std_logic_vector(18312, 16),
28073 => conv_std_logic_vector(18421, 16),
28074 => conv_std_logic_vector(18530, 16),
28075 => conv_std_logic_vector(18639, 16),
28076 => conv_std_logic_vector(18748, 16),
28077 => conv_std_logic_vector(18857, 16),
28078 => conv_std_logic_vector(18966, 16),
28079 => conv_std_logic_vector(19075, 16),
28080 => conv_std_logic_vector(19184, 16),
28081 => conv_std_logic_vector(19293, 16),
28082 => conv_std_logic_vector(19402, 16),
28083 => conv_std_logic_vector(19511, 16),
28084 => conv_std_logic_vector(19620, 16),
28085 => conv_std_logic_vector(19729, 16),
28086 => conv_std_logic_vector(19838, 16),
28087 => conv_std_logic_vector(19947, 16),
28088 => conv_std_logic_vector(20056, 16),
28089 => conv_std_logic_vector(20165, 16),
28090 => conv_std_logic_vector(20274, 16),
28091 => conv_std_logic_vector(20383, 16),
28092 => conv_std_logic_vector(20492, 16),
28093 => conv_std_logic_vector(20601, 16),
28094 => conv_std_logic_vector(20710, 16),
28095 => conv_std_logic_vector(20819, 16),
28096 => conv_std_logic_vector(20928, 16),
28097 => conv_std_logic_vector(21037, 16),
28098 => conv_std_logic_vector(21146, 16),
28099 => conv_std_logic_vector(21255, 16),
28100 => conv_std_logic_vector(21364, 16),
28101 => conv_std_logic_vector(21473, 16),
28102 => conv_std_logic_vector(21582, 16),
28103 => conv_std_logic_vector(21691, 16),
28104 => conv_std_logic_vector(21800, 16),
28105 => conv_std_logic_vector(21909, 16),
28106 => conv_std_logic_vector(22018, 16),
28107 => conv_std_logic_vector(22127, 16),
28108 => conv_std_logic_vector(22236, 16),
28109 => conv_std_logic_vector(22345, 16),
28110 => conv_std_logic_vector(22454, 16),
28111 => conv_std_logic_vector(22563, 16),
28112 => conv_std_logic_vector(22672, 16),
28113 => conv_std_logic_vector(22781, 16),
28114 => conv_std_logic_vector(22890, 16),
28115 => conv_std_logic_vector(22999, 16),
28116 => conv_std_logic_vector(23108, 16),
28117 => conv_std_logic_vector(23217, 16),
28118 => conv_std_logic_vector(23326, 16),
28119 => conv_std_logic_vector(23435, 16),
28120 => conv_std_logic_vector(23544, 16),
28121 => conv_std_logic_vector(23653, 16),
28122 => conv_std_logic_vector(23762, 16),
28123 => conv_std_logic_vector(23871, 16),
28124 => conv_std_logic_vector(23980, 16),
28125 => conv_std_logic_vector(24089, 16),
28126 => conv_std_logic_vector(24198, 16),
28127 => conv_std_logic_vector(24307, 16),
28128 => conv_std_logic_vector(24416, 16),
28129 => conv_std_logic_vector(24525, 16),
28130 => conv_std_logic_vector(24634, 16),
28131 => conv_std_logic_vector(24743, 16),
28132 => conv_std_logic_vector(24852, 16),
28133 => conv_std_logic_vector(24961, 16),
28134 => conv_std_logic_vector(25070, 16),
28135 => conv_std_logic_vector(25179, 16),
28136 => conv_std_logic_vector(25288, 16),
28137 => conv_std_logic_vector(25397, 16),
28138 => conv_std_logic_vector(25506, 16),
28139 => conv_std_logic_vector(25615, 16),
28140 => conv_std_logic_vector(25724, 16),
28141 => conv_std_logic_vector(25833, 16),
28142 => conv_std_logic_vector(25942, 16),
28143 => conv_std_logic_vector(26051, 16),
28144 => conv_std_logic_vector(26160, 16),
28145 => conv_std_logic_vector(26269, 16),
28146 => conv_std_logic_vector(26378, 16),
28147 => conv_std_logic_vector(26487, 16),
28148 => conv_std_logic_vector(26596, 16),
28149 => conv_std_logic_vector(26705, 16),
28150 => conv_std_logic_vector(26814, 16),
28151 => conv_std_logic_vector(26923, 16),
28152 => conv_std_logic_vector(27032, 16),
28153 => conv_std_logic_vector(27141, 16),
28154 => conv_std_logic_vector(27250, 16),
28155 => conv_std_logic_vector(27359, 16),
28156 => conv_std_logic_vector(27468, 16),
28157 => conv_std_logic_vector(27577, 16),
28158 => conv_std_logic_vector(27686, 16),
28159 => conv_std_logic_vector(27795, 16),
28160 => conv_std_logic_vector(0, 16),
28161 => conv_std_logic_vector(110, 16),
28162 => conv_std_logic_vector(220, 16),
28163 => conv_std_logic_vector(330, 16),
28164 => conv_std_logic_vector(440, 16),
28165 => conv_std_logic_vector(550, 16),
28166 => conv_std_logic_vector(660, 16),
28167 => conv_std_logic_vector(770, 16),
28168 => conv_std_logic_vector(880, 16),
28169 => conv_std_logic_vector(990, 16),
28170 => conv_std_logic_vector(1100, 16),
28171 => conv_std_logic_vector(1210, 16),
28172 => conv_std_logic_vector(1320, 16),
28173 => conv_std_logic_vector(1430, 16),
28174 => conv_std_logic_vector(1540, 16),
28175 => conv_std_logic_vector(1650, 16),
28176 => conv_std_logic_vector(1760, 16),
28177 => conv_std_logic_vector(1870, 16),
28178 => conv_std_logic_vector(1980, 16),
28179 => conv_std_logic_vector(2090, 16),
28180 => conv_std_logic_vector(2200, 16),
28181 => conv_std_logic_vector(2310, 16),
28182 => conv_std_logic_vector(2420, 16),
28183 => conv_std_logic_vector(2530, 16),
28184 => conv_std_logic_vector(2640, 16),
28185 => conv_std_logic_vector(2750, 16),
28186 => conv_std_logic_vector(2860, 16),
28187 => conv_std_logic_vector(2970, 16),
28188 => conv_std_logic_vector(3080, 16),
28189 => conv_std_logic_vector(3190, 16),
28190 => conv_std_logic_vector(3300, 16),
28191 => conv_std_logic_vector(3410, 16),
28192 => conv_std_logic_vector(3520, 16),
28193 => conv_std_logic_vector(3630, 16),
28194 => conv_std_logic_vector(3740, 16),
28195 => conv_std_logic_vector(3850, 16),
28196 => conv_std_logic_vector(3960, 16),
28197 => conv_std_logic_vector(4070, 16),
28198 => conv_std_logic_vector(4180, 16),
28199 => conv_std_logic_vector(4290, 16),
28200 => conv_std_logic_vector(4400, 16),
28201 => conv_std_logic_vector(4510, 16),
28202 => conv_std_logic_vector(4620, 16),
28203 => conv_std_logic_vector(4730, 16),
28204 => conv_std_logic_vector(4840, 16),
28205 => conv_std_logic_vector(4950, 16),
28206 => conv_std_logic_vector(5060, 16),
28207 => conv_std_logic_vector(5170, 16),
28208 => conv_std_logic_vector(5280, 16),
28209 => conv_std_logic_vector(5390, 16),
28210 => conv_std_logic_vector(5500, 16),
28211 => conv_std_logic_vector(5610, 16),
28212 => conv_std_logic_vector(5720, 16),
28213 => conv_std_logic_vector(5830, 16),
28214 => conv_std_logic_vector(5940, 16),
28215 => conv_std_logic_vector(6050, 16),
28216 => conv_std_logic_vector(6160, 16),
28217 => conv_std_logic_vector(6270, 16),
28218 => conv_std_logic_vector(6380, 16),
28219 => conv_std_logic_vector(6490, 16),
28220 => conv_std_logic_vector(6600, 16),
28221 => conv_std_logic_vector(6710, 16),
28222 => conv_std_logic_vector(6820, 16),
28223 => conv_std_logic_vector(6930, 16),
28224 => conv_std_logic_vector(7040, 16),
28225 => conv_std_logic_vector(7150, 16),
28226 => conv_std_logic_vector(7260, 16),
28227 => conv_std_logic_vector(7370, 16),
28228 => conv_std_logic_vector(7480, 16),
28229 => conv_std_logic_vector(7590, 16),
28230 => conv_std_logic_vector(7700, 16),
28231 => conv_std_logic_vector(7810, 16),
28232 => conv_std_logic_vector(7920, 16),
28233 => conv_std_logic_vector(8030, 16),
28234 => conv_std_logic_vector(8140, 16),
28235 => conv_std_logic_vector(8250, 16),
28236 => conv_std_logic_vector(8360, 16),
28237 => conv_std_logic_vector(8470, 16),
28238 => conv_std_logic_vector(8580, 16),
28239 => conv_std_logic_vector(8690, 16),
28240 => conv_std_logic_vector(8800, 16),
28241 => conv_std_logic_vector(8910, 16),
28242 => conv_std_logic_vector(9020, 16),
28243 => conv_std_logic_vector(9130, 16),
28244 => conv_std_logic_vector(9240, 16),
28245 => conv_std_logic_vector(9350, 16),
28246 => conv_std_logic_vector(9460, 16),
28247 => conv_std_logic_vector(9570, 16),
28248 => conv_std_logic_vector(9680, 16),
28249 => conv_std_logic_vector(9790, 16),
28250 => conv_std_logic_vector(9900, 16),
28251 => conv_std_logic_vector(10010, 16),
28252 => conv_std_logic_vector(10120, 16),
28253 => conv_std_logic_vector(10230, 16),
28254 => conv_std_logic_vector(10340, 16),
28255 => conv_std_logic_vector(10450, 16),
28256 => conv_std_logic_vector(10560, 16),
28257 => conv_std_logic_vector(10670, 16),
28258 => conv_std_logic_vector(10780, 16),
28259 => conv_std_logic_vector(10890, 16),
28260 => conv_std_logic_vector(11000, 16),
28261 => conv_std_logic_vector(11110, 16),
28262 => conv_std_logic_vector(11220, 16),
28263 => conv_std_logic_vector(11330, 16),
28264 => conv_std_logic_vector(11440, 16),
28265 => conv_std_logic_vector(11550, 16),
28266 => conv_std_logic_vector(11660, 16),
28267 => conv_std_logic_vector(11770, 16),
28268 => conv_std_logic_vector(11880, 16),
28269 => conv_std_logic_vector(11990, 16),
28270 => conv_std_logic_vector(12100, 16),
28271 => conv_std_logic_vector(12210, 16),
28272 => conv_std_logic_vector(12320, 16),
28273 => conv_std_logic_vector(12430, 16),
28274 => conv_std_logic_vector(12540, 16),
28275 => conv_std_logic_vector(12650, 16),
28276 => conv_std_logic_vector(12760, 16),
28277 => conv_std_logic_vector(12870, 16),
28278 => conv_std_logic_vector(12980, 16),
28279 => conv_std_logic_vector(13090, 16),
28280 => conv_std_logic_vector(13200, 16),
28281 => conv_std_logic_vector(13310, 16),
28282 => conv_std_logic_vector(13420, 16),
28283 => conv_std_logic_vector(13530, 16),
28284 => conv_std_logic_vector(13640, 16),
28285 => conv_std_logic_vector(13750, 16),
28286 => conv_std_logic_vector(13860, 16),
28287 => conv_std_logic_vector(13970, 16),
28288 => conv_std_logic_vector(14080, 16),
28289 => conv_std_logic_vector(14190, 16),
28290 => conv_std_logic_vector(14300, 16),
28291 => conv_std_logic_vector(14410, 16),
28292 => conv_std_logic_vector(14520, 16),
28293 => conv_std_logic_vector(14630, 16),
28294 => conv_std_logic_vector(14740, 16),
28295 => conv_std_logic_vector(14850, 16),
28296 => conv_std_logic_vector(14960, 16),
28297 => conv_std_logic_vector(15070, 16),
28298 => conv_std_logic_vector(15180, 16),
28299 => conv_std_logic_vector(15290, 16),
28300 => conv_std_logic_vector(15400, 16),
28301 => conv_std_logic_vector(15510, 16),
28302 => conv_std_logic_vector(15620, 16),
28303 => conv_std_logic_vector(15730, 16),
28304 => conv_std_logic_vector(15840, 16),
28305 => conv_std_logic_vector(15950, 16),
28306 => conv_std_logic_vector(16060, 16),
28307 => conv_std_logic_vector(16170, 16),
28308 => conv_std_logic_vector(16280, 16),
28309 => conv_std_logic_vector(16390, 16),
28310 => conv_std_logic_vector(16500, 16),
28311 => conv_std_logic_vector(16610, 16),
28312 => conv_std_logic_vector(16720, 16),
28313 => conv_std_logic_vector(16830, 16),
28314 => conv_std_logic_vector(16940, 16),
28315 => conv_std_logic_vector(17050, 16),
28316 => conv_std_logic_vector(17160, 16),
28317 => conv_std_logic_vector(17270, 16),
28318 => conv_std_logic_vector(17380, 16),
28319 => conv_std_logic_vector(17490, 16),
28320 => conv_std_logic_vector(17600, 16),
28321 => conv_std_logic_vector(17710, 16),
28322 => conv_std_logic_vector(17820, 16),
28323 => conv_std_logic_vector(17930, 16),
28324 => conv_std_logic_vector(18040, 16),
28325 => conv_std_logic_vector(18150, 16),
28326 => conv_std_logic_vector(18260, 16),
28327 => conv_std_logic_vector(18370, 16),
28328 => conv_std_logic_vector(18480, 16),
28329 => conv_std_logic_vector(18590, 16),
28330 => conv_std_logic_vector(18700, 16),
28331 => conv_std_logic_vector(18810, 16),
28332 => conv_std_logic_vector(18920, 16),
28333 => conv_std_logic_vector(19030, 16),
28334 => conv_std_logic_vector(19140, 16),
28335 => conv_std_logic_vector(19250, 16),
28336 => conv_std_logic_vector(19360, 16),
28337 => conv_std_logic_vector(19470, 16),
28338 => conv_std_logic_vector(19580, 16),
28339 => conv_std_logic_vector(19690, 16),
28340 => conv_std_logic_vector(19800, 16),
28341 => conv_std_logic_vector(19910, 16),
28342 => conv_std_logic_vector(20020, 16),
28343 => conv_std_logic_vector(20130, 16),
28344 => conv_std_logic_vector(20240, 16),
28345 => conv_std_logic_vector(20350, 16),
28346 => conv_std_logic_vector(20460, 16),
28347 => conv_std_logic_vector(20570, 16),
28348 => conv_std_logic_vector(20680, 16),
28349 => conv_std_logic_vector(20790, 16),
28350 => conv_std_logic_vector(20900, 16),
28351 => conv_std_logic_vector(21010, 16),
28352 => conv_std_logic_vector(21120, 16),
28353 => conv_std_logic_vector(21230, 16),
28354 => conv_std_logic_vector(21340, 16),
28355 => conv_std_logic_vector(21450, 16),
28356 => conv_std_logic_vector(21560, 16),
28357 => conv_std_logic_vector(21670, 16),
28358 => conv_std_logic_vector(21780, 16),
28359 => conv_std_logic_vector(21890, 16),
28360 => conv_std_logic_vector(22000, 16),
28361 => conv_std_logic_vector(22110, 16),
28362 => conv_std_logic_vector(22220, 16),
28363 => conv_std_logic_vector(22330, 16),
28364 => conv_std_logic_vector(22440, 16),
28365 => conv_std_logic_vector(22550, 16),
28366 => conv_std_logic_vector(22660, 16),
28367 => conv_std_logic_vector(22770, 16),
28368 => conv_std_logic_vector(22880, 16),
28369 => conv_std_logic_vector(22990, 16),
28370 => conv_std_logic_vector(23100, 16),
28371 => conv_std_logic_vector(23210, 16),
28372 => conv_std_logic_vector(23320, 16),
28373 => conv_std_logic_vector(23430, 16),
28374 => conv_std_logic_vector(23540, 16),
28375 => conv_std_logic_vector(23650, 16),
28376 => conv_std_logic_vector(23760, 16),
28377 => conv_std_logic_vector(23870, 16),
28378 => conv_std_logic_vector(23980, 16),
28379 => conv_std_logic_vector(24090, 16),
28380 => conv_std_logic_vector(24200, 16),
28381 => conv_std_logic_vector(24310, 16),
28382 => conv_std_logic_vector(24420, 16),
28383 => conv_std_logic_vector(24530, 16),
28384 => conv_std_logic_vector(24640, 16),
28385 => conv_std_logic_vector(24750, 16),
28386 => conv_std_logic_vector(24860, 16),
28387 => conv_std_logic_vector(24970, 16),
28388 => conv_std_logic_vector(25080, 16),
28389 => conv_std_logic_vector(25190, 16),
28390 => conv_std_logic_vector(25300, 16),
28391 => conv_std_logic_vector(25410, 16),
28392 => conv_std_logic_vector(25520, 16),
28393 => conv_std_logic_vector(25630, 16),
28394 => conv_std_logic_vector(25740, 16),
28395 => conv_std_logic_vector(25850, 16),
28396 => conv_std_logic_vector(25960, 16),
28397 => conv_std_logic_vector(26070, 16),
28398 => conv_std_logic_vector(26180, 16),
28399 => conv_std_logic_vector(26290, 16),
28400 => conv_std_logic_vector(26400, 16),
28401 => conv_std_logic_vector(26510, 16),
28402 => conv_std_logic_vector(26620, 16),
28403 => conv_std_logic_vector(26730, 16),
28404 => conv_std_logic_vector(26840, 16),
28405 => conv_std_logic_vector(26950, 16),
28406 => conv_std_logic_vector(27060, 16),
28407 => conv_std_logic_vector(27170, 16),
28408 => conv_std_logic_vector(27280, 16),
28409 => conv_std_logic_vector(27390, 16),
28410 => conv_std_logic_vector(27500, 16),
28411 => conv_std_logic_vector(27610, 16),
28412 => conv_std_logic_vector(27720, 16),
28413 => conv_std_logic_vector(27830, 16),
28414 => conv_std_logic_vector(27940, 16),
28415 => conv_std_logic_vector(28050, 16),
28416 => conv_std_logic_vector(0, 16),
28417 => conv_std_logic_vector(111, 16),
28418 => conv_std_logic_vector(222, 16),
28419 => conv_std_logic_vector(333, 16),
28420 => conv_std_logic_vector(444, 16),
28421 => conv_std_logic_vector(555, 16),
28422 => conv_std_logic_vector(666, 16),
28423 => conv_std_logic_vector(777, 16),
28424 => conv_std_logic_vector(888, 16),
28425 => conv_std_logic_vector(999, 16),
28426 => conv_std_logic_vector(1110, 16),
28427 => conv_std_logic_vector(1221, 16),
28428 => conv_std_logic_vector(1332, 16),
28429 => conv_std_logic_vector(1443, 16),
28430 => conv_std_logic_vector(1554, 16),
28431 => conv_std_logic_vector(1665, 16),
28432 => conv_std_logic_vector(1776, 16),
28433 => conv_std_logic_vector(1887, 16),
28434 => conv_std_logic_vector(1998, 16),
28435 => conv_std_logic_vector(2109, 16),
28436 => conv_std_logic_vector(2220, 16),
28437 => conv_std_logic_vector(2331, 16),
28438 => conv_std_logic_vector(2442, 16),
28439 => conv_std_logic_vector(2553, 16),
28440 => conv_std_logic_vector(2664, 16),
28441 => conv_std_logic_vector(2775, 16),
28442 => conv_std_logic_vector(2886, 16),
28443 => conv_std_logic_vector(2997, 16),
28444 => conv_std_logic_vector(3108, 16),
28445 => conv_std_logic_vector(3219, 16),
28446 => conv_std_logic_vector(3330, 16),
28447 => conv_std_logic_vector(3441, 16),
28448 => conv_std_logic_vector(3552, 16),
28449 => conv_std_logic_vector(3663, 16),
28450 => conv_std_logic_vector(3774, 16),
28451 => conv_std_logic_vector(3885, 16),
28452 => conv_std_logic_vector(3996, 16),
28453 => conv_std_logic_vector(4107, 16),
28454 => conv_std_logic_vector(4218, 16),
28455 => conv_std_logic_vector(4329, 16),
28456 => conv_std_logic_vector(4440, 16),
28457 => conv_std_logic_vector(4551, 16),
28458 => conv_std_logic_vector(4662, 16),
28459 => conv_std_logic_vector(4773, 16),
28460 => conv_std_logic_vector(4884, 16),
28461 => conv_std_logic_vector(4995, 16),
28462 => conv_std_logic_vector(5106, 16),
28463 => conv_std_logic_vector(5217, 16),
28464 => conv_std_logic_vector(5328, 16),
28465 => conv_std_logic_vector(5439, 16),
28466 => conv_std_logic_vector(5550, 16),
28467 => conv_std_logic_vector(5661, 16),
28468 => conv_std_logic_vector(5772, 16),
28469 => conv_std_logic_vector(5883, 16),
28470 => conv_std_logic_vector(5994, 16),
28471 => conv_std_logic_vector(6105, 16),
28472 => conv_std_logic_vector(6216, 16),
28473 => conv_std_logic_vector(6327, 16),
28474 => conv_std_logic_vector(6438, 16),
28475 => conv_std_logic_vector(6549, 16),
28476 => conv_std_logic_vector(6660, 16),
28477 => conv_std_logic_vector(6771, 16),
28478 => conv_std_logic_vector(6882, 16),
28479 => conv_std_logic_vector(6993, 16),
28480 => conv_std_logic_vector(7104, 16),
28481 => conv_std_logic_vector(7215, 16),
28482 => conv_std_logic_vector(7326, 16),
28483 => conv_std_logic_vector(7437, 16),
28484 => conv_std_logic_vector(7548, 16),
28485 => conv_std_logic_vector(7659, 16),
28486 => conv_std_logic_vector(7770, 16),
28487 => conv_std_logic_vector(7881, 16),
28488 => conv_std_logic_vector(7992, 16),
28489 => conv_std_logic_vector(8103, 16),
28490 => conv_std_logic_vector(8214, 16),
28491 => conv_std_logic_vector(8325, 16),
28492 => conv_std_logic_vector(8436, 16),
28493 => conv_std_logic_vector(8547, 16),
28494 => conv_std_logic_vector(8658, 16),
28495 => conv_std_logic_vector(8769, 16),
28496 => conv_std_logic_vector(8880, 16),
28497 => conv_std_logic_vector(8991, 16),
28498 => conv_std_logic_vector(9102, 16),
28499 => conv_std_logic_vector(9213, 16),
28500 => conv_std_logic_vector(9324, 16),
28501 => conv_std_logic_vector(9435, 16),
28502 => conv_std_logic_vector(9546, 16),
28503 => conv_std_logic_vector(9657, 16),
28504 => conv_std_logic_vector(9768, 16),
28505 => conv_std_logic_vector(9879, 16),
28506 => conv_std_logic_vector(9990, 16),
28507 => conv_std_logic_vector(10101, 16),
28508 => conv_std_logic_vector(10212, 16),
28509 => conv_std_logic_vector(10323, 16),
28510 => conv_std_logic_vector(10434, 16),
28511 => conv_std_logic_vector(10545, 16),
28512 => conv_std_logic_vector(10656, 16),
28513 => conv_std_logic_vector(10767, 16),
28514 => conv_std_logic_vector(10878, 16),
28515 => conv_std_logic_vector(10989, 16),
28516 => conv_std_logic_vector(11100, 16),
28517 => conv_std_logic_vector(11211, 16),
28518 => conv_std_logic_vector(11322, 16),
28519 => conv_std_logic_vector(11433, 16),
28520 => conv_std_logic_vector(11544, 16),
28521 => conv_std_logic_vector(11655, 16),
28522 => conv_std_logic_vector(11766, 16),
28523 => conv_std_logic_vector(11877, 16),
28524 => conv_std_logic_vector(11988, 16),
28525 => conv_std_logic_vector(12099, 16),
28526 => conv_std_logic_vector(12210, 16),
28527 => conv_std_logic_vector(12321, 16),
28528 => conv_std_logic_vector(12432, 16),
28529 => conv_std_logic_vector(12543, 16),
28530 => conv_std_logic_vector(12654, 16),
28531 => conv_std_logic_vector(12765, 16),
28532 => conv_std_logic_vector(12876, 16),
28533 => conv_std_logic_vector(12987, 16),
28534 => conv_std_logic_vector(13098, 16),
28535 => conv_std_logic_vector(13209, 16),
28536 => conv_std_logic_vector(13320, 16),
28537 => conv_std_logic_vector(13431, 16),
28538 => conv_std_logic_vector(13542, 16),
28539 => conv_std_logic_vector(13653, 16),
28540 => conv_std_logic_vector(13764, 16),
28541 => conv_std_logic_vector(13875, 16),
28542 => conv_std_logic_vector(13986, 16),
28543 => conv_std_logic_vector(14097, 16),
28544 => conv_std_logic_vector(14208, 16),
28545 => conv_std_logic_vector(14319, 16),
28546 => conv_std_logic_vector(14430, 16),
28547 => conv_std_logic_vector(14541, 16),
28548 => conv_std_logic_vector(14652, 16),
28549 => conv_std_logic_vector(14763, 16),
28550 => conv_std_logic_vector(14874, 16),
28551 => conv_std_logic_vector(14985, 16),
28552 => conv_std_logic_vector(15096, 16),
28553 => conv_std_logic_vector(15207, 16),
28554 => conv_std_logic_vector(15318, 16),
28555 => conv_std_logic_vector(15429, 16),
28556 => conv_std_logic_vector(15540, 16),
28557 => conv_std_logic_vector(15651, 16),
28558 => conv_std_logic_vector(15762, 16),
28559 => conv_std_logic_vector(15873, 16),
28560 => conv_std_logic_vector(15984, 16),
28561 => conv_std_logic_vector(16095, 16),
28562 => conv_std_logic_vector(16206, 16),
28563 => conv_std_logic_vector(16317, 16),
28564 => conv_std_logic_vector(16428, 16),
28565 => conv_std_logic_vector(16539, 16),
28566 => conv_std_logic_vector(16650, 16),
28567 => conv_std_logic_vector(16761, 16),
28568 => conv_std_logic_vector(16872, 16),
28569 => conv_std_logic_vector(16983, 16),
28570 => conv_std_logic_vector(17094, 16),
28571 => conv_std_logic_vector(17205, 16),
28572 => conv_std_logic_vector(17316, 16),
28573 => conv_std_logic_vector(17427, 16),
28574 => conv_std_logic_vector(17538, 16),
28575 => conv_std_logic_vector(17649, 16),
28576 => conv_std_logic_vector(17760, 16),
28577 => conv_std_logic_vector(17871, 16),
28578 => conv_std_logic_vector(17982, 16),
28579 => conv_std_logic_vector(18093, 16),
28580 => conv_std_logic_vector(18204, 16),
28581 => conv_std_logic_vector(18315, 16),
28582 => conv_std_logic_vector(18426, 16),
28583 => conv_std_logic_vector(18537, 16),
28584 => conv_std_logic_vector(18648, 16),
28585 => conv_std_logic_vector(18759, 16),
28586 => conv_std_logic_vector(18870, 16),
28587 => conv_std_logic_vector(18981, 16),
28588 => conv_std_logic_vector(19092, 16),
28589 => conv_std_logic_vector(19203, 16),
28590 => conv_std_logic_vector(19314, 16),
28591 => conv_std_logic_vector(19425, 16),
28592 => conv_std_logic_vector(19536, 16),
28593 => conv_std_logic_vector(19647, 16),
28594 => conv_std_logic_vector(19758, 16),
28595 => conv_std_logic_vector(19869, 16),
28596 => conv_std_logic_vector(19980, 16),
28597 => conv_std_logic_vector(20091, 16),
28598 => conv_std_logic_vector(20202, 16),
28599 => conv_std_logic_vector(20313, 16),
28600 => conv_std_logic_vector(20424, 16),
28601 => conv_std_logic_vector(20535, 16),
28602 => conv_std_logic_vector(20646, 16),
28603 => conv_std_logic_vector(20757, 16),
28604 => conv_std_logic_vector(20868, 16),
28605 => conv_std_logic_vector(20979, 16),
28606 => conv_std_logic_vector(21090, 16),
28607 => conv_std_logic_vector(21201, 16),
28608 => conv_std_logic_vector(21312, 16),
28609 => conv_std_logic_vector(21423, 16),
28610 => conv_std_logic_vector(21534, 16),
28611 => conv_std_logic_vector(21645, 16),
28612 => conv_std_logic_vector(21756, 16),
28613 => conv_std_logic_vector(21867, 16),
28614 => conv_std_logic_vector(21978, 16),
28615 => conv_std_logic_vector(22089, 16),
28616 => conv_std_logic_vector(22200, 16),
28617 => conv_std_logic_vector(22311, 16),
28618 => conv_std_logic_vector(22422, 16),
28619 => conv_std_logic_vector(22533, 16),
28620 => conv_std_logic_vector(22644, 16),
28621 => conv_std_logic_vector(22755, 16),
28622 => conv_std_logic_vector(22866, 16),
28623 => conv_std_logic_vector(22977, 16),
28624 => conv_std_logic_vector(23088, 16),
28625 => conv_std_logic_vector(23199, 16),
28626 => conv_std_logic_vector(23310, 16),
28627 => conv_std_logic_vector(23421, 16),
28628 => conv_std_logic_vector(23532, 16),
28629 => conv_std_logic_vector(23643, 16),
28630 => conv_std_logic_vector(23754, 16),
28631 => conv_std_logic_vector(23865, 16),
28632 => conv_std_logic_vector(23976, 16),
28633 => conv_std_logic_vector(24087, 16),
28634 => conv_std_logic_vector(24198, 16),
28635 => conv_std_logic_vector(24309, 16),
28636 => conv_std_logic_vector(24420, 16),
28637 => conv_std_logic_vector(24531, 16),
28638 => conv_std_logic_vector(24642, 16),
28639 => conv_std_logic_vector(24753, 16),
28640 => conv_std_logic_vector(24864, 16),
28641 => conv_std_logic_vector(24975, 16),
28642 => conv_std_logic_vector(25086, 16),
28643 => conv_std_logic_vector(25197, 16),
28644 => conv_std_logic_vector(25308, 16),
28645 => conv_std_logic_vector(25419, 16),
28646 => conv_std_logic_vector(25530, 16),
28647 => conv_std_logic_vector(25641, 16),
28648 => conv_std_logic_vector(25752, 16),
28649 => conv_std_logic_vector(25863, 16),
28650 => conv_std_logic_vector(25974, 16),
28651 => conv_std_logic_vector(26085, 16),
28652 => conv_std_logic_vector(26196, 16),
28653 => conv_std_logic_vector(26307, 16),
28654 => conv_std_logic_vector(26418, 16),
28655 => conv_std_logic_vector(26529, 16),
28656 => conv_std_logic_vector(26640, 16),
28657 => conv_std_logic_vector(26751, 16),
28658 => conv_std_logic_vector(26862, 16),
28659 => conv_std_logic_vector(26973, 16),
28660 => conv_std_logic_vector(27084, 16),
28661 => conv_std_logic_vector(27195, 16),
28662 => conv_std_logic_vector(27306, 16),
28663 => conv_std_logic_vector(27417, 16),
28664 => conv_std_logic_vector(27528, 16),
28665 => conv_std_logic_vector(27639, 16),
28666 => conv_std_logic_vector(27750, 16),
28667 => conv_std_logic_vector(27861, 16),
28668 => conv_std_logic_vector(27972, 16),
28669 => conv_std_logic_vector(28083, 16),
28670 => conv_std_logic_vector(28194, 16),
28671 => conv_std_logic_vector(28305, 16),
28672 => conv_std_logic_vector(0, 16),
28673 => conv_std_logic_vector(112, 16),
28674 => conv_std_logic_vector(224, 16),
28675 => conv_std_logic_vector(336, 16),
28676 => conv_std_logic_vector(448, 16),
28677 => conv_std_logic_vector(560, 16),
28678 => conv_std_logic_vector(672, 16),
28679 => conv_std_logic_vector(784, 16),
28680 => conv_std_logic_vector(896, 16),
28681 => conv_std_logic_vector(1008, 16),
28682 => conv_std_logic_vector(1120, 16),
28683 => conv_std_logic_vector(1232, 16),
28684 => conv_std_logic_vector(1344, 16),
28685 => conv_std_logic_vector(1456, 16),
28686 => conv_std_logic_vector(1568, 16),
28687 => conv_std_logic_vector(1680, 16),
28688 => conv_std_logic_vector(1792, 16),
28689 => conv_std_logic_vector(1904, 16),
28690 => conv_std_logic_vector(2016, 16),
28691 => conv_std_logic_vector(2128, 16),
28692 => conv_std_logic_vector(2240, 16),
28693 => conv_std_logic_vector(2352, 16),
28694 => conv_std_logic_vector(2464, 16),
28695 => conv_std_logic_vector(2576, 16),
28696 => conv_std_logic_vector(2688, 16),
28697 => conv_std_logic_vector(2800, 16),
28698 => conv_std_logic_vector(2912, 16),
28699 => conv_std_logic_vector(3024, 16),
28700 => conv_std_logic_vector(3136, 16),
28701 => conv_std_logic_vector(3248, 16),
28702 => conv_std_logic_vector(3360, 16),
28703 => conv_std_logic_vector(3472, 16),
28704 => conv_std_logic_vector(3584, 16),
28705 => conv_std_logic_vector(3696, 16),
28706 => conv_std_logic_vector(3808, 16),
28707 => conv_std_logic_vector(3920, 16),
28708 => conv_std_logic_vector(4032, 16),
28709 => conv_std_logic_vector(4144, 16),
28710 => conv_std_logic_vector(4256, 16),
28711 => conv_std_logic_vector(4368, 16),
28712 => conv_std_logic_vector(4480, 16),
28713 => conv_std_logic_vector(4592, 16),
28714 => conv_std_logic_vector(4704, 16),
28715 => conv_std_logic_vector(4816, 16),
28716 => conv_std_logic_vector(4928, 16),
28717 => conv_std_logic_vector(5040, 16),
28718 => conv_std_logic_vector(5152, 16),
28719 => conv_std_logic_vector(5264, 16),
28720 => conv_std_logic_vector(5376, 16),
28721 => conv_std_logic_vector(5488, 16),
28722 => conv_std_logic_vector(5600, 16),
28723 => conv_std_logic_vector(5712, 16),
28724 => conv_std_logic_vector(5824, 16),
28725 => conv_std_logic_vector(5936, 16),
28726 => conv_std_logic_vector(6048, 16),
28727 => conv_std_logic_vector(6160, 16),
28728 => conv_std_logic_vector(6272, 16),
28729 => conv_std_logic_vector(6384, 16),
28730 => conv_std_logic_vector(6496, 16),
28731 => conv_std_logic_vector(6608, 16),
28732 => conv_std_logic_vector(6720, 16),
28733 => conv_std_logic_vector(6832, 16),
28734 => conv_std_logic_vector(6944, 16),
28735 => conv_std_logic_vector(7056, 16),
28736 => conv_std_logic_vector(7168, 16),
28737 => conv_std_logic_vector(7280, 16),
28738 => conv_std_logic_vector(7392, 16),
28739 => conv_std_logic_vector(7504, 16),
28740 => conv_std_logic_vector(7616, 16),
28741 => conv_std_logic_vector(7728, 16),
28742 => conv_std_logic_vector(7840, 16),
28743 => conv_std_logic_vector(7952, 16),
28744 => conv_std_logic_vector(8064, 16),
28745 => conv_std_logic_vector(8176, 16),
28746 => conv_std_logic_vector(8288, 16),
28747 => conv_std_logic_vector(8400, 16),
28748 => conv_std_logic_vector(8512, 16),
28749 => conv_std_logic_vector(8624, 16),
28750 => conv_std_logic_vector(8736, 16),
28751 => conv_std_logic_vector(8848, 16),
28752 => conv_std_logic_vector(8960, 16),
28753 => conv_std_logic_vector(9072, 16),
28754 => conv_std_logic_vector(9184, 16),
28755 => conv_std_logic_vector(9296, 16),
28756 => conv_std_logic_vector(9408, 16),
28757 => conv_std_logic_vector(9520, 16),
28758 => conv_std_logic_vector(9632, 16),
28759 => conv_std_logic_vector(9744, 16),
28760 => conv_std_logic_vector(9856, 16),
28761 => conv_std_logic_vector(9968, 16),
28762 => conv_std_logic_vector(10080, 16),
28763 => conv_std_logic_vector(10192, 16),
28764 => conv_std_logic_vector(10304, 16),
28765 => conv_std_logic_vector(10416, 16),
28766 => conv_std_logic_vector(10528, 16),
28767 => conv_std_logic_vector(10640, 16),
28768 => conv_std_logic_vector(10752, 16),
28769 => conv_std_logic_vector(10864, 16),
28770 => conv_std_logic_vector(10976, 16),
28771 => conv_std_logic_vector(11088, 16),
28772 => conv_std_logic_vector(11200, 16),
28773 => conv_std_logic_vector(11312, 16),
28774 => conv_std_logic_vector(11424, 16),
28775 => conv_std_logic_vector(11536, 16),
28776 => conv_std_logic_vector(11648, 16),
28777 => conv_std_logic_vector(11760, 16),
28778 => conv_std_logic_vector(11872, 16),
28779 => conv_std_logic_vector(11984, 16),
28780 => conv_std_logic_vector(12096, 16),
28781 => conv_std_logic_vector(12208, 16),
28782 => conv_std_logic_vector(12320, 16),
28783 => conv_std_logic_vector(12432, 16),
28784 => conv_std_logic_vector(12544, 16),
28785 => conv_std_logic_vector(12656, 16),
28786 => conv_std_logic_vector(12768, 16),
28787 => conv_std_logic_vector(12880, 16),
28788 => conv_std_logic_vector(12992, 16),
28789 => conv_std_logic_vector(13104, 16),
28790 => conv_std_logic_vector(13216, 16),
28791 => conv_std_logic_vector(13328, 16),
28792 => conv_std_logic_vector(13440, 16),
28793 => conv_std_logic_vector(13552, 16),
28794 => conv_std_logic_vector(13664, 16),
28795 => conv_std_logic_vector(13776, 16),
28796 => conv_std_logic_vector(13888, 16),
28797 => conv_std_logic_vector(14000, 16),
28798 => conv_std_logic_vector(14112, 16),
28799 => conv_std_logic_vector(14224, 16),
28800 => conv_std_logic_vector(14336, 16),
28801 => conv_std_logic_vector(14448, 16),
28802 => conv_std_logic_vector(14560, 16),
28803 => conv_std_logic_vector(14672, 16),
28804 => conv_std_logic_vector(14784, 16),
28805 => conv_std_logic_vector(14896, 16),
28806 => conv_std_logic_vector(15008, 16),
28807 => conv_std_logic_vector(15120, 16),
28808 => conv_std_logic_vector(15232, 16),
28809 => conv_std_logic_vector(15344, 16),
28810 => conv_std_logic_vector(15456, 16),
28811 => conv_std_logic_vector(15568, 16),
28812 => conv_std_logic_vector(15680, 16),
28813 => conv_std_logic_vector(15792, 16),
28814 => conv_std_logic_vector(15904, 16),
28815 => conv_std_logic_vector(16016, 16),
28816 => conv_std_logic_vector(16128, 16),
28817 => conv_std_logic_vector(16240, 16),
28818 => conv_std_logic_vector(16352, 16),
28819 => conv_std_logic_vector(16464, 16),
28820 => conv_std_logic_vector(16576, 16),
28821 => conv_std_logic_vector(16688, 16),
28822 => conv_std_logic_vector(16800, 16),
28823 => conv_std_logic_vector(16912, 16),
28824 => conv_std_logic_vector(17024, 16),
28825 => conv_std_logic_vector(17136, 16),
28826 => conv_std_logic_vector(17248, 16),
28827 => conv_std_logic_vector(17360, 16),
28828 => conv_std_logic_vector(17472, 16),
28829 => conv_std_logic_vector(17584, 16),
28830 => conv_std_logic_vector(17696, 16),
28831 => conv_std_logic_vector(17808, 16),
28832 => conv_std_logic_vector(17920, 16),
28833 => conv_std_logic_vector(18032, 16),
28834 => conv_std_logic_vector(18144, 16),
28835 => conv_std_logic_vector(18256, 16),
28836 => conv_std_logic_vector(18368, 16),
28837 => conv_std_logic_vector(18480, 16),
28838 => conv_std_logic_vector(18592, 16),
28839 => conv_std_logic_vector(18704, 16),
28840 => conv_std_logic_vector(18816, 16),
28841 => conv_std_logic_vector(18928, 16),
28842 => conv_std_logic_vector(19040, 16),
28843 => conv_std_logic_vector(19152, 16),
28844 => conv_std_logic_vector(19264, 16),
28845 => conv_std_logic_vector(19376, 16),
28846 => conv_std_logic_vector(19488, 16),
28847 => conv_std_logic_vector(19600, 16),
28848 => conv_std_logic_vector(19712, 16),
28849 => conv_std_logic_vector(19824, 16),
28850 => conv_std_logic_vector(19936, 16),
28851 => conv_std_logic_vector(20048, 16),
28852 => conv_std_logic_vector(20160, 16),
28853 => conv_std_logic_vector(20272, 16),
28854 => conv_std_logic_vector(20384, 16),
28855 => conv_std_logic_vector(20496, 16),
28856 => conv_std_logic_vector(20608, 16),
28857 => conv_std_logic_vector(20720, 16),
28858 => conv_std_logic_vector(20832, 16),
28859 => conv_std_logic_vector(20944, 16),
28860 => conv_std_logic_vector(21056, 16),
28861 => conv_std_logic_vector(21168, 16),
28862 => conv_std_logic_vector(21280, 16),
28863 => conv_std_logic_vector(21392, 16),
28864 => conv_std_logic_vector(21504, 16),
28865 => conv_std_logic_vector(21616, 16),
28866 => conv_std_logic_vector(21728, 16),
28867 => conv_std_logic_vector(21840, 16),
28868 => conv_std_logic_vector(21952, 16),
28869 => conv_std_logic_vector(22064, 16),
28870 => conv_std_logic_vector(22176, 16),
28871 => conv_std_logic_vector(22288, 16),
28872 => conv_std_logic_vector(22400, 16),
28873 => conv_std_logic_vector(22512, 16),
28874 => conv_std_logic_vector(22624, 16),
28875 => conv_std_logic_vector(22736, 16),
28876 => conv_std_logic_vector(22848, 16),
28877 => conv_std_logic_vector(22960, 16),
28878 => conv_std_logic_vector(23072, 16),
28879 => conv_std_logic_vector(23184, 16),
28880 => conv_std_logic_vector(23296, 16),
28881 => conv_std_logic_vector(23408, 16),
28882 => conv_std_logic_vector(23520, 16),
28883 => conv_std_logic_vector(23632, 16),
28884 => conv_std_logic_vector(23744, 16),
28885 => conv_std_logic_vector(23856, 16),
28886 => conv_std_logic_vector(23968, 16),
28887 => conv_std_logic_vector(24080, 16),
28888 => conv_std_logic_vector(24192, 16),
28889 => conv_std_logic_vector(24304, 16),
28890 => conv_std_logic_vector(24416, 16),
28891 => conv_std_logic_vector(24528, 16),
28892 => conv_std_logic_vector(24640, 16),
28893 => conv_std_logic_vector(24752, 16),
28894 => conv_std_logic_vector(24864, 16),
28895 => conv_std_logic_vector(24976, 16),
28896 => conv_std_logic_vector(25088, 16),
28897 => conv_std_logic_vector(25200, 16),
28898 => conv_std_logic_vector(25312, 16),
28899 => conv_std_logic_vector(25424, 16),
28900 => conv_std_logic_vector(25536, 16),
28901 => conv_std_logic_vector(25648, 16),
28902 => conv_std_logic_vector(25760, 16),
28903 => conv_std_logic_vector(25872, 16),
28904 => conv_std_logic_vector(25984, 16),
28905 => conv_std_logic_vector(26096, 16),
28906 => conv_std_logic_vector(26208, 16),
28907 => conv_std_logic_vector(26320, 16),
28908 => conv_std_logic_vector(26432, 16),
28909 => conv_std_logic_vector(26544, 16),
28910 => conv_std_logic_vector(26656, 16),
28911 => conv_std_logic_vector(26768, 16),
28912 => conv_std_logic_vector(26880, 16),
28913 => conv_std_logic_vector(26992, 16),
28914 => conv_std_logic_vector(27104, 16),
28915 => conv_std_logic_vector(27216, 16),
28916 => conv_std_logic_vector(27328, 16),
28917 => conv_std_logic_vector(27440, 16),
28918 => conv_std_logic_vector(27552, 16),
28919 => conv_std_logic_vector(27664, 16),
28920 => conv_std_logic_vector(27776, 16),
28921 => conv_std_logic_vector(27888, 16),
28922 => conv_std_logic_vector(28000, 16),
28923 => conv_std_logic_vector(28112, 16),
28924 => conv_std_logic_vector(28224, 16),
28925 => conv_std_logic_vector(28336, 16),
28926 => conv_std_logic_vector(28448, 16),
28927 => conv_std_logic_vector(28560, 16),
28928 => conv_std_logic_vector(0, 16),
28929 => conv_std_logic_vector(113, 16),
28930 => conv_std_logic_vector(226, 16),
28931 => conv_std_logic_vector(339, 16),
28932 => conv_std_logic_vector(452, 16),
28933 => conv_std_logic_vector(565, 16),
28934 => conv_std_logic_vector(678, 16),
28935 => conv_std_logic_vector(791, 16),
28936 => conv_std_logic_vector(904, 16),
28937 => conv_std_logic_vector(1017, 16),
28938 => conv_std_logic_vector(1130, 16),
28939 => conv_std_logic_vector(1243, 16),
28940 => conv_std_logic_vector(1356, 16),
28941 => conv_std_logic_vector(1469, 16),
28942 => conv_std_logic_vector(1582, 16),
28943 => conv_std_logic_vector(1695, 16),
28944 => conv_std_logic_vector(1808, 16),
28945 => conv_std_logic_vector(1921, 16),
28946 => conv_std_logic_vector(2034, 16),
28947 => conv_std_logic_vector(2147, 16),
28948 => conv_std_logic_vector(2260, 16),
28949 => conv_std_logic_vector(2373, 16),
28950 => conv_std_logic_vector(2486, 16),
28951 => conv_std_logic_vector(2599, 16),
28952 => conv_std_logic_vector(2712, 16),
28953 => conv_std_logic_vector(2825, 16),
28954 => conv_std_logic_vector(2938, 16),
28955 => conv_std_logic_vector(3051, 16),
28956 => conv_std_logic_vector(3164, 16),
28957 => conv_std_logic_vector(3277, 16),
28958 => conv_std_logic_vector(3390, 16),
28959 => conv_std_logic_vector(3503, 16),
28960 => conv_std_logic_vector(3616, 16),
28961 => conv_std_logic_vector(3729, 16),
28962 => conv_std_logic_vector(3842, 16),
28963 => conv_std_logic_vector(3955, 16),
28964 => conv_std_logic_vector(4068, 16),
28965 => conv_std_logic_vector(4181, 16),
28966 => conv_std_logic_vector(4294, 16),
28967 => conv_std_logic_vector(4407, 16),
28968 => conv_std_logic_vector(4520, 16),
28969 => conv_std_logic_vector(4633, 16),
28970 => conv_std_logic_vector(4746, 16),
28971 => conv_std_logic_vector(4859, 16),
28972 => conv_std_logic_vector(4972, 16),
28973 => conv_std_logic_vector(5085, 16),
28974 => conv_std_logic_vector(5198, 16),
28975 => conv_std_logic_vector(5311, 16),
28976 => conv_std_logic_vector(5424, 16),
28977 => conv_std_logic_vector(5537, 16),
28978 => conv_std_logic_vector(5650, 16),
28979 => conv_std_logic_vector(5763, 16),
28980 => conv_std_logic_vector(5876, 16),
28981 => conv_std_logic_vector(5989, 16),
28982 => conv_std_logic_vector(6102, 16),
28983 => conv_std_logic_vector(6215, 16),
28984 => conv_std_logic_vector(6328, 16),
28985 => conv_std_logic_vector(6441, 16),
28986 => conv_std_logic_vector(6554, 16),
28987 => conv_std_logic_vector(6667, 16),
28988 => conv_std_logic_vector(6780, 16),
28989 => conv_std_logic_vector(6893, 16),
28990 => conv_std_logic_vector(7006, 16),
28991 => conv_std_logic_vector(7119, 16),
28992 => conv_std_logic_vector(7232, 16),
28993 => conv_std_logic_vector(7345, 16),
28994 => conv_std_logic_vector(7458, 16),
28995 => conv_std_logic_vector(7571, 16),
28996 => conv_std_logic_vector(7684, 16),
28997 => conv_std_logic_vector(7797, 16),
28998 => conv_std_logic_vector(7910, 16),
28999 => conv_std_logic_vector(8023, 16),
29000 => conv_std_logic_vector(8136, 16),
29001 => conv_std_logic_vector(8249, 16),
29002 => conv_std_logic_vector(8362, 16),
29003 => conv_std_logic_vector(8475, 16),
29004 => conv_std_logic_vector(8588, 16),
29005 => conv_std_logic_vector(8701, 16),
29006 => conv_std_logic_vector(8814, 16),
29007 => conv_std_logic_vector(8927, 16),
29008 => conv_std_logic_vector(9040, 16),
29009 => conv_std_logic_vector(9153, 16),
29010 => conv_std_logic_vector(9266, 16),
29011 => conv_std_logic_vector(9379, 16),
29012 => conv_std_logic_vector(9492, 16),
29013 => conv_std_logic_vector(9605, 16),
29014 => conv_std_logic_vector(9718, 16),
29015 => conv_std_logic_vector(9831, 16),
29016 => conv_std_logic_vector(9944, 16),
29017 => conv_std_logic_vector(10057, 16),
29018 => conv_std_logic_vector(10170, 16),
29019 => conv_std_logic_vector(10283, 16),
29020 => conv_std_logic_vector(10396, 16),
29021 => conv_std_logic_vector(10509, 16),
29022 => conv_std_logic_vector(10622, 16),
29023 => conv_std_logic_vector(10735, 16),
29024 => conv_std_logic_vector(10848, 16),
29025 => conv_std_logic_vector(10961, 16),
29026 => conv_std_logic_vector(11074, 16),
29027 => conv_std_logic_vector(11187, 16),
29028 => conv_std_logic_vector(11300, 16),
29029 => conv_std_logic_vector(11413, 16),
29030 => conv_std_logic_vector(11526, 16),
29031 => conv_std_logic_vector(11639, 16),
29032 => conv_std_logic_vector(11752, 16),
29033 => conv_std_logic_vector(11865, 16),
29034 => conv_std_logic_vector(11978, 16),
29035 => conv_std_logic_vector(12091, 16),
29036 => conv_std_logic_vector(12204, 16),
29037 => conv_std_logic_vector(12317, 16),
29038 => conv_std_logic_vector(12430, 16),
29039 => conv_std_logic_vector(12543, 16),
29040 => conv_std_logic_vector(12656, 16),
29041 => conv_std_logic_vector(12769, 16),
29042 => conv_std_logic_vector(12882, 16),
29043 => conv_std_logic_vector(12995, 16),
29044 => conv_std_logic_vector(13108, 16),
29045 => conv_std_logic_vector(13221, 16),
29046 => conv_std_logic_vector(13334, 16),
29047 => conv_std_logic_vector(13447, 16),
29048 => conv_std_logic_vector(13560, 16),
29049 => conv_std_logic_vector(13673, 16),
29050 => conv_std_logic_vector(13786, 16),
29051 => conv_std_logic_vector(13899, 16),
29052 => conv_std_logic_vector(14012, 16),
29053 => conv_std_logic_vector(14125, 16),
29054 => conv_std_logic_vector(14238, 16),
29055 => conv_std_logic_vector(14351, 16),
29056 => conv_std_logic_vector(14464, 16),
29057 => conv_std_logic_vector(14577, 16),
29058 => conv_std_logic_vector(14690, 16),
29059 => conv_std_logic_vector(14803, 16),
29060 => conv_std_logic_vector(14916, 16),
29061 => conv_std_logic_vector(15029, 16),
29062 => conv_std_logic_vector(15142, 16),
29063 => conv_std_logic_vector(15255, 16),
29064 => conv_std_logic_vector(15368, 16),
29065 => conv_std_logic_vector(15481, 16),
29066 => conv_std_logic_vector(15594, 16),
29067 => conv_std_logic_vector(15707, 16),
29068 => conv_std_logic_vector(15820, 16),
29069 => conv_std_logic_vector(15933, 16),
29070 => conv_std_logic_vector(16046, 16),
29071 => conv_std_logic_vector(16159, 16),
29072 => conv_std_logic_vector(16272, 16),
29073 => conv_std_logic_vector(16385, 16),
29074 => conv_std_logic_vector(16498, 16),
29075 => conv_std_logic_vector(16611, 16),
29076 => conv_std_logic_vector(16724, 16),
29077 => conv_std_logic_vector(16837, 16),
29078 => conv_std_logic_vector(16950, 16),
29079 => conv_std_logic_vector(17063, 16),
29080 => conv_std_logic_vector(17176, 16),
29081 => conv_std_logic_vector(17289, 16),
29082 => conv_std_logic_vector(17402, 16),
29083 => conv_std_logic_vector(17515, 16),
29084 => conv_std_logic_vector(17628, 16),
29085 => conv_std_logic_vector(17741, 16),
29086 => conv_std_logic_vector(17854, 16),
29087 => conv_std_logic_vector(17967, 16),
29088 => conv_std_logic_vector(18080, 16),
29089 => conv_std_logic_vector(18193, 16),
29090 => conv_std_logic_vector(18306, 16),
29091 => conv_std_logic_vector(18419, 16),
29092 => conv_std_logic_vector(18532, 16),
29093 => conv_std_logic_vector(18645, 16),
29094 => conv_std_logic_vector(18758, 16),
29095 => conv_std_logic_vector(18871, 16),
29096 => conv_std_logic_vector(18984, 16),
29097 => conv_std_logic_vector(19097, 16),
29098 => conv_std_logic_vector(19210, 16),
29099 => conv_std_logic_vector(19323, 16),
29100 => conv_std_logic_vector(19436, 16),
29101 => conv_std_logic_vector(19549, 16),
29102 => conv_std_logic_vector(19662, 16),
29103 => conv_std_logic_vector(19775, 16),
29104 => conv_std_logic_vector(19888, 16),
29105 => conv_std_logic_vector(20001, 16),
29106 => conv_std_logic_vector(20114, 16),
29107 => conv_std_logic_vector(20227, 16),
29108 => conv_std_logic_vector(20340, 16),
29109 => conv_std_logic_vector(20453, 16),
29110 => conv_std_logic_vector(20566, 16),
29111 => conv_std_logic_vector(20679, 16),
29112 => conv_std_logic_vector(20792, 16),
29113 => conv_std_logic_vector(20905, 16),
29114 => conv_std_logic_vector(21018, 16),
29115 => conv_std_logic_vector(21131, 16),
29116 => conv_std_logic_vector(21244, 16),
29117 => conv_std_logic_vector(21357, 16),
29118 => conv_std_logic_vector(21470, 16),
29119 => conv_std_logic_vector(21583, 16),
29120 => conv_std_logic_vector(21696, 16),
29121 => conv_std_logic_vector(21809, 16),
29122 => conv_std_logic_vector(21922, 16),
29123 => conv_std_logic_vector(22035, 16),
29124 => conv_std_logic_vector(22148, 16),
29125 => conv_std_logic_vector(22261, 16),
29126 => conv_std_logic_vector(22374, 16),
29127 => conv_std_logic_vector(22487, 16),
29128 => conv_std_logic_vector(22600, 16),
29129 => conv_std_logic_vector(22713, 16),
29130 => conv_std_logic_vector(22826, 16),
29131 => conv_std_logic_vector(22939, 16),
29132 => conv_std_logic_vector(23052, 16),
29133 => conv_std_logic_vector(23165, 16),
29134 => conv_std_logic_vector(23278, 16),
29135 => conv_std_logic_vector(23391, 16),
29136 => conv_std_logic_vector(23504, 16),
29137 => conv_std_logic_vector(23617, 16),
29138 => conv_std_logic_vector(23730, 16),
29139 => conv_std_logic_vector(23843, 16),
29140 => conv_std_logic_vector(23956, 16),
29141 => conv_std_logic_vector(24069, 16),
29142 => conv_std_logic_vector(24182, 16),
29143 => conv_std_logic_vector(24295, 16),
29144 => conv_std_logic_vector(24408, 16),
29145 => conv_std_logic_vector(24521, 16),
29146 => conv_std_logic_vector(24634, 16),
29147 => conv_std_logic_vector(24747, 16),
29148 => conv_std_logic_vector(24860, 16),
29149 => conv_std_logic_vector(24973, 16),
29150 => conv_std_logic_vector(25086, 16),
29151 => conv_std_logic_vector(25199, 16),
29152 => conv_std_logic_vector(25312, 16),
29153 => conv_std_logic_vector(25425, 16),
29154 => conv_std_logic_vector(25538, 16),
29155 => conv_std_logic_vector(25651, 16),
29156 => conv_std_logic_vector(25764, 16),
29157 => conv_std_logic_vector(25877, 16),
29158 => conv_std_logic_vector(25990, 16),
29159 => conv_std_logic_vector(26103, 16),
29160 => conv_std_logic_vector(26216, 16),
29161 => conv_std_logic_vector(26329, 16),
29162 => conv_std_logic_vector(26442, 16),
29163 => conv_std_logic_vector(26555, 16),
29164 => conv_std_logic_vector(26668, 16),
29165 => conv_std_logic_vector(26781, 16),
29166 => conv_std_logic_vector(26894, 16),
29167 => conv_std_logic_vector(27007, 16),
29168 => conv_std_logic_vector(27120, 16),
29169 => conv_std_logic_vector(27233, 16),
29170 => conv_std_logic_vector(27346, 16),
29171 => conv_std_logic_vector(27459, 16),
29172 => conv_std_logic_vector(27572, 16),
29173 => conv_std_logic_vector(27685, 16),
29174 => conv_std_logic_vector(27798, 16),
29175 => conv_std_logic_vector(27911, 16),
29176 => conv_std_logic_vector(28024, 16),
29177 => conv_std_logic_vector(28137, 16),
29178 => conv_std_logic_vector(28250, 16),
29179 => conv_std_logic_vector(28363, 16),
29180 => conv_std_logic_vector(28476, 16),
29181 => conv_std_logic_vector(28589, 16),
29182 => conv_std_logic_vector(28702, 16),
29183 => conv_std_logic_vector(28815, 16),
29184 => conv_std_logic_vector(0, 16),
29185 => conv_std_logic_vector(114, 16),
29186 => conv_std_logic_vector(228, 16),
29187 => conv_std_logic_vector(342, 16),
29188 => conv_std_logic_vector(456, 16),
29189 => conv_std_logic_vector(570, 16),
29190 => conv_std_logic_vector(684, 16),
29191 => conv_std_logic_vector(798, 16),
29192 => conv_std_logic_vector(912, 16),
29193 => conv_std_logic_vector(1026, 16),
29194 => conv_std_logic_vector(1140, 16),
29195 => conv_std_logic_vector(1254, 16),
29196 => conv_std_logic_vector(1368, 16),
29197 => conv_std_logic_vector(1482, 16),
29198 => conv_std_logic_vector(1596, 16),
29199 => conv_std_logic_vector(1710, 16),
29200 => conv_std_logic_vector(1824, 16),
29201 => conv_std_logic_vector(1938, 16),
29202 => conv_std_logic_vector(2052, 16),
29203 => conv_std_logic_vector(2166, 16),
29204 => conv_std_logic_vector(2280, 16),
29205 => conv_std_logic_vector(2394, 16),
29206 => conv_std_logic_vector(2508, 16),
29207 => conv_std_logic_vector(2622, 16),
29208 => conv_std_logic_vector(2736, 16),
29209 => conv_std_logic_vector(2850, 16),
29210 => conv_std_logic_vector(2964, 16),
29211 => conv_std_logic_vector(3078, 16),
29212 => conv_std_logic_vector(3192, 16),
29213 => conv_std_logic_vector(3306, 16),
29214 => conv_std_logic_vector(3420, 16),
29215 => conv_std_logic_vector(3534, 16),
29216 => conv_std_logic_vector(3648, 16),
29217 => conv_std_logic_vector(3762, 16),
29218 => conv_std_logic_vector(3876, 16),
29219 => conv_std_logic_vector(3990, 16),
29220 => conv_std_logic_vector(4104, 16),
29221 => conv_std_logic_vector(4218, 16),
29222 => conv_std_logic_vector(4332, 16),
29223 => conv_std_logic_vector(4446, 16),
29224 => conv_std_logic_vector(4560, 16),
29225 => conv_std_logic_vector(4674, 16),
29226 => conv_std_logic_vector(4788, 16),
29227 => conv_std_logic_vector(4902, 16),
29228 => conv_std_logic_vector(5016, 16),
29229 => conv_std_logic_vector(5130, 16),
29230 => conv_std_logic_vector(5244, 16),
29231 => conv_std_logic_vector(5358, 16),
29232 => conv_std_logic_vector(5472, 16),
29233 => conv_std_logic_vector(5586, 16),
29234 => conv_std_logic_vector(5700, 16),
29235 => conv_std_logic_vector(5814, 16),
29236 => conv_std_logic_vector(5928, 16),
29237 => conv_std_logic_vector(6042, 16),
29238 => conv_std_logic_vector(6156, 16),
29239 => conv_std_logic_vector(6270, 16),
29240 => conv_std_logic_vector(6384, 16),
29241 => conv_std_logic_vector(6498, 16),
29242 => conv_std_logic_vector(6612, 16),
29243 => conv_std_logic_vector(6726, 16),
29244 => conv_std_logic_vector(6840, 16),
29245 => conv_std_logic_vector(6954, 16),
29246 => conv_std_logic_vector(7068, 16),
29247 => conv_std_logic_vector(7182, 16),
29248 => conv_std_logic_vector(7296, 16),
29249 => conv_std_logic_vector(7410, 16),
29250 => conv_std_logic_vector(7524, 16),
29251 => conv_std_logic_vector(7638, 16),
29252 => conv_std_logic_vector(7752, 16),
29253 => conv_std_logic_vector(7866, 16),
29254 => conv_std_logic_vector(7980, 16),
29255 => conv_std_logic_vector(8094, 16),
29256 => conv_std_logic_vector(8208, 16),
29257 => conv_std_logic_vector(8322, 16),
29258 => conv_std_logic_vector(8436, 16),
29259 => conv_std_logic_vector(8550, 16),
29260 => conv_std_logic_vector(8664, 16),
29261 => conv_std_logic_vector(8778, 16),
29262 => conv_std_logic_vector(8892, 16),
29263 => conv_std_logic_vector(9006, 16),
29264 => conv_std_logic_vector(9120, 16),
29265 => conv_std_logic_vector(9234, 16),
29266 => conv_std_logic_vector(9348, 16),
29267 => conv_std_logic_vector(9462, 16),
29268 => conv_std_logic_vector(9576, 16),
29269 => conv_std_logic_vector(9690, 16),
29270 => conv_std_logic_vector(9804, 16),
29271 => conv_std_logic_vector(9918, 16),
29272 => conv_std_logic_vector(10032, 16),
29273 => conv_std_logic_vector(10146, 16),
29274 => conv_std_logic_vector(10260, 16),
29275 => conv_std_logic_vector(10374, 16),
29276 => conv_std_logic_vector(10488, 16),
29277 => conv_std_logic_vector(10602, 16),
29278 => conv_std_logic_vector(10716, 16),
29279 => conv_std_logic_vector(10830, 16),
29280 => conv_std_logic_vector(10944, 16),
29281 => conv_std_logic_vector(11058, 16),
29282 => conv_std_logic_vector(11172, 16),
29283 => conv_std_logic_vector(11286, 16),
29284 => conv_std_logic_vector(11400, 16),
29285 => conv_std_logic_vector(11514, 16),
29286 => conv_std_logic_vector(11628, 16),
29287 => conv_std_logic_vector(11742, 16),
29288 => conv_std_logic_vector(11856, 16),
29289 => conv_std_logic_vector(11970, 16),
29290 => conv_std_logic_vector(12084, 16),
29291 => conv_std_logic_vector(12198, 16),
29292 => conv_std_logic_vector(12312, 16),
29293 => conv_std_logic_vector(12426, 16),
29294 => conv_std_logic_vector(12540, 16),
29295 => conv_std_logic_vector(12654, 16),
29296 => conv_std_logic_vector(12768, 16),
29297 => conv_std_logic_vector(12882, 16),
29298 => conv_std_logic_vector(12996, 16),
29299 => conv_std_logic_vector(13110, 16),
29300 => conv_std_logic_vector(13224, 16),
29301 => conv_std_logic_vector(13338, 16),
29302 => conv_std_logic_vector(13452, 16),
29303 => conv_std_logic_vector(13566, 16),
29304 => conv_std_logic_vector(13680, 16),
29305 => conv_std_logic_vector(13794, 16),
29306 => conv_std_logic_vector(13908, 16),
29307 => conv_std_logic_vector(14022, 16),
29308 => conv_std_logic_vector(14136, 16),
29309 => conv_std_logic_vector(14250, 16),
29310 => conv_std_logic_vector(14364, 16),
29311 => conv_std_logic_vector(14478, 16),
29312 => conv_std_logic_vector(14592, 16),
29313 => conv_std_logic_vector(14706, 16),
29314 => conv_std_logic_vector(14820, 16),
29315 => conv_std_logic_vector(14934, 16),
29316 => conv_std_logic_vector(15048, 16),
29317 => conv_std_logic_vector(15162, 16),
29318 => conv_std_logic_vector(15276, 16),
29319 => conv_std_logic_vector(15390, 16),
29320 => conv_std_logic_vector(15504, 16),
29321 => conv_std_logic_vector(15618, 16),
29322 => conv_std_logic_vector(15732, 16),
29323 => conv_std_logic_vector(15846, 16),
29324 => conv_std_logic_vector(15960, 16),
29325 => conv_std_logic_vector(16074, 16),
29326 => conv_std_logic_vector(16188, 16),
29327 => conv_std_logic_vector(16302, 16),
29328 => conv_std_logic_vector(16416, 16),
29329 => conv_std_logic_vector(16530, 16),
29330 => conv_std_logic_vector(16644, 16),
29331 => conv_std_logic_vector(16758, 16),
29332 => conv_std_logic_vector(16872, 16),
29333 => conv_std_logic_vector(16986, 16),
29334 => conv_std_logic_vector(17100, 16),
29335 => conv_std_logic_vector(17214, 16),
29336 => conv_std_logic_vector(17328, 16),
29337 => conv_std_logic_vector(17442, 16),
29338 => conv_std_logic_vector(17556, 16),
29339 => conv_std_logic_vector(17670, 16),
29340 => conv_std_logic_vector(17784, 16),
29341 => conv_std_logic_vector(17898, 16),
29342 => conv_std_logic_vector(18012, 16),
29343 => conv_std_logic_vector(18126, 16),
29344 => conv_std_logic_vector(18240, 16),
29345 => conv_std_logic_vector(18354, 16),
29346 => conv_std_logic_vector(18468, 16),
29347 => conv_std_logic_vector(18582, 16),
29348 => conv_std_logic_vector(18696, 16),
29349 => conv_std_logic_vector(18810, 16),
29350 => conv_std_logic_vector(18924, 16),
29351 => conv_std_logic_vector(19038, 16),
29352 => conv_std_logic_vector(19152, 16),
29353 => conv_std_logic_vector(19266, 16),
29354 => conv_std_logic_vector(19380, 16),
29355 => conv_std_logic_vector(19494, 16),
29356 => conv_std_logic_vector(19608, 16),
29357 => conv_std_logic_vector(19722, 16),
29358 => conv_std_logic_vector(19836, 16),
29359 => conv_std_logic_vector(19950, 16),
29360 => conv_std_logic_vector(20064, 16),
29361 => conv_std_logic_vector(20178, 16),
29362 => conv_std_logic_vector(20292, 16),
29363 => conv_std_logic_vector(20406, 16),
29364 => conv_std_logic_vector(20520, 16),
29365 => conv_std_logic_vector(20634, 16),
29366 => conv_std_logic_vector(20748, 16),
29367 => conv_std_logic_vector(20862, 16),
29368 => conv_std_logic_vector(20976, 16),
29369 => conv_std_logic_vector(21090, 16),
29370 => conv_std_logic_vector(21204, 16),
29371 => conv_std_logic_vector(21318, 16),
29372 => conv_std_logic_vector(21432, 16),
29373 => conv_std_logic_vector(21546, 16),
29374 => conv_std_logic_vector(21660, 16),
29375 => conv_std_logic_vector(21774, 16),
29376 => conv_std_logic_vector(21888, 16),
29377 => conv_std_logic_vector(22002, 16),
29378 => conv_std_logic_vector(22116, 16),
29379 => conv_std_logic_vector(22230, 16),
29380 => conv_std_logic_vector(22344, 16),
29381 => conv_std_logic_vector(22458, 16),
29382 => conv_std_logic_vector(22572, 16),
29383 => conv_std_logic_vector(22686, 16),
29384 => conv_std_logic_vector(22800, 16),
29385 => conv_std_logic_vector(22914, 16),
29386 => conv_std_logic_vector(23028, 16),
29387 => conv_std_logic_vector(23142, 16),
29388 => conv_std_logic_vector(23256, 16),
29389 => conv_std_logic_vector(23370, 16),
29390 => conv_std_logic_vector(23484, 16),
29391 => conv_std_logic_vector(23598, 16),
29392 => conv_std_logic_vector(23712, 16),
29393 => conv_std_logic_vector(23826, 16),
29394 => conv_std_logic_vector(23940, 16),
29395 => conv_std_logic_vector(24054, 16),
29396 => conv_std_logic_vector(24168, 16),
29397 => conv_std_logic_vector(24282, 16),
29398 => conv_std_logic_vector(24396, 16),
29399 => conv_std_logic_vector(24510, 16),
29400 => conv_std_logic_vector(24624, 16),
29401 => conv_std_logic_vector(24738, 16),
29402 => conv_std_logic_vector(24852, 16),
29403 => conv_std_logic_vector(24966, 16),
29404 => conv_std_logic_vector(25080, 16),
29405 => conv_std_logic_vector(25194, 16),
29406 => conv_std_logic_vector(25308, 16),
29407 => conv_std_logic_vector(25422, 16),
29408 => conv_std_logic_vector(25536, 16),
29409 => conv_std_logic_vector(25650, 16),
29410 => conv_std_logic_vector(25764, 16),
29411 => conv_std_logic_vector(25878, 16),
29412 => conv_std_logic_vector(25992, 16),
29413 => conv_std_logic_vector(26106, 16),
29414 => conv_std_logic_vector(26220, 16),
29415 => conv_std_logic_vector(26334, 16),
29416 => conv_std_logic_vector(26448, 16),
29417 => conv_std_logic_vector(26562, 16),
29418 => conv_std_logic_vector(26676, 16),
29419 => conv_std_logic_vector(26790, 16),
29420 => conv_std_logic_vector(26904, 16),
29421 => conv_std_logic_vector(27018, 16),
29422 => conv_std_logic_vector(27132, 16),
29423 => conv_std_logic_vector(27246, 16),
29424 => conv_std_logic_vector(27360, 16),
29425 => conv_std_logic_vector(27474, 16),
29426 => conv_std_logic_vector(27588, 16),
29427 => conv_std_logic_vector(27702, 16),
29428 => conv_std_logic_vector(27816, 16),
29429 => conv_std_logic_vector(27930, 16),
29430 => conv_std_logic_vector(28044, 16),
29431 => conv_std_logic_vector(28158, 16),
29432 => conv_std_logic_vector(28272, 16),
29433 => conv_std_logic_vector(28386, 16),
29434 => conv_std_logic_vector(28500, 16),
29435 => conv_std_logic_vector(28614, 16),
29436 => conv_std_logic_vector(28728, 16),
29437 => conv_std_logic_vector(28842, 16),
29438 => conv_std_logic_vector(28956, 16),
29439 => conv_std_logic_vector(29070, 16),
29440 => conv_std_logic_vector(0, 16),
29441 => conv_std_logic_vector(115, 16),
29442 => conv_std_logic_vector(230, 16),
29443 => conv_std_logic_vector(345, 16),
29444 => conv_std_logic_vector(460, 16),
29445 => conv_std_logic_vector(575, 16),
29446 => conv_std_logic_vector(690, 16),
29447 => conv_std_logic_vector(805, 16),
29448 => conv_std_logic_vector(920, 16),
29449 => conv_std_logic_vector(1035, 16),
29450 => conv_std_logic_vector(1150, 16),
29451 => conv_std_logic_vector(1265, 16),
29452 => conv_std_logic_vector(1380, 16),
29453 => conv_std_logic_vector(1495, 16),
29454 => conv_std_logic_vector(1610, 16),
29455 => conv_std_logic_vector(1725, 16),
29456 => conv_std_logic_vector(1840, 16),
29457 => conv_std_logic_vector(1955, 16),
29458 => conv_std_logic_vector(2070, 16),
29459 => conv_std_logic_vector(2185, 16),
29460 => conv_std_logic_vector(2300, 16),
29461 => conv_std_logic_vector(2415, 16),
29462 => conv_std_logic_vector(2530, 16),
29463 => conv_std_logic_vector(2645, 16),
29464 => conv_std_logic_vector(2760, 16),
29465 => conv_std_logic_vector(2875, 16),
29466 => conv_std_logic_vector(2990, 16),
29467 => conv_std_logic_vector(3105, 16),
29468 => conv_std_logic_vector(3220, 16),
29469 => conv_std_logic_vector(3335, 16),
29470 => conv_std_logic_vector(3450, 16),
29471 => conv_std_logic_vector(3565, 16),
29472 => conv_std_logic_vector(3680, 16),
29473 => conv_std_logic_vector(3795, 16),
29474 => conv_std_logic_vector(3910, 16),
29475 => conv_std_logic_vector(4025, 16),
29476 => conv_std_logic_vector(4140, 16),
29477 => conv_std_logic_vector(4255, 16),
29478 => conv_std_logic_vector(4370, 16),
29479 => conv_std_logic_vector(4485, 16),
29480 => conv_std_logic_vector(4600, 16),
29481 => conv_std_logic_vector(4715, 16),
29482 => conv_std_logic_vector(4830, 16),
29483 => conv_std_logic_vector(4945, 16),
29484 => conv_std_logic_vector(5060, 16),
29485 => conv_std_logic_vector(5175, 16),
29486 => conv_std_logic_vector(5290, 16),
29487 => conv_std_logic_vector(5405, 16),
29488 => conv_std_logic_vector(5520, 16),
29489 => conv_std_logic_vector(5635, 16),
29490 => conv_std_logic_vector(5750, 16),
29491 => conv_std_logic_vector(5865, 16),
29492 => conv_std_logic_vector(5980, 16),
29493 => conv_std_logic_vector(6095, 16),
29494 => conv_std_logic_vector(6210, 16),
29495 => conv_std_logic_vector(6325, 16),
29496 => conv_std_logic_vector(6440, 16),
29497 => conv_std_logic_vector(6555, 16),
29498 => conv_std_logic_vector(6670, 16),
29499 => conv_std_logic_vector(6785, 16),
29500 => conv_std_logic_vector(6900, 16),
29501 => conv_std_logic_vector(7015, 16),
29502 => conv_std_logic_vector(7130, 16),
29503 => conv_std_logic_vector(7245, 16),
29504 => conv_std_logic_vector(7360, 16),
29505 => conv_std_logic_vector(7475, 16),
29506 => conv_std_logic_vector(7590, 16),
29507 => conv_std_logic_vector(7705, 16),
29508 => conv_std_logic_vector(7820, 16),
29509 => conv_std_logic_vector(7935, 16),
29510 => conv_std_logic_vector(8050, 16),
29511 => conv_std_logic_vector(8165, 16),
29512 => conv_std_logic_vector(8280, 16),
29513 => conv_std_logic_vector(8395, 16),
29514 => conv_std_logic_vector(8510, 16),
29515 => conv_std_logic_vector(8625, 16),
29516 => conv_std_logic_vector(8740, 16),
29517 => conv_std_logic_vector(8855, 16),
29518 => conv_std_logic_vector(8970, 16),
29519 => conv_std_logic_vector(9085, 16),
29520 => conv_std_logic_vector(9200, 16),
29521 => conv_std_logic_vector(9315, 16),
29522 => conv_std_logic_vector(9430, 16),
29523 => conv_std_logic_vector(9545, 16),
29524 => conv_std_logic_vector(9660, 16),
29525 => conv_std_logic_vector(9775, 16),
29526 => conv_std_logic_vector(9890, 16),
29527 => conv_std_logic_vector(10005, 16),
29528 => conv_std_logic_vector(10120, 16),
29529 => conv_std_logic_vector(10235, 16),
29530 => conv_std_logic_vector(10350, 16),
29531 => conv_std_logic_vector(10465, 16),
29532 => conv_std_logic_vector(10580, 16),
29533 => conv_std_logic_vector(10695, 16),
29534 => conv_std_logic_vector(10810, 16),
29535 => conv_std_logic_vector(10925, 16),
29536 => conv_std_logic_vector(11040, 16),
29537 => conv_std_logic_vector(11155, 16),
29538 => conv_std_logic_vector(11270, 16),
29539 => conv_std_logic_vector(11385, 16),
29540 => conv_std_logic_vector(11500, 16),
29541 => conv_std_logic_vector(11615, 16),
29542 => conv_std_logic_vector(11730, 16),
29543 => conv_std_logic_vector(11845, 16),
29544 => conv_std_logic_vector(11960, 16),
29545 => conv_std_logic_vector(12075, 16),
29546 => conv_std_logic_vector(12190, 16),
29547 => conv_std_logic_vector(12305, 16),
29548 => conv_std_logic_vector(12420, 16),
29549 => conv_std_logic_vector(12535, 16),
29550 => conv_std_logic_vector(12650, 16),
29551 => conv_std_logic_vector(12765, 16),
29552 => conv_std_logic_vector(12880, 16),
29553 => conv_std_logic_vector(12995, 16),
29554 => conv_std_logic_vector(13110, 16),
29555 => conv_std_logic_vector(13225, 16),
29556 => conv_std_logic_vector(13340, 16),
29557 => conv_std_logic_vector(13455, 16),
29558 => conv_std_logic_vector(13570, 16),
29559 => conv_std_logic_vector(13685, 16),
29560 => conv_std_logic_vector(13800, 16),
29561 => conv_std_logic_vector(13915, 16),
29562 => conv_std_logic_vector(14030, 16),
29563 => conv_std_logic_vector(14145, 16),
29564 => conv_std_logic_vector(14260, 16),
29565 => conv_std_logic_vector(14375, 16),
29566 => conv_std_logic_vector(14490, 16),
29567 => conv_std_logic_vector(14605, 16),
29568 => conv_std_logic_vector(14720, 16),
29569 => conv_std_logic_vector(14835, 16),
29570 => conv_std_logic_vector(14950, 16),
29571 => conv_std_logic_vector(15065, 16),
29572 => conv_std_logic_vector(15180, 16),
29573 => conv_std_logic_vector(15295, 16),
29574 => conv_std_logic_vector(15410, 16),
29575 => conv_std_logic_vector(15525, 16),
29576 => conv_std_logic_vector(15640, 16),
29577 => conv_std_logic_vector(15755, 16),
29578 => conv_std_logic_vector(15870, 16),
29579 => conv_std_logic_vector(15985, 16),
29580 => conv_std_logic_vector(16100, 16),
29581 => conv_std_logic_vector(16215, 16),
29582 => conv_std_logic_vector(16330, 16),
29583 => conv_std_logic_vector(16445, 16),
29584 => conv_std_logic_vector(16560, 16),
29585 => conv_std_logic_vector(16675, 16),
29586 => conv_std_logic_vector(16790, 16),
29587 => conv_std_logic_vector(16905, 16),
29588 => conv_std_logic_vector(17020, 16),
29589 => conv_std_logic_vector(17135, 16),
29590 => conv_std_logic_vector(17250, 16),
29591 => conv_std_logic_vector(17365, 16),
29592 => conv_std_logic_vector(17480, 16),
29593 => conv_std_logic_vector(17595, 16),
29594 => conv_std_logic_vector(17710, 16),
29595 => conv_std_logic_vector(17825, 16),
29596 => conv_std_logic_vector(17940, 16),
29597 => conv_std_logic_vector(18055, 16),
29598 => conv_std_logic_vector(18170, 16),
29599 => conv_std_logic_vector(18285, 16),
29600 => conv_std_logic_vector(18400, 16),
29601 => conv_std_logic_vector(18515, 16),
29602 => conv_std_logic_vector(18630, 16),
29603 => conv_std_logic_vector(18745, 16),
29604 => conv_std_logic_vector(18860, 16),
29605 => conv_std_logic_vector(18975, 16),
29606 => conv_std_logic_vector(19090, 16),
29607 => conv_std_logic_vector(19205, 16),
29608 => conv_std_logic_vector(19320, 16),
29609 => conv_std_logic_vector(19435, 16),
29610 => conv_std_logic_vector(19550, 16),
29611 => conv_std_logic_vector(19665, 16),
29612 => conv_std_logic_vector(19780, 16),
29613 => conv_std_logic_vector(19895, 16),
29614 => conv_std_logic_vector(20010, 16),
29615 => conv_std_logic_vector(20125, 16),
29616 => conv_std_logic_vector(20240, 16),
29617 => conv_std_logic_vector(20355, 16),
29618 => conv_std_logic_vector(20470, 16),
29619 => conv_std_logic_vector(20585, 16),
29620 => conv_std_logic_vector(20700, 16),
29621 => conv_std_logic_vector(20815, 16),
29622 => conv_std_logic_vector(20930, 16),
29623 => conv_std_logic_vector(21045, 16),
29624 => conv_std_logic_vector(21160, 16),
29625 => conv_std_logic_vector(21275, 16),
29626 => conv_std_logic_vector(21390, 16),
29627 => conv_std_logic_vector(21505, 16),
29628 => conv_std_logic_vector(21620, 16),
29629 => conv_std_logic_vector(21735, 16),
29630 => conv_std_logic_vector(21850, 16),
29631 => conv_std_logic_vector(21965, 16),
29632 => conv_std_logic_vector(22080, 16),
29633 => conv_std_logic_vector(22195, 16),
29634 => conv_std_logic_vector(22310, 16),
29635 => conv_std_logic_vector(22425, 16),
29636 => conv_std_logic_vector(22540, 16),
29637 => conv_std_logic_vector(22655, 16),
29638 => conv_std_logic_vector(22770, 16),
29639 => conv_std_logic_vector(22885, 16),
29640 => conv_std_logic_vector(23000, 16),
29641 => conv_std_logic_vector(23115, 16),
29642 => conv_std_logic_vector(23230, 16),
29643 => conv_std_logic_vector(23345, 16),
29644 => conv_std_logic_vector(23460, 16),
29645 => conv_std_logic_vector(23575, 16),
29646 => conv_std_logic_vector(23690, 16),
29647 => conv_std_logic_vector(23805, 16),
29648 => conv_std_logic_vector(23920, 16),
29649 => conv_std_logic_vector(24035, 16),
29650 => conv_std_logic_vector(24150, 16),
29651 => conv_std_logic_vector(24265, 16),
29652 => conv_std_logic_vector(24380, 16),
29653 => conv_std_logic_vector(24495, 16),
29654 => conv_std_logic_vector(24610, 16),
29655 => conv_std_logic_vector(24725, 16),
29656 => conv_std_logic_vector(24840, 16),
29657 => conv_std_logic_vector(24955, 16),
29658 => conv_std_logic_vector(25070, 16),
29659 => conv_std_logic_vector(25185, 16),
29660 => conv_std_logic_vector(25300, 16),
29661 => conv_std_logic_vector(25415, 16),
29662 => conv_std_logic_vector(25530, 16),
29663 => conv_std_logic_vector(25645, 16),
29664 => conv_std_logic_vector(25760, 16),
29665 => conv_std_logic_vector(25875, 16),
29666 => conv_std_logic_vector(25990, 16),
29667 => conv_std_logic_vector(26105, 16),
29668 => conv_std_logic_vector(26220, 16),
29669 => conv_std_logic_vector(26335, 16),
29670 => conv_std_logic_vector(26450, 16),
29671 => conv_std_logic_vector(26565, 16),
29672 => conv_std_logic_vector(26680, 16),
29673 => conv_std_logic_vector(26795, 16),
29674 => conv_std_logic_vector(26910, 16),
29675 => conv_std_logic_vector(27025, 16),
29676 => conv_std_logic_vector(27140, 16),
29677 => conv_std_logic_vector(27255, 16),
29678 => conv_std_logic_vector(27370, 16),
29679 => conv_std_logic_vector(27485, 16),
29680 => conv_std_logic_vector(27600, 16),
29681 => conv_std_logic_vector(27715, 16),
29682 => conv_std_logic_vector(27830, 16),
29683 => conv_std_logic_vector(27945, 16),
29684 => conv_std_logic_vector(28060, 16),
29685 => conv_std_logic_vector(28175, 16),
29686 => conv_std_logic_vector(28290, 16),
29687 => conv_std_logic_vector(28405, 16),
29688 => conv_std_logic_vector(28520, 16),
29689 => conv_std_logic_vector(28635, 16),
29690 => conv_std_logic_vector(28750, 16),
29691 => conv_std_logic_vector(28865, 16),
29692 => conv_std_logic_vector(28980, 16),
29693 => conv_std_logic_vector(29095, 16),
29694 => conv_std_logic_vector(29210, 16),
29695 => conv_std_logic_vector(29325, 16),
29696 => conv_std_logic_vector(0, 16),
29697 => conv_std_logic_vector(116, 16),
29698 => conv_std_logic_vector(232, 16),
29699 => conv_std_logic_vector(348, 16),
29700 => conv_std_logic_vector(464, 16),
29701 => conv_std_logic_vector(580, 16),
29702 => conv_std_logic_vector(696, 16),
29703 => conv_std_logic_vector(812, 16),
29704 => conv_std_logic_vector(928, 16),
29705 => conv_std_logic_vector(1044, 16),
29706 => conv_std_logic_vector(1160, 16),
29707 => conv_std_logic_vector(1276, 16),
29708 => conv_std_logic_vector(1392, 16),
29709 => conv_std_logic_vector(1508, 16),
29710 => conv_std_logic_vector(1624, 16),
29711 => conv_std_logic_vector(1740, 16),
29712 => conv_std_logic_vector(1856, 16),
29713 => conv_std_logic_vector(1972, 16),
29714 => conv_std_logic_vector(2088, 16),
29715 => conv_std_logic_vector(2204, 16),
29716 => conv_std_logic_vector(2320, 16),
29717 => conv_std_logic_vector(2436, 16),
29718 => conv_std_logic_vector(2552, 16),
29719 => conv_std_logic_vector(2668, 16),
29720 => conv_std_logic_vector(2784, 16),
29721 => conv_std_logic_vector(2900, 16),
29722 => conv_std_logic_vector(3016, 16),
29723 => conv_std_logic_vector(3132, 16),
29724 => conv_std_logic_vector(3248, 16),
29725 => conv_std_logic_vector(3364, 16),
29726 => conv_std_logic_vector(3480, 16),
29727 => conv_std_logic_vector(3596, 16),
29728 => conv_std_logic_vector(3712, 16),
29729 => conv_std_logic_vector(3828, 16),
29730 => conv_std_logic_vector(3944, 16),
29731 => conv_std_logic_vector(4060, 16),
29732 => conv_std_logic_vector(4176, 16),
29733 => conv_std_logic_vector(4292, 16),
29734 => conv_std_logic_vector(4408, 16),
29735 => conv_std_logic_vector(4524, 16),
29736 => conv_std_logic_vector(4640, 16),
29737 => conv_std_logic_vector(4756, 16),
29738 => conv_std_logic_vector(4872, 16),
29739 => conv_std_logic_vector(4988, 16),
29740 => conv_std_logic_vector(5104, 16),
29741 => conv_std_logic_vector(5220, 16),
29742 => conv_std_logic_vector(5336, 16),
29743 => conv_std_logic_vector(5452, 16),
29744 => conv_std_logic_vector(5568, 16),
29745 => conv_std_logic_vector(5684, 16),
29746 => conv_std_logic_vector(5800, 16),
29747 => conv_std_logic_vector(5916, 16),
29748 => conv_std_logic_vector(6032, 16),
29749 => conv_std_logic_vector(6148, 16),
29750 => conv_std_logic_vector(6264, 16),
29751 => conv_std_logic_vector(6380, 16),
29752 => conv_std_logic_vector(6496, 16),
29753 => conv_std_logic_vector(6612, 16),
29754 => conv_std_logic_vector(6728, 16),
29755 => conv_std_logic_vector(6844, 16),
29756 => conv_std_logic_vector(6960, 16),
29757 => conv_std_logic_vector(7076, 16),
29758 => conv_std_logic_vector(7192, 16),
29759 => conv_std_logic_vector(7308, 16),
29760 => conv_std_logic_vector(7424, 16),
29761 => conv_std_logic_vector(7540, 16),
29762 => conv_std_logic_vector(7656, 16),
29763 => conv_std_logic_vector(7772, 16),
29764 => conv_std_logic_vector(7888, 16),
29765 => conv_std_logic_vector(8004, 16),
29766 => conv_std_logic_vector(8120, 16),
29767 => conv_std_logic_vector(8236, 16),
29768 => conv_std_logic_vector(8352, 16),
29769 => conv_std_logic_vector(8468, 16),
29770 => conv_std_logic_vector(8584, 16),
29771 => conv_std_logic_vector(8700, 16),
29772 => conv_std_logic_vector(8816, 16),
29773 => conv_std_logic_vector(8932, 16),
29774 => conv_std_logic_vector(9048, 16),
29775 => conv_std_logic_vector(9164, 16),
29776 => conv_std_logic_vector(9280, 16),
29777 => conv_std_logic_vector(9396, 16),
29778 => conv_std_logic_vector(9512, 16),
29779 => conv_std_logic_vector(9628, 16),
29780 => conv_std_logic_vector(9744, 16),
29781 => conv_std_logic_vector(9860, 16),
29782 => conv_std_logic_vector(9976, 16),
29783 => conv_std_logic_vector(10092, 16),
29784 => conv_std_logic_vector(10208, 16),
29785 => conv_std_logic_vector(10324, 16),
29786 => conv_std_logic_vector(10440, 16),
29787 => conv_std_logic_vector(10556, 16),
29788 => conv_std_logic_vector(10672, 16),
29789 => conv_std_logic_vector(10788, 16),
29790 => conv_std_logic_vector(10904, 16),
29791 => conv_std_logic_vector(11020, 16),
29792 => conv_std_logic_vector(11136, 16),
29793 => conv_std_logic_vector(11252, 16),
29794 => conv_std_logic_vector(11368, 16),
29795 => conv_std_logic_vector(11484, 16),
29796 => conv_std_logic_vector(11600, 16),
29797 => conv_std_logic_vector(11716, 16),
29798 => conv_std_logic_vector(11832, 16),
29799 => conv_std_logic_vector(11948, 16),
29800 => conv_std_logic_vector(12064, 16),
29801 => conv_std_logic_vector(12180, 16),
29802 => conv_std_logic_vector(12296, 16),
29803 => conv_std_logic_vector(12412, 16),
29804 => conv_std_logic_vector(12528, 16),
29805 => conv_std_logic_vector(12644, 16),
29806 => conv_std_logic_vector(12760, 16),
29807 => conv_std_logic_vector(12876, 16),
29808 => conv_std_logic_vector(12992, 16),
29809 => conv_std_logic_vector(13108, 16),
29810 => conv_std_logic_vector(13224, 16),
29811 => conv_std_logic_vector(13340, 16),
29812 => conv_std_logic_vector(13456, 16),
29813 => conv_std_logic_vector(13572, 16),
29814 => conv_std_logic_vector(13688, 16),
29815 => conv_std_logic_vector(13804, 16),
29816 => conv_std_logic_vector(13920, 16),
29817 => conv_std_logic_vector(14036, 16),
29818 => conv_std_logic_vector(14152, 16),
29819 => conv_std_logic_vector(14268, 16),
29820 => conv_std_logic_vector(14384, 16),
29821 => conv_std_logic_vector(14500, 16),
29822 => conv_std_logic_vector(14616, 16),
29823 => conv_std_logic_vector(14732, 16),
29824 => conv_std_logic_vector(14848, 16),
29825 => conv_std_logic_vector(14964, 16),
29826 => conv_std_logic_vector(15080, 16),
29827 => conv_std_logic_vector(15196, 16),
29828 => conv_std_logic_vector(15312, 16),
29829 => conv_std_logic_vector(15428, 16),
29830 => conv_std_logic_vector(15544, 16),
29831 => conv_std_logic_vector(15660, 16),
29832 => conv_std_logic_vector(15776, 16),
29833 => conv_std_logic_vector(15892, 16),
29834 => conv_std_logic_vector(16008, 16),
29835 => conv_std_logic_vector(16124, 16),
29836 => conv_std_logic_vector(16240, 16),
29837 => conv_std_logic_vector(16356, 16),
29838 => conv_std_logic_vector(16472, 16),
29839 => conv_std_logic_vector(16588, 16),
29840 => conv_std_logic_vector(16704, 16),
29841 => conv_std_logic_vector(16820, 16),
29842 => conv_std_logic_vector(16936, 16),
29843 => conv_std_logic_vector(17052, 16),
29844 => conv_std_logic_vector(17168, 16),
29845 => conv_std_logic_vector(17284, 16),
29846 => conv_std_logic_vector(17400, 16),
29847 => conv_std_logic_vector(17516, 16),
29848 => conv_std_logic_vector(17632, 16),
29849 => conv_std_logic_vector(17748, 16),
29850 => conv_std_logic_vector(17864, 16),
29851 => conv_std_logic_vector(17980, 16),
29852 => conv_std_logic_vector(18096, 16),
29853 => conv_std_logic_vector(18212, 16),
29854 => conv_std_logic_vector(18328, 16),
29855 => conv_std_logic_vector(18444, 16),
29856 => conv_std_logic_vector(18560, 16),
29857 => conv_std_logic_vector(18676, 16),
29858 => conv_std_logic_vector(18792, 16),
29859 => conv_std_logic_vector(18908, 16),
29860 => conv_std_logic_vector(19024, 16),
29861 => conv_std_logic_vector(19140, 16),
29862 => conv_std_logic_vector(19256, 16),
29863 => conv_std_logic_vector(19372, 16),
29864 => conv_std_logic_vector(19488, 16),
29865 => conv_std_logic_vector(19604, 16),
29866 => conv_std_logic_vector(19720, 16),
29867 => conv_std_logic_vector(19836, 16),
29868 => conv_std_logic_vector(19952, 16),
29869 => conv_std_logic_vector(20068, 16),
29870 => conv_std_logic_vector(20184, 16),
29871 => conv_std_logic_vector(20300, 16),
29872 => conv_std_logic_vector(20416, 16),
29873 => conv_std_logic_vector(20532, 16),
29874 => conv_std_logic_vector(20648, 16),
29875 => conv_std_logic_vector(20764, 16),
29876 => conv_std_logic_vector(20880, 16),
29877 => conv_std_logic_vector(20996, 16),
29878 => conv_std_logic_vector(21112, 16),
29879 => conv_std_logic_vector(21228, 16),
29880 => conv_std_logic_vector(21344, 16),
29881 => conv_std_logic_vector(21460, 16),
29882 => conv_std_logic_vector(21576, 16),
29883 => conv_std_logic_vector(21692, 16),
29884 => conv_std_logic_vector(21808, 16),
29885 => conv_std_logic_vector(21924, 16),
29886 => conv_std_logic_vector(22040, 16),
29887 => conv_std_logic_vector(22156, 16),
29888 => conv_std_logic_vector(22272, 16),
29889 => conv_std_logic_vector(22388, 16),
29890 => conv_std_logic_vector(22504, 16),
29891 => conv_std_logic_vector(22620, 16),
29892 => conv_std_logic_vector(22736, 16),
29893 => conv_std_logic_vector(22852, 16),
29894 => conv_std_logic_vector(22968, 16),
29895 => conv_std_logic_vector(23084, 16),
29896 => conv_std_logic_vector(23200, 16),
29897 => conv_std_logic_vector(23316, 16),
29898 => conv_std_logic_vector(23432, 16),
29899 => conv_std_logic_vector(23548, 16),
29900 => conv_std_logic_vector(23664, 16),
29901 => conv_std_logic_vector(23780, 16),
29902 => conv_std_logic_vector(23896, 16),
29903 => conv_std_logic_vector(24012, 16),
29904 => conv_std_logic_vector(24128, 16),
29905 => conv_std_logic_vector(24244, 16),
29906 => conv_std_logic_vector(24360, 16),
29907 => conv_std_logic_vector(24476, 16),
29908 => conv_std_logic_vector(24592, 16),
29909 => conv_std_logic_vector(24708, 16),
29910 => conv_std_logic_vector(24824, 16),
29911 => conv_std_logic_vector(24940, 16),
29912 => conv_std_logic_vector(25056, 16),
29913 => conv_std_logic_vector(25172, 16),
29914 => conv_std_logic_vector(25288, 16),
29915 => conv_std_logic_vector(25404, 16),
29916 => conv_std_logic_vector(25520, 16),
29917 => conv_std_logic_vector(25636, 16),
29918 => conv_std_logic_vector(25752, 16),
29919 => conv_std_logic_vector(25868, 16),
29920 => conv_std_logic_vector(25984, 16),
29921 => conv_std_logic_vector(26100, 16),
29922 => conv_std_logic_vector(26216, 16),
29923 => conv_std_logic_vector(26332, 16),
29924 => conv_std_logic_vector(26448, 16),
29925 => conv_std_logic_vector(26564, 16),
29926 => conv_std_logic_vector(26680, 16),
29927 => conv_std_logic_vector(26796, 16),
29928 => conv_std_logic_vector(26912, 16),
29929 => conv_std_logic_vector(27028, 16),
29930 => conv_std_logic_vector(27144, 16),
29931 => conv_std_logic_vector(27260, 16),
29932 => conv_std_logic_vector(27376, 16),
29933 => conv_std_logic_vector(27492, 16),
29934 => conv_std_logic_vector(27608, 16),
29935 => conv_std_logic_vector(27724, 16),
29936 => conv_std_logic_vector(27840, 16),
29937 => conv_std_logic_vector(27956, 16),
29938 => conv_std_logic_vector(28072, 16),
29939 => conv_std_logic_vector(28188, 16),
29940 => conv_std_logic_vector(28304, 16),
29941 => conv_std_logic_vector(28420, 16),
29942 => conv_std_logic_vector(28536, 16),
29943 => conv_std_logic_vector(28652, 16),
29944 => conv_std_logic_vector(28768, 16),
29945 => conv_std_logic_vector(28884, 16),
29946 => conv_std_logic_vector(29000, 16),
29947 => conv_std_logic_vector(29116, 16),
29948 => conv_std_logic_vector(29232, 16),
29949 => conv_std_logic_vector(29348, 16),
29950 => conv_std_logic_vector(29464, 16),
29951 => conv_std_logic_vector(29580, 16),
29952 => conv_std_logic_vector(0, 16),
29953 => conv_std_logic_vector(117, 16),
29954 => conv_std_logic_vector(234, 16),
29955 => conv_std_logic_vector(351, 16),
29956 => conv_std_logic_vector(468, 16),
29957 => conv_std_logic_vector(585, 16),
29958 => conv_std_logic_vector(702, 16),
29959 => conv_std_logic_vector(819, 16),
29960 => conv_std_logic_vector(936, 16),
29961 => conv_std_logic_vector(1053, 16),
29962 => conv_std_logic_vector(1170, 16),
29963 => conv_std_logic_vector(1287, 16),
29964 => conv_std_logic_vector(1404, 16),
29965 => conv_std_logic_vector(1521, 16),
29966 => conv_std_logic_vector(1638, 16),
29967 => conv_std_logic_vector(1755, 16),
29968 => conv_std_logic_vector(1872, 16),
29969 => conv_std_logic_vector(1989, 16),
29970 => conv_std_logic_vector(2106, 16),
29971 => conv_std_logic_vector(2223, 16),
29972 => conv_std_logic_vector(2340, 16),
29973 => conv_std_logic_vector(2457, 16),
29974 => conv_std_logic_vector(2574, 16),
29975 => conv_std_logic_vector(2691, 16),
29976 => conv_std_logic_vector(2808, 16),
29977 => conv_std_logic_vector(2925, 16),
29978 => conv_std_logic_vector(3042, 16),
29979 => conv_std_logic_vector(3159, 16),
29980 => conv_std_logic_vector(3276, 16),
29981 => conv_std_logic_vector(3393, 16),
29982 => conv_std_logic_vector(3510, 16),
29983 => conv_std_logic_vector(3627, 16),
29984 => conv_std_logic_vector(3744, 16),
29985 => conv_std_logic_vector(3861, 16),
29986 => conv_std_logic_vector(3978, 16),
29987 => conv_std_logic_vector(4095, 16),
29988 => conv_std_logic_vector(4212, 16),
29989 => conv_std_logic_vector(4329, 16),
29990 => conv_std_logic_vector(4446, 16),
29991 => conv_std_logic_vector(4563, 16),
29992 => conv_std_logic_vector(4680, 16),
29993 => conv_std_logic_vector(4797, 16),
29994 => conv_std_logic_vector(4914, 16),
29995 => conv_std_logic_vector(5031, 16),
29996 => conv_std_logic_vector(5148, 16),
29997 => conv_std_logic_vector(5265, 16),
29998 => conv_std_logic_vector(5382, 16),
29999 => conv_std_logic_vector(5499, 16),
30000 => conv_std_logic_vector(5616, 16),
30001 => conv_std_logic_vector(5733, 16),
30002 => conv_std_logic_vector(5850, 16),
30003 => conv_std_logic_vector(5967, 16),
30004 => conv_std_logic_vector(6084, 16),
30005 => conv_std_logic_vector(6201, 16),
30006 => conv_std_logic_vector(6318, 16),
30007 => conv_std_logic_vector(6435, 16),
30008 => conv_std_logic_vector(6552, 16),
30009 => conv_std_logic_vector(6669, 16),
30010 => conv_std_logic_vector(6786, 16),
30011 => conv_std_logic_vector(6903, 16),
30012 => conv_std_logic_vector(7020, 16),
30013 => conv_std_logic_vector(7137, 16),
30014 => conv_std_logic_vector(7254, 16),
30015 => conv_std_logic_vector(7371, 16),
30016 => conv_std_logic_vector(7488, 16),
30017 => conv_std_logic_vector(7605, 16),
30018 => conv_std_logic_vector(7722, 16),
30019 => conv_std_logic_vector(7839, 16),
30020 => conv_std_logic_vector(7956, 16),
30021 => conv_std_logic_vector(8073, 16),
30022 => conv_std_logic_vector(8190, 16),
30023 => conv_std_logic_vector(8307, 16),
30024 => conv_std_logic_vector(8424, 16),
30025 => conv_std_logic_vector(8541, 16),
30026 => conv_std_logic_vector(8658, 16),
30027 => conv_std_logic_vector(8775, 16),
30028 => conv_std_logic_vector(8892, 16),
30029 => conv_std_logic_vector(9009, 16),
30030 => conv_std_logic_vector(9126, 16),
30031 => conv_std_logic_vector(9243, 16),
30032 => conv_std_logic_vector(9360, 16),
30033 => conv_std_logic_vector(9477, 16),
30034 => conv_std_logic_vector(9594, 16),
30035 => conv_std_logic_vector(9711, 16),
30036 => conv_std_logic_vector(9828, 16),
30037 => conv_std_logic_vector(9945, 16),
30038 => conv_std_logic_vector(10062, 16),
30039 => conv_std_logic_vector(10179, 16),
30040 => conv_std_logic_vector(10296, 16),
30041 => conv_std_logic_vector(10413, 16),
30042 => conv_std_logic_vector(10530, 16),
30043 => conv_std_logic_vector(10647, 16),
30044 => conv_std_logic_vector(10764, 16),
30045 => conv_std_logic_vector(10881, 16),
30046 => conv_std_logic_vector(10998, 16),
30047 => conv_std_logic_vector(11115, 16),
30048 => conv_std_logic_vector(11232, 16),
30049 => conv_std_logic_vector(11349, 16),
30050 => conv_std_logic_vector(11466, 16),
30051 => conv_std_logic_vector(11583, 16),
30052 => conv_std_logic_vector(11700, 16),
30053 => conv_std_logic_vector(11817, 16),
30054 => conv_std_logic_vector(11934, 16),
30055 => conv_std_logic_vector(12051, 16),
30056 => conv_std_logic_vector(12168, 16),
30057 => conv_std_logic_vector(12285, 16),
30058 => conv_std_logic_vector(12402, 16),
30059 => conv_std_logic_vector(12519, 16),
30060 => conv_std_logic_vector(12636, 16),
30061 => conv_std_logic_vector(12753, 16),
30062 => conv_std_logic_vector(12870, 16),
30063 => conv_std_logic_vector(12987, 16),
30064 => conv_std_logic_vector(13104, 16),
30065 => conv_std_logic_vector(13221, 16),
30066 => conv_std_logic_vector(13338, 16),
30067 => conv_std_logic_vector(13455, 16),
30068 => conv_std_logic_vector(13572, 16),
30069 => conv_std_logic_vector(13689, 16),
30070 => conv_std_logic_vector(13806, 16),
30071 => conv_std_logic_vector(13923, 16),
30072 => conv_std_logic_vector(14040, 16),
30073 => conv_std_logic_vector(14157, 16),
30074 => conv_std_logic_vector(14274, 16),
30075 => conv_std_logic_vector(14391, 16),
30076 => conv_std_logic_vector(14508, 16),
30077 => conv_std_logic_vector(14625, 16),
30078 => conv_std_logic_vector(14742, 16),
30079 => conv_std_logic_vector(14859, 16),
30080 => conv_std_logic_vector(14976, 16),
30081 => conv_std_logic_vector(15093, 16),
30082 => conv_std_logic_vector(15210, 16),
30083 => conv_std_logic_vector(15327, 16),
30084 => conv_std_logic_vector(15444, 16),
30085 => conv_std_logic_vector(15561, 16),
30086 => conv_std_logic_vector(15678, 16),
30087 => conv_std_logic_vector(15795, 16),
30088 => conv_std_logic_vector(15912, 16),
30089 => conv_std_logic_vector(16029, 16),
30090 => conv_std_logic_vector(16146, 16),
30091 => conv_std_logic_vector(16263, 16),
30092 => conv_std_logic_vector(16380, 16),
30093 => conv_std_logic_vector(16497, 16),
30094 => conv_std_logic_vector(16614, 16),
30095 => conv_std_logic_vector(16731, 16),
30096 => conv_std_logic_vector(16848, 16),
30097 => conv_std_logic_vector(16965, 16),
30098 => conv_std_logic_vector(17082, 16),
30099 => conv_std_logic_vector(17199, 16),
30100 => conv_std_logic_vector(17316, 16),
30101 => conv_std_logic_vector(17433, 16),
30102 => conv_std_logic_vector(17550, 16),
30103 => conv_std_logic_vector(17667, 16),
30104 => conv_std_logic_vector(17784, 16),
30105 => conv_std_logic_vector(17901, 16),
30106 => conv_std_logic_vector(18018, 16),
30107 => conv_std_logic_vector(18135, 16),
30108 => conv_std_logic_vector(18252, 16),
30109 => conv_std_logic_vector(18369, 16),
30110 => conv_std_logic_vector(18486, 16),
30111 => conv_std_logic_vector(18603, 16),
30112 => conv_std_logic_vector(18720, 16),
30113 => conv_std_logic_vector(18837, 16),
30114 => conv_std_logic_vector(18954, 16),
30115 => conv_std_logic_vector(19071, 16),
30116 => conv_std_logic_vector(19188, 16),
30117 => conv_std_logic_vector(19305, 16),
30118 => conv_std_logic_vector(19422, 16),
30119 => conv_std_logic_vector(19539, 16),
30120 => conv_std_logic_vector(19656, 16),
30121 => conv_std_logic_vector(19773, 16),
30122 => conv_std_logic_vector(19890, 16),
30123 => conv_std_logic_vector(20007, 16),
30124 => conv_std_logic_vector(20124, 16),
30125 => conv_std_logic_vector(20241, 16),
30126 => conv_std_logic_vector(20358, 16),
30127 => conv_std_logic_vector(20475, 16),
30128 => conv_std_logic_vector(20592, 16),
30129 => conv_std_logic_vector(20709, 16),
30130 => conv_std_logic_vector(20826, 16),
30131 => conv_std_logic_vector(20943, 16),
30132 => conv_std_logic_vector(21060, 16),
30133 => conv_std_logic_vector(21177, 16),
30134 => conv_std_logic_vector(21294, 16),
30135 => conv_std_logic_vector(21411, 16),
30136 => conv_std_logic_vector(21528, 16),
30137 => conv_std_logic_vector(21645, 16),
30138 => conv_std_logic_vector(21762, 16),
30139 => conv_std_logic_vector(21879, 16),
30140 => conv_std_logic_vector(21996, 16),
30141 => conv_std_logic_vector(22113, 16),
30142 => conv_std_logic_vector(22230, 16),
30143 => conv_std_logic_vector(22347, 16),
30144 => conv_std_logic_vector(22464, 16),
30145 => conv_std_logic_vector(22581, 16),
30146 => conv_std_logic_vector(22698, 16),
30147 => conv_std_logic_vector(22815, 16),
30148 => conv_std_logic_vector(22932, 16),
30149 => conv_std_logic_vector(23049, 16),
30150 => conv_std_logic_vector(23166, 16),
30151 => conv_std_logic_vector(23283, 16),
30152 => conv_std_logic_vector(23400, 16),
30153 => conv_std_logic_vector(23517, 16),
30154 => conv_std_logic_vector(23634, 16),
30155 => conv_std_logic_vector(23751, 16),
30156 => conv_std_logic_vector(23868, 16),
30157 => conv_std_logic_vector(23985, 16),
30158 => conv_std_logic_vector(24102, 16),
30159 => conv_std_logic_vector(24219, 16),
30160 => conv_std_logic_vector(24336, 16),
30161 => conv_std_logic_vector(24453, 16),
30162 => conv_std_logic_vector(24570, 16),
30163 => conv_std_logic_vector(24687, 16),
30164 => conv_std_logic_vector(24804, 16),
30165 => conv_std_logic_vector(24921, 16),
30166 => conv_std_logic_vector(25038, 16),
30167 => conv_std_logic_vector(25155, 16),
30168 => conv_std_logic_vector(25272, 16),
30169 => conv_std_logic_vector(25389, 16),
30170 => conv_std_logic_vector(25506, 16),
30171 => conv_std_logic_vector(25623, 16),
30172 => conv_std_logic_vector(25740, 16),
30173 => conv_std_logic_vector(25857, 16),
30174 => conv_std_logic_vector(25974, 16),
30175 => conv_std_logic_vector(26091, 16),
30176 => conv_std_logic_vector(26208, 16),
30177 => conv_std_logic_vector(26325, 16),
30178 => conv_std_logic_vector(26442, 16),
30179 => conv_std_logic_vector(26559, 16),
30180 => conv_std_logic_vector(26676, 16),
30181 => conv_std_logic_vector(26793, 16),
30182 => conv_std_logic_vector(26910, 16),
30183 => conv_std_logic_vector(27027, 16),
30184 => conv_std_logic_vector(27144, 16),
30185 => conv_std_logic_vector(27261, 16),
30186 => conv_std_logic_vector(27378, 16),
30187 => conv_std_logic_vector(27495, 16),
30188 => conv_std_logic_vector(27612, 16),
30189 => conv_std_logic_vector(27729, 16),
30190 => conv_std_logic_vector(27846, 16),
30191 => conv_std_logic_vector(27963, 16),
30192 => conv_std_logic_vector(28080, 16),
30193 => conv_std_logic_vector(28197, 16),
30194 => conv_std_logic_vector(28314, 16),
30195 => conv_std_logic_vector(28431, 16),
30196 => conv_std_logic_vector(28548, 16),
30197 => conv_std_logic_vector(28665, 16),
30198 => conv_std_logic_vector(28782, 16),
30199 => conv_std_logic_vector(28899, 16),
30200 => conv_std_logic_vector(29016, 16),
30201 => conv_std_logic_vector(29133, 16),
30202 => conv_std_logic_vector(29250, 16),
30203 => conv_std_logic_vector(29367, 16),
30204 => conv_std_logic_vector(29484, 16),
30205 => conv_std_logic_vector(29601, 16),
30206 => conv_std_logic_vector(29718, 16),
30207 => conv_std_logic_vector(29835, 16),
30208 => conv_std_logic_vector(0, 16),
30209 => conv_std_logic_vector(118, 16),
30210 => conv_std_logic_vector(236, 16),
30211 => conv_std_logic_vector(354, 16),
30212 => conv_std_logic_vector(472, 16),
30213 => conv_std_logic_vector(590, 16),
30214 => conv_std_logic_vector(708, 16),
30215 => conv_std_logic_vector(826, 16),
30216 => conv_std_logic_vector(944, 16),
30217 => conv_std_logic_vector(1062, 16),
30218 => conv_std_logic_vector(1180, 16),
30219 => conv_std_logic_vector(1298, 16),
30220 => conv_std_logic_vector(1416, 16),
30221 => conv_std_logic_vector(1534, 16),
30222 => conv_std_logic_vector(1652, 16),
30223 => conv_std_logic_vector(1770, 16),
30224 => conv_std_logic_vector(1888, 16),
30225 => conv_std_logic_vector(2006, 16),
30226 => conv_std_logic_vector(2124, 16),
30227 => conv_std_logic_vector(2242, 16),
30228 => conv_std_logic_vector(2360, 16),
30229 => conv_std_logic_vector(2478, 16),
30230 => conv_std_logic_vector(2596, 16),
30231 => conv_std_logic_vector(2714, 16),
30232 => conv_std_logic_vector(2832, 16),
30233 => conv_std_logic_vector(2950, 16),
30234 => conv_std_logic_vector(3068, 16),
30235 => conv_std_logic_vector(3186, 16),
30236 => conv_std_logic_vector(3304, 16),
30237 => conv_std_logic_vector(3422, 16),
30238 => conv_std_logic_vector(3540, 16),
30239 => conv_std_logic_vector(3658, 16),
30240 => conv_std_logic_vector(3776, 16),
30241 => conv_std_logic_vector(3894, 16),
30242 => conv_std_logic_vector(4012, 16),
30243 => conv_std_logic_vector(4130, 16),
30244 => conv_std_logic_vector(4248, 16),
30245 => conv_std_logic_vector(4366, 16),
30246 => conv_std_logic_vector(4484, 16),
30247 => conv_std_logic_vector(4602, 16),
30248 => conv_std_logic_vector(4720, 16),
30249 => conv_std_logic_vector(4838, 16),
30250 => conv_std_logic_vector(4956, 16),
30251 => conv_std_logic_vector(5074, 16),
30252 => conv_std_logic_vector(5192, 16),
30253 => conv_std_logic_vector(5310, 16),
30254 => conv_std_logic_vector(5428, 16),
30255 => conv_std_logic_vector(5546, 16),
30256 => conv_std_logic_vector(5664, 16),
30257 => conv_std_logic_vector(5782, 16),
30258 => conv_std_logic_vector(5900, 16),
30259 => conv_std_logic_vector(6018, 16),
30260 => conv_std_logic_vector(6136, 16),
30261 => conv_std_logic_vector(6254, 16),
30262 => conv_std_logic_vector(6372, 16),
30263 => conv_std_logic_vector(6490, 16),
30264 => conv_std_logic_vector(6608, 16),
30265 => conv_std_logic_vector(6726, 16),
30266 => conv_std_logic_vector(6844, 16),
30267 => conv_std_logic_vector(6962, 16),
30268 => conv_std_logic_vector(7080, 16),
30269 => conv_std_logic_vector(7198, 16),
30270 => conv_std_logic_vector(7316, 16),
30271 => conv_std_logic_vector(7434, 16),
30272 => conv_std_logic_vector(7552, 16),
30273 => conv_std_logic_vector(7670, 16),
30274 => conv_std_logic_vector(7788, 16),
30275 => conv_std_logic_vector(7906, 16),
30276 => conv_std_logic_vector(8024, 16),
30277 => conv_std_logic_vector(8142, 16),
30278 => conv_std_logic_vector(8260, 16),
30279 => conv_std_logic_vector(8378, 16),
30280 => conv_std_logic_vector(8496, 16),
30281 => conv_std_logic_vector(8614, 16),
30282 => conv_std_logic_vector(8732, 16),
30283 => conv_std_logic_vector(8850, 16),
30284 => conv_std_logic_vector(8968, 16),
30285 => conv_std_logic_vector(9086, 16),
30286 => conv_std_logic_vector(9204, 16),
30287 => conv_std_logic_vector(9322, 16),
30288 => conv_std_logic_vector(9440, 16),
30289 => conv_std_logic_vector(9558, 16),
30290 => conv_std_logic_vector(9676, 16),
30291 => conv_std_logic_vector(9794, 16),
30292 => conv_std_logic_vector(9912, 16),
30293 => conv_std_logic_vector(10030, 16),
30294 => conv_std_logic_vector(10148, 16),
30295 => conv_std_logic_vector(10266, 16),
30296 => conv_std_logic_vector(10384, 16),
30297 => conv_std_logic_vector(10502, 16),
30298 => conv_std_logic_vector(10620, 16),
30299 => conv_std_logic_vector(10738, 16),
30300 => conv_std_logic_vector(10856, 16),
30301 => conv_std_logic_vector(10974, 16),
30302 => conv_std_logic_vector(11092, 16),
30303 => conv_std_logic_vector(11210, 16),
30304 => conv_std_logic_vector(11328, 16),
30305 => conv_std_logic_vector(11446, 16),
30306 => conv_std_logic_vector(11564, 16),
30307 => conv_std_logic_vector(11682, 16),
30308 => conv_std_logic_vector(11800, 16),
30309 => conv_std_logic_vector(11918, 16),
30310 => conv_std_logic_vector(12036, 16),
30311 => conv_std_logic_vector(12154, 16),
30312 => conv_std_logic_vector(12272, 16),
30313 => conv_std_logic_vector(12390, 16),
30314 => conv_std_logic_vector(12508, 16),
30315 => conv_std_logic_vector(12626, 16),
30316 => conv_std_logic_vector(12744, 16),
30317 => conv_std_logic_vector(12862, 16),
30318 => conv_std_logic_vector(12980, 16),
30319 => conv_std_logic_vector(13098, 16),
30320 => conv_std_logic_vector(13216, 16),
30321 => conv_std_logic_vector(13334, 16),
30322 => conv_std_logic_vector(13452, 16),
30323 => conv_std_logic_vector(13570, 16),
30324 => conv_std_logic_vector(13688, 16),
30325 => conv_std_logic_vector(13806, 16),
30326 => conv_std_logic_vector(13924, 16),
30327 => conv_std_logic_vector(14042, 16),
30328 => conv_std_logic_vector(14160, 16),
30329 => conv_std_logic_vector(14278, 16),
30330 => conv_std_logic_vector(14396, 16),
30331 => conv_std_logic_vector(14514, 16),
30332 => conv_std_logic_vector(14632, 16),
30333 => conv_std_logic_vector(14750, 16),
30334 => conv_std_logic_vector(14868, 16),
30335 => conv_std_logic_vector(14986, 16),
30336 => conv_std_logic_vector(15104, 16),
30337 => conv_std_logic_vector(15222, 16),
30338 => conv_std_logic_vector(15340, 16),
30339 => conv_std_logic_vector(15458, 16),
30340 => conv_std_logic_vector(15576, 16),
30341 => conv_std_logic_vector(15694, 16),
30342 => conv_std_logic_vector(15812, 16),
30343 => conv_std_logic_vector(15930, 16),
30344 => conv_std_logic_vector(16048, 16),
30345 => conv_std_logic_vector(16166, 16),
30346 => conv_std_logic_vector(16284, 16),
30347 => conv_std_logic_vector(16402, 16),
30348 => conv_std_logic_vector(16520, 16),
30349 => conv_std_logic_vector(16638, 16),
30350 => conv_std_logic_vector(16756, 16),
30351 => conv_std_logic_vector(16874, 16),
30352 => conv_std_logic_vector(16992, 16),
30353 => conv_std_logic_vector(17110, 16),
30354 => conv_std_logic_vector(17228, 16),
30355 => conv_std_logic_vector(17346, 16),
30356 => conv_std_logic_vector(17464, 16),
30357 => conv_std_logic_vector(17582, 16),
30358 => conv_std_logic_vector(17700, 16),
30359 => conv_std_logic_vector(17818, 16),
30360 => conv_std_logic_vector(17936, 16),
30361 => conv_std_logic_vector(18054, 16),
30362 => conv_std_logic_vector(18172, 16),
30363 => conv_std_logic_vector(18290, 16),
30364 => conv_std_logic_vector(18408, 16),
30365 => conv_std_logic_vector(18526, 16),
30366 => conv_std_logic_vector(18644, 16),
30367 => conv_std_logic_vector(18762, 16),
30368 => conv_std_logic_vector(18880, 16),
30369 => conv_std_logic_vector(18998, 16),
30370 => conv_std_logic_vector(19116, 16),
30371 => conv_std_logic_vector(19234, 16),
30372 => conv_std_logic_vector(19352, 16),
30373 => conv_std_logic_vector(19470, 16),
30374 => conv_std_logic_vector(19588, 16),
30375 => conv_std_logic_vector(19706, 16),
30376 => conv_std_logic_vector(19824, 16),
30377 => conv_std_logic_vector(19942, 16),
30378 => conv_std_logic_vector(20060, 16),
30379 => conv_std_logic_vector(20178, 16),
30380 => conv_std_logic_vector(20296, 16),
30381 => conv_std_logic_vector(20414, 16),
30382 => conv_std_logic_vector(20532, 16),
30383 => conv_std_logic_vector(20650, 16),
30384 => conv_std_logic_vector(20768, 16),
30385 => conv_std_logic_vector(20886, 16),
30386 => conv_std_logic_vector(21004, 16),
30387 => conv_std_logic_vector(21122, 16),
30388 => conv_std_logic_vector(21240, 16),
30389 => conv_std_logic_vector(21358, 16),
30390 => conv_std_logic_vector(21476, 16),
30391 => conv_std_logic_vector(21594, 16),
30392 => conv_std_logic_vector(21712, 16),
30393 => conv_std_logic_vector(21830, 16),
30394 => conv_std_logic_vector(21948, 16),
30395 => conv_std_logic_vector(22066, 16),
30396 => conv_std_logic_vector(22184, 16),
30397 => conv_std_logic_vector(22302, 16),
30398 => conv_std_logic_vector(22420, 16),
30399 => conv_std_logic_vector(22538, 16),
30400 => conv_std_logic_vector(22656, 16),
30401 => conv_std_logic_vector(22774, 16),
30402 => conv_std_logic_vector(22892, 16),
30403 => conv_std_logic_vector(23010, 16),
30404 => conv_std_logic_vector(23128, 16),
30405 => conv_std_logic_vector(23246, 16),
30406 => conv_std_logic_vector(23364, 16),
30407 => conv_std_logic_vector(23482, 16),
30408 => conv_std_logic_vector(23600, 16),
30409 => conv_std_logic_vector(23718, 16),
30410 => conv_std_logic_vector(23836, 16),
30411 => conv_std_logic_vector(23954, 16),
30412 => conv_std_logic_vector(24072, 16),
30413 => conv_std_logic_vector(24190, 16),
30414 => conv_std_logic_vector(24308, 16),
30415 => conv_std_logic_vector(24426, 16),
30416 => conv_std_logic_vector(24544, 16),
30417 => conv_std_logic_vector(24662, 16),
30418 => conv_std_logic_vector(24780, 16),
30419 => conv_std_logic_vector(24898, 16),
30420 => conv_std_logic_vector(25016, 16),
30421 => conv_std_logic_vector(25134, 16),
30422 => conv_std_logic_vector(25252, 16),
30423 => conv_std_logic_vector(25370, 16),
30424 => conv_std_logic_vector(25488, 16),
30425 => conv_std_logic_vector(25606, 16),
30426 => conv_std_logic_vector(25724, 16),
30427 => conv_std_logic_vector(25842, 16),
30428 => conv_std_logic_vector(25960, 16),
30429 => conv_std_logic_vector(26078, 16),
30430 => conv_std_logic_vector(26196, 16),
30431 => conv_std_logic_vector(26314, 16),
30432 => conv_std_logic_vector(26432, 16),
30433 => conv_std_logic_vector(26550, 16),
30434 => conv_std_logic_vector(26668, 16),
30435 => conv_std_logic_vector(26786, 16),
30436 => conv_std_logic_vector(26904, 16),
30437 => conv_std_logic_vector(27022, 16),
30438 => conv_std_logic_vector(27140, 16),
30439 => conv_std_logic_vector(27258, 16),
30440 => conv_std_logic_vector(27376, 16),
30441 => conv_std_logic_vector(27494, 16),
30442 => conv_std_logic_vector(27612, 16),
30443 => conv_std_logic_vector(27730, 16),
30444 => conv_std_logic_vector(27848, 16),
30445 => conv_std_logic_vector(27966, 16),
30446 => conv_std_logic_vector(28084, 16),
30447 => conv_std_logic_vector(28202, 16),
30448 => conv_std_logic_vector(28320, 16),
30449 => conv_std_logic_vector(28438, 16),
30450 => conv_std_logic_vector(28556, 16),
30451 => conv_std_logic_vector(28674, 16),
30452 => conv_std_logic_vector(28792, 16),
30453 => conv_std_logic_vector(28910, 16),
30454 => conv_std_logic_vector(29028, 16),
30455 => conv_std_logic_vector(29146, 16),
30456 => conv_std_logic_vector(29264, 16),
30457 => conv_std_logic_vector(29382, 16),
30458 => conv_std_logic_vector(29500, 16),
30459 => conv_std_logic_vector(29618, 16),
30460 => conv_std_logic_vector(29736, 16),
30461 => conv_std_logic_vector(29854, 16),
30462 => conv_std_logic_vector(29972, 16),
30463 => conv_std_logic_vector(30090, 16),
30464 => conv_std_logic_vector(0, 16),
30465 => conv_std_logic_vector(119, 16),
30466 => conv_std_logic_vector(238, 16),
30467 => conv_std_logic_vector(357, 16),
30468 => conv_std_logic_vector(476, 16),
30469 => conv_std_logic_vector(595, 16),
30470 => conv_std_logic_vector(714, 16),
30471 => conv_std_logic_vector(833, 16),
30472 => conv_std_logic_vector(952, 16),
30473 => conv_std_logic_vector(1071, 16),
30474 => conv_std_logic_vector(1190, 16),
30475 => conv_std_logic_vector(1309, 16),
30476 => conv_std_logic_vector(1428, 16),
30477 => conv_std_logic_vector(1547, 16),
30478 => conv_std_logic_vector(1666, 16),
30479 => conv_std_logic_vector(1785, 16),
30480 => conv_std_logic_vector(1904, 16),
30481 => conv_std_logic_vector(2023, 16),
30482 => conv_std_logic_vector(2142, 16),
30483 => conv_std_logic_vector(2261, 16),
30484 => conv_std_logic_vector(2380, 16),
30485 => conv_std_logic_vector(2499, 16),
30486 => conv_std_logic_vector(2618, 16),
30487 => conv_std_logic_vector(2737, 16),
30488 => conv_std_logic_vector(2856, 16),
30489 => conv_std_logic_vector(2975, 16),
30490 => conv_std_logic_vector(3094, 16),
30491 => conv_std_logic_vector(3213, 16),
30492 => conv_std_logic_vector(3332, 16),
30493 => conv_std_logic_vector(3451, 16),
30494 => conv_std_logic_vector(3570, 16),
30495 => conv_std_logic_vector(3689, 16),
30496 => conv_std_logic_vector(3808, 16),
30497 => conv_std_logic_vector(3927, 16),
30498 => conv_std_logic_vector(4046, 16),
30499 => conv_std_logic_vector(4165, 16),
30500 => conv_std_logic_vector(4284, 16),
30501 => conv_std_logic_vector(4403, 16),
30502 => conv_std_logic_vector(4522, 16),
30503 => conv_std_logic_vector(4641, 16),
30504 => conv_std_logic_vector(4760, 16),
30505 => conv_std_logic_vector(4879, 16),
30506 => conv_std_logic_vector(4998, 16),
30507 => conv_std_logic_vector(5117, 16),
30508 => conv_std_logic_vector(5236, 16),
30509 => conv_std_logic_vector(5355, 16),
30510 => conv_std_logic_vector(5474, 16),
30511 => conv_std_logic_vector(5593, 16),
30512 => conv_std_logic_vector(5712, 16),
30513 => conv_std_logic_vector(5831, 16),
30514 => conv_std_logic_vector(5950, 16),
30515 => conv_std_logic_vector(6069, 16),
30516 => conv_std_logic_vector(6188, 16),
30517 => conv_std_logic_vector(6307, 16),
30518 => conv_std_logic_vector(6426, 16),
30519 => conv_std_logic_vector(6545, 16),
30520 => conv_std_logic_vector(6664, 16),
30521 => conv_std_logic_vector(6783, 16),
30522 => conv_std_logic_vector(6902, 16),
30523 => conv_std_logic_vector(7021, 16),
30524 => conv_std_logic_vector(7140, 16),
30525 => conv_std_logic_vector(7259, 16),
30526 => conv_std_logic_vector(7378, 16),
30527 => conv_std_logic_vector(7497, 16),
30528 => conv_std_logic_vector(7616, 16),
30529 => conv_std_logic_vector(7735, 16),
30530 => conv_std_logic_vector(7854, 16),
30531 => conv_std_logic_vector(7973, 16),
30532 => conv_std_logic_vector(8092, 16),
30533 => conv_std_logic_vector(8211, 16),
30534 => conv_std_logic_vector(8330, 16),
30535 => conv_std_logic_vector(8449, 16),
30536 => conv_std_logic_vector(8568, 16),
30537 => conv_std_logic_vector(8687, 16),
30538 => conv_std_logic_vector(8806, 16),
30539 => conv_std_logic_vector(8925, 16),
30540 => conv_std_logic_vector(9044, 16),
30541 => conv_std_logic_vector(9163, 16),
30542 => conv_std_logic_vector(9282, 16),
30543 => conv_std_logic_vector(9401, 16),
30544 => conv_std_logic_vector(9520, 16),
30545 => conv_std_logic_vector(9639, 16),
30546 => conv_std_logic_vector(9758, 16),
30547 => conv_std_logic_vector(9877, 16),
30548 => conv_std_logic_vector(9996, 16),
30549 => conv_std_logic_vector(10115, 16),
30550 => conv_std_logic_vector(10234, 16),
30551 => conv_std_logic_vector(10353, 16),
30552 => conv_std_logic_vector(10472, 16),
30553 => conv_std_logic_vector(10591, 16),
30554 => conv_std_logic_vector(10710, 16),
30555 => conv_std_logic_vector(10829, 16),
30556 => conv_std_logic_vector(10948, 16),
30557 => conv_std_logic_vector(11067, 16),
30558 => conv_std_logic_vector(11186, 16),
30559 => conv_std_logic_vector(11305, 16),
30560 => conv_std_logic_vector(11424, 16),
30561 => conv_std_logic_vector(11543, 16),
30562 => conv_std_logic_vector(11662, 16),
30563 => conv_std_logic_vector(11781, 16),
30564 => conv_std_logic_vector(11900, 16),
30565 => conv_std_logic_vector(12019, 16),
30566 => conv_std_logic_vector(12138, 16),
30567 => conv_std_logic_vector(12257, 16),
30568 => conv_std_logic_vector(12376, 16),
30569 => conv_std_logic_vector(12495, 16),
30570 => conv_std_logic_vector(12614, 16),
30571 => conv_std_logic_vector(12733, 16),
30572 => conv_std_logic_vector(12852, 16),
30573 => conv_std_logic_vector(12971, 16),
30574 => conv_std_logic_vector(13090, 16),
30575 => conv_std_logic_vector(13209, 16),
30576 => conv_std_logic_vector(13328, 16),
30577 => conv_std_logic_vector(13447, 16),
30578 => conv_std_logic_vector(13566, 16),
30579 => conv_std_logic_vector(13685, 16),
30580 => conv_std_logic_vector(13804, 16),
30581 => conv_std_logic_vector(13923, 16),
30582 => conv_std_logic_vector(14042, 16),
30583 => conv_std_logic_vector(14161, 16),
30584 => conv_std_logic_vector(14280, 16),
30585 => conv_std_logic_vector(14399, 16),
30586 => conv_std_logic_vector(14518, 16),
30587 => conv_std_logic_vector(14637, 16),
30588 => conv_std_logic_vector(14756, 16),
30589 => conv_std_logic_vector(14875, 16),
30590 => conv_std_logic_vector(14994, 16),
30591 => conv_std_logic_vector(15113, 16),
30592 => conv_std_logic_vector(15232, 16),
30593 => conv_std_logic_vector(15351, 16),
30594 => conv_std_logic_vector(15470, 16),
30595 => conv_std_logic_vector(15589, 16),
30596 => conv_std_logic_vector(15708, 16),
30597 => conv_std_logic_vector(15827, 16),
30598 => conv_std_logic_vector(15946, 16),
30599 => conv_std_logic_vector(16065, 16),
30600 => conv_std_logic_vector(16184, 16),
30601 => conv_std_logic_vector(16303, 16),
30602 => conv_std_logic_vector(16422, 16),
30603 => conv_std_logic_vector(16541, 16),
30604 => conv_std_logic_vector(16660, 16),
30605 => conv_std_logic_vector(16779, 16),
30606 => conv_std_logic_vector(16898, 16),
30607 => conv_std_logic_vector(17017, 16),
30608 => conv_std_logic_vector(17136, 16),
30609 => conv_std_logic_vector(17255, 16),
30610 => conv_std_logic_vector(17374, 16),
30611 => conv_std_logic_vector(17493, 16),
30612 => conv_std_logic_vector(17612, 16),
30613 => conv_std_logic_vector(17731, 16),
30614 => conv_std_logic_vector(17850, 16),
30615 => conv_std_logic_vector(17969, 16),
30616 => conv_std_logic_vector(18088, 16),
30617 => conv_std_logic_vector(18207, 16),
30618 => conv_std_logic_vector(18326, 16),
30619 => conv_std_logic_vector(18445, 16),
30620 => conv_std_logic_vector(18564, 16),
30621 => conv_std_logic_vector(18683, 16),
30622 => conv_std_logic_vector(18802, 16),
30623 => conv_std_logic_vector(18921, 16),
30624 => conv_std_logic_vector(19040, 16),
30625 => conv_std_logic_vector(19159, 16),
30626 => conv_std_logic_vector(19278, 16),
30627 => conv_std_logic_vector(19397, 16),
30628 => conv_std_logic_vector(19516, 16),
30629 => conv_std_logic_vector(19635, 16),
30630 => conv_std_logic_vector(19754, 16),
30631 => conv_std_logic_vector(19873, 16),
30632 => conv_std_logic_vector(19992, 16),
30633 => conv_std_logic_vector(20111, 16),
30634 => conv_std_logic_vector(20230, 16),
30635 => conv_std_logic_vector(20349, 16),
30636 => conv_std_logic_vector(20468, 16),
30637 => conv_std_logic_vector(20587, 16),
30638 => conv_std_logic_vector(20706, 16),
30639 => conv_std_logic_vector(20825, 16),
30640 => conv_std_logic_vector(20944, 16),
30641 => conv_std_logic_vector(21063, 16),
30642 => conv_std_logic_vector(21182, 16),
30643 => conv_std_logic_vector(21301, 16),
30644 => conv_std_logic_vector(21420, 16),
30645 => conv_std_logic_vector(21539, 16),
30646 => conv_std_logic_vector(21658, 16),
30647 => conv_std_logic_vector(21777, 16),
30648 => conv_std_logic_vector(21896, 16),
30649 => conv_std_logic_vector(22015, 16),
30650 => conv_std_logic_vector(22134, 16),
30651 => conv_std_logic_vector(22253, 16),
30652 => conv_std_logic_vector(22372, 16),
30653 => conv_std_logic_vector(22491, 16),
30654 => conv_std_logic_vector(22610, 16),
30655 => conv_std_logic_vector(22729, 16),
30656 => conv_std_logic_vector(22848, 16),
30657 => conv_std_logic_vector(22967, 16),
30658 => conv_std_logic_vector(23086, 16),
30659 => conv_std_logic_vector(23205, 16),
30660 => conv_std_logic_vector(23324, 16),
30661 => conv_std_logic_vector(23443, 16),
30662 => conv_std_logic_vector(23562, 16),
30663 => conv_std_logic_vector(23681, 16),
30664 => conv_std_logic_vector(23800, 16),
30665 => conv_std_logic_vector(23919, 16),
30666 => conv_std_logic_vector(24038, 16),
30667 => conv_std_logic_vector(24157, 16),
30668 => conv_std_logic_vector(24276, 16),
30669 => conv_std_logic_vector(24395, 16),
30670 => conv_std_logic_vector(24514, 16),
30671 => conv_std_logic_vector(24633, 16),
30672 => conv_std_logic_vector(24752, 16),
30673 => conv_std_logic_vector(24871, 16),
30674 => conv_std_logic_vector(24990, 16),
30675 => conv_std_logic_vector(25109, 16),
30676 => conv_std_logic_vector(25228, 16),
30677 => conv_std_logic_vector(25347, 16),
30678 => conv_std_logic_vector(25466, 16),
30679 => conv_std_logic_vector(25585, 16),
30680 => conv_std_logic_vector(25704, 16),
30681 => conv_std_logic_vector(25823, 16),
30682 => conv_std_logic_vector(25942, 16),
30683 => conv_std_logic_vector(26061, 16),
30684 => conv_std_logic_vector(26180, 16),
30685 => conv_std_logic_vector(26299, 16),
30686 => conv_std_logic_vector(26418, 16),
30687 => conv_std_logic_vector(26537, 16),
30688 => conv_std_logic_vector(26656, 16),
30689 => conv_std_logic_vector(26775, 16),
30690 => conv_std_logic_vector(26894, 16),
30691 => conv_std_logic_vector(27013, 16),
30692 => conv_std_logic_vector(27132, 16),
30693 => conv_std_logic_vector(27251, 16),
30694 => conv_std_logic_vector(27370, 16),
30695 => conv_std_logic_vector(27489, 16),
30696 => conv_std_logic_vector(27608, 16),
30697 => conv_std_logic_vector(27727, 16),
30698 => conv_std_logic_vector(27846, 16),
30699 => conv_std_logic_vector(27965, 16),
30700 => conv_std_logic_vector(28084, 16),
30701 => conv_std_logic_vector(28203, 16),
30702 => conv_std_logic_vector(28322, 16),
30703 => conv_std_logic_vector(28441, 16),
30704 => conv_std_logic_vector(28560, 16),
30705 => conv_std_logic_vector(28679, 16),
30706 => conv_std_logic_vector(28798, 16),
30707 => conv_std_logic_vector(28917, 16),
30708 => conv_std_logic_vector(29036, 16),
30709 => conv_std_logic_vector(29155, 16),
30710 => conv_std_logic_vector(29274, 16),
30711 => conv_std_logic_vector(29393, 16),
30712 => conv_std_logic_vector(29512, 16),
30713 => conv_std_logic_vector(29631, 16),
30714 => conv_std_logic_vector(29750, 16),
30715 => conv_std_logic_vector(29869, 16),
30716 => conv_std_logic_vector(29988, 16),
30717 => conv_std_logic_vector(30107, 16),
30718 => conv_std_logic_vector(30226, 16),
30719 => conv_std_logic_vector(30345, 16),
30720 => conv_std_logic_vector(0, 16),
30721 => conv_std_logic_vector(120, 16),
30722 => conv_std_logic_vector(240, 16),
30723 => conv_std_logic_vector(360, 16),
30724 => conv_std_logic_vector(480, 16),
30725 => conv_std_logic_vector(600, 16),
30726 => conv_std_logic_vector(720, 16),
30727 => conv_std_logic_vector(840, 16),
30728 => conv_std_logic_vector(960, 16),
30729 => conv_std_logic_vector(1080, 16),
30730 => conv_std_logic_vector(1200, 16),
30731 => conv_std_logic_vector(1320, 16),
30732 => conv_std_logic_vector(1440, 16),
30733 => conv_std_logic_vector(1560, 16),
30734 => conv_std_logic_vector(1680, 16),
30735 => conv_std_logic_vector(1800, 16),
30736 => conv_std_logic_vector(1920, 16),
30737 => conv_std_logic_vector(2040, 16),
30738 => conv_std_logic_vector(2160, 16),
30739 => conv_std_logic_vector(2280, 16),
30740 => conv_std_logic_vector(2400, 16),
30741 => conv_std_logic_vector(2520, 16),
30742 => conv_std_logic_vector(2640, 16),
30743 => conv_std_logic_vector(2760, 16),
30744 => conv_std_logic_vector(2880, 16),
30745 => conv_std_logic_vector(3000, 16),
30746 => conv_std_logic_vector(3120, 16),
30747 => conv_std_logic_vector(3240, 16),
30748 => conv_std_logic_vector(3360, 16),
30749 => conv_std_logic_vector(3480, 16),
30750 => conv_std_logic_vector(3600, 16),
30751 => conv_std_logic_vector(3720, 16),
30752 => conv_std_logic_vector(3840, 16),
30753 => conv_std_logic_vector(3960, 16),
30754 => conv_std_logic_vector(4080, 16),
30755 => conv_std_logic_vector(4200, 16),
30756 => conv_std_logic_vector(4320, 16),
30757 => conv_std_logic_vector(4440, 16),
30758 => conv_std_logic_vector(4560, 16),
30759 => conv_std_logic_vector(4680, 16),
30760 => conv_std_logic_vector(4800, 16),
30761 => conv_std_logic_vector(4920, 16),
30762 => conv_std_logic_vector(5040, 16),
30763 => conv_std_logic_vector(5160, 16),
30764 => conv_std_logic_vector(5280, 16),
30765 => conv_std_logic_vector(5400, 16),
30766 => conv_std_logic_vector(5520, 16),
30767 => conv_std_logic_vector(5640, 16),
30768 => conv_std_logic_vector(5760, 16),
30769 => conv_std_logic_vector(5880, 16),
30770 => conv_std_logic_vector(6000, 16),
30771 => conv_std_logic_vector(6120, 16),
30772 => conv_std_logic_vector(6240, 16),
30773 => conv_std_logic_vector(6360, 16),
30774 => conv_std_logic_vector(6480, 16),
30775 => conv_std_logic_vector(6600, 16),
30776 => conv_std_logic_vector(6720, 16),
30777 => conv_std_logic_vector(6840, 16),
30778 => conv_std_logic_vector(6960, 16),
30779 => conv_std_logic_vector(7080, 16),
30780 => conv_std_logic_vector(7200, 16),
30781 => conv_std_logic_vector(7320, 16),
30782 => conv_std_logic_vector(7440, 16),
30783 => conv_std_logic_vector(7560, 16),
30784 => conv_std_logic_vector(7680, 16),
30785 => conv_std_logic_vector(7800, 16),
30786 => conv_std_logic_vector(7920, 16),
30787 => conv_std_logic_vector(8040, 16),
30788 => conv_std_logic_vector(8160, 16),
30789 => conv_std_logic_vector(8280, 16),
30790 => conv_std_logic_vector(8400, 16),
30791 => conv_std_logic_vector(8520, 16),
30792 => conv_std_logic_vector(8640, 16),
30793 => conv_std_logic_vector(8760, 16),
30794 => conv_std_logic_vector(8880, 16),
30795 => conv_std_logic_vector(9000, 16),
30796 => conv_std_logic_vector(9120, 16),
30797 => conv_std_logic_vector(9240, 16),
30798 => conv_std_logic_vector(9360, 16),
30799 => conv_std_logic_vector(9480, 16),
30800 => conv_std_logic_vector(9600, 16),
30801 => conv_std_logic_vector(9720, 16),
30802 => conv_std_logic_vector(9840, 16),
30803 => conv_std_logic_vector(9960, 16),
30804 => conv_std_logic_vector(10080, 16),
30805 => conv_std_logic_vector(10200, 16),
30806 => conv_std_logic_vector(10320, 16),
30807 => conv_std_logic_vector(10440, 16),
30808 => conv_std_logic_vector(10560, 16),
30809 => conv_std_logic_vector(10680, 16),
30810 => conv_std_logic_vector(10800, 16),
30811 => conv_std_logic_vector(10920, 16),
30812 => conv_std_logic_vector(11040, 16),
30813 => conv_std_logic_vector(11160, 16),
30814 => conv_std_logic_vector(11280, 16),
30815 => conv_std_logic_vector(11400, 16),
30816 => conv_std_logic_vector(11520, 16),
30817 => conv_std_logic_vector(11640, 16),
30818 => conv_std_logic_vector(11760, 16),
30819 => conv_std_logic_vector(11880, 16),
30820 => conv_std_logic_vector(12000, 16),
30821 => conv_std_logic_vector(12120, 16),
30822 => conv_std_logic_vector(12240, 16),
30823 => conv_std_logic_vector(12360, 16),
30824 => conv_std_logic_vector(12480, 16),
30825 => conv_std_logic_vector(12600, 16),
30826 => conv_std_logic_vector(12720, 16),
30827 => conv_std_logic_vector(12840, 16),
30828 => conv_std_logic_vector(12960, 16),
30829 => conv_std_logic_vector(13080, 16),
30830 => conv_std_logic_vector(13200, 16),
30831 => conv_std_logic_vector(13320, 16),
30832 => conv_std_logic_vector(13440, 16),
30833 => conv_std_logic_vector(13560, 16),
30834 => conv_std_logic_vector(13680, 16),
30835 => conv_std_logic_vector(13800, 16),
30836 => conv_std_logic_vector(13920, 16),
30837 => conv_std_logic_vector(14040, 16),
30838 => conv_std_logic_vector(14160, 16),
30839 => conv_std_logic_vector(14280, 16),
30840 => conv_std_logic_vector(14400, 16),
30841 => conv_std_logic_vector(14520, 16),
30842 => conv_std_logic_vector(14640, 16),
30843 => conv_std_logic_vector(14760, 16),
30844 => conv_std_logic_vector(14880, 16),
30845 => conv_std_logic_vector(15000, 16),
30846 => conv_std_logic_vector(15120, 16),
30847 => conv_std_logic_vector(15240, 16),
30848 => conv_std_logic_vector(15360, 16),
30849 => conv_std_logic_vector(15480, 16),
30850 => conv_std_logic_vector(15600, 16),
30851 => conv_std_logic_vector(15720, 16),
30852 => conv_std_logic_vector(15840, 16),
30853 => conv_std_logic_vector(15960, 16),
30854 => conv_std_logic_vector(16080, 16),
30855 => conv_std_logic_vector(16200, 16),
30856 => conv_std_logic_vector(16320, 16),
30857 => conv_std_logic_vector(16440, 16),
30858 => conv_std_logic_vector(16560, 16),
30859 => conv_std_logic_vector(16680, 16),
30860 => conv_std_logic_vector(16800, 16),
30861 => conv_std_logic_vector(16920, 16),
30862 => conv_std_logic_vector(17040, 16),
30863 => conv_std_logic_vector(17160, 16),
30864 => conv_std_logic_vector(17280, 16),
30865 => conv_std_logic_vector(17400, 16),
30866 => conv_std_logic_vector(17520, 16),
30867 => conv_std_logic_vector(17640, 16),
30868 => conv_std_logic_vector(17760, 16),
30869 => conv_std_logic_vector(17880, 16),
30870 => conv_std_logic_vector(18000, 16),
30871 => conv_std_logic_vector(18120, 16),
30872 => conv_std_logic_vector(18240, 16),
30873 => conv_std_logic_vector(18360, 16),
30874 => conv_std_logic_vector(18480, 16),
30875 => conv_std_logic_vector(18600, 16),
30876 => conv_std_logic_vector(18720, 16),
30877 => conv_std_logic_vector(18840, 16),
30878 => conv_std_logic_vector(18960, 16),
30879 => conv_std_logic_vector(19080, 16),
30880 => conv_std_logic_vector(19200, 16),
30881 => conv_std_logic_vector(19320, 16),
30882 => conv_std_logic_vector(19440, 16),
30883 => conv_std_logic_vector(19560, 16),
30884 => conv_std_logic_vector(19680, 16),
30885 => conv_std_logic_vector(19800, 16),
30886 => conv_std_logic_vector(19920, 16),
30887 => conv_std_logic_vector(20040, 16),
30888 => conv_std_logic_vector(20160, 16),
30889 => conv_std_logic_vector(20280, 16),
30890 => conv_std_logic_vector(20400, 16),
30891 => conv_std_logic_vector(20520, 16),
30892 => conv_std_logic_vector(20640, 16),
30893 => conv_std_logic_vector(20760, 16),
30894 => conv_std_logic_vector(20880, 16),
30895 => conv_std_logic_vector(21000, 16),
30896 => conv_std_logic_vector(21120, 16),
30897 => conv_std_logic_vector(21240, 16),
30898 => conv_std_logic_vector(21360, 16),
30899 => conv_std_logic_vector(21480, 16),
30900 => conv_std_logic_vector(21600, 16),
30901 => conv_std_logic_vector(21720, 16),
30902 => conv_std_logic_vector(21840, 16),
30903 => conv_std_logic_vector(21960, 16),
30904 => conv_std_logic_vector(22080, 16),
30905 => conv_std_logic_vector(22200, 16),
30906 => conv_std_logic_vector(22320, 16),
30907 => conv_std_logic_vector(22440, 16),
30908 => conv_std_logic_vector(22560, 16),
30909 => conv_std_logic_vector(22680, 16),
30910 => conv_std_logic_vector(22800, 16),
30911 => conv_std_logic_vector(22920, 16),
30912 => conv_std_logic_vector(23040, 16),
30913 => conv_std_logic_vector(23160, 16),
30914 => conv_std_logic_vector(23280, 16),
30915 => conv_std_logic_vector(23400, 16),
30916 => conv_std_logic_vector(23520, 16),
30917 => conv_std_logic_vector(23640, 16),
30918 => conv_std_logic_vector(23760, 16),
30919 => conv_std_logic_vector(23880, 16),
30920 => conv_std_logic_vector(24000, 16),
30921 => conv_std_logic_vector(24120, 16),
30922 => conv_std_logic_vector(24240, 16),
30923 => conv_std_logic_vector(24360, 16),
30924 => conv_std_logic_vector(24480, 16),
30925 => conv_std_logic_vector(24600, 16),
30926 => conv_std_logic_vector(24720, 16),
30927 => conv_std_logic_vector(24840, 16),
30928 => conv_std_logic_vector(24960, 16),
30929 => conv_std_logic_vector(25080, 16),
30930 => conv_std_logic_vector(25200, 16),
30931 => conv_std_logic_vector(25320, 16),
30932 => conv_std_logic_vector(25440, 16),
30933 => conv_std_logic_vector(25560, 16),
30934 => conv_std_logic_vector(25680, 16),
30935 => conv_std_logic_vector(25800, 16),
30936 => conv_std_logic_vector(25920, 16),
30937 => conv_std_logic_vector(26040, 16),
30938 => conv_std_logic_vector(26160, 16),
30939 => conv_std_logic_vector(26280, 16),
30940 => conv_std_logic_vector(26400, 16),
30941 => conv_std_logic_vector(26520, 16),
30942 => conv_std_logic_vector(26640, 16),
30943 => conv_std_logic_vector(26760, 16),
30944 => conv_std_logic_vector(26880, 16),
30945 => conv_std_logic_vector(27000, 16),
30946 => conv_std_logic_vector(27120, 16),
30947 => conv_std_logic_vector(27240, 16),
30948 => conv_std_logic_vector(27360, 16),
30949 => conv_std_logic_vector(27480, 16),
30950 => conv_std_logic_vector(27600, 16),
30951 => conv_std_logic_vector(27720, 16),
30952 => conv_std_logic_vector(27840, 16),
30953 => conv_std_logic_vector(27960, 16),
30954 => conv_std_logic_vector(28080, 16),
30955 => conv_std_logic_vector(28200, 16),
30956 => conv_std_logic_vector(28320, 16),
30957 => conv_std_logic_vector(28440, 16),
30958 => conv_std_logic_vector(28560, 16),
30959 => conv_std_logic_vector(28680, 16),
30960 => conv_std_logic_vector(28800, 16),
30961 => conv_std_logic_vector(28920, 16),
30962 => conv_std_logic_vector(29040, 16),
30963 => conv_std_logic_vector(29160, 16),
30964 => conv_std_logic_vector(29280, 16),
30965 => conv_std_logic_vector(29400, 16),
30966 => conv_std_logic_vector(29520, 16),
30967 => conv_std_logic_vector(29640, 16),
30968 => conv_std_logic_vector(29760, 16),
30969 => conv_std_logic_vector(29880, 16),
30970 => conv_std_logic_vector(30000, 16),
30971 => conv_std_logic_vector(30120, 16),
30972 => conv_std_logic_vector(30240, 16),
30973 => conv_std_logic_vector(30360, 16),
30974 => conv_std_logic_vector(30480, 16),
30975 => conv_std_logic_vector(30600, 16),
30976 => conv_std_logic_vector(0, 16),
30977 => conv_std_logic_vector(121, 16),
30978 => conv_std_logic_vector(242, 16),
30979 => conv_std_logic_vector(363, 16),
30980 => conv_std_logic_vector(484, 16),
30981 => conv_std_logic_vector(605, 16),
30982 => conv_std_logic_vector(726, 16),
30983 => conv_std_logic_vector(847, 16),
30984 => conv_std_logic_vector(968, 16),
30985 => conv_std_logic_vector(1089, 16),
30986 => conv_std_logic_vector(1210, 16),
30987 => conv_std_logic_vector(1331, 16),
30988 => conv_std_logic_vector(1452, 16),
30989 => conv_std_logic_vector(1573, 16),
30990 => conv_std_logic_vector(1694, 16),
30991 => conv_std_logic_vector(1815, 16),
30992 => conv_std_logic_vector(1936, 16),
30993 => conv_std_logic_vector(2057, 16),
30994 => conv_std_logic_vector(2178, 16),
30995 => conv_std_logic_vector(2299, 16),
30996 => conv_std_logic_vector(2420, 16),
30997 => conv_std_logic_vector(2541, 16),
30998 => conv_std_logic_vector(2662, 16),
30999 => conv_std_logic_vector(2783, 16),
31000 => conv_std_logic_vector(2904, 16),
31001 => conv_std_logic_vector(3025, 16),
31002 => conv_std_logic_vector(3146, 16),
31003 => conv_std_logic_vector(3267, 16),
31004 => conv_std_logic_vector(3388, 16),
31005 => conv_std_logic_vector(3509, 16),
31006 => conv_std_logic_vector(3630, 16),
31007 => conv_std_logic_vector(3751, 16),
31008 => conv_std_logic_vector(3872, 16),
31009 => conv_std_logic_vector(3993, 16),
31010 => conv_std_logic_vector(4114, 16),
31011 => conv_std_logic_vector(4235, 16),
31012 => conv_std_logic_vector(4356, 16),
31013 => conv_std_logic_vector(4477, 16),
31014 => conv_std_logic_vector(4598, 16),
31015 => conv_std_logic_vector(4719, 16),
31016 => conv_std_logic_vector(4840, 16),
31017 => conv_std_logic_vector(4961, 16),
31018 => conv_std_logic_vector(5082, 16),
31019 => conv_std_logic_vector(5203, 16),
31020 => conv_std_logic_vector(5324, 16),
31021 => conv_std_logic_vector(5445, 16),
31022 => conv_std_logic_vector(5566, 16),
31023 => conv_std_logic_vector(5687, 16),
31024 => conv_std_logic_vector(5808, 16),
31025 => conv_std_logic_vector(5929, 16),
31026 => conv_std_logic_vector(6050, 16),
31027 => conv_std_logic_vector(6171, 16),
31028 => conv_std_logic_vector(6292, 16),
31029 => conv_std_logic_vector(6413, 16),
31030 => conv_std_logic_vector(6534, 16),
31031 => conv_std_logic_vector(6655, 16),
31032 => conv_std_logic_vector(6776, 16),
31033 => conv_std_logic_vector(6897, 16),
31034 => conv_std_logic_vector(7018, 16),
31035 => conv_std_logic_vector(7139, 16),
31036 => conv_std_logic_vector(7260, 16),
31037 => conv_std_logic_vector(7381, 16),
31038 => conv_std_logic_vector(7502, 16),
31039 => conv_std_logic_vector(7623, 16),
31040 => conv_std_logic_vector(7744, 16),
31041 => conv_std_logic_vector(7865, 16),
31042 => conv_std_logic_vector(7986, 16),
31043 => conv_std_logic_vector(8107, 16),
31044 => conv_std_logic_vector(8228, 16),
31045 => conv_std_logic_vector(8349, 16),
31046 => conv_std_logic_vector(8470, 16),
31047 => conv_std_logic_vector(8591, 16),
31048 => conv_std_logic_vector(8712, 16),
31049 => conv_std_logic_vector(8833, 16),
31050 => conv_std_logic_vector(8954, 16),
31051 => conv_std_logic_vector(9075, 16),
31052 => conv_std_logic_vector(9196, 16),
31053 => conv_std_logic_vector(9317, 16),
31054 => conv_std_logic_vector(9438, 16),
31055 => conv_std_logic_vector(9559, 16),
31056 => conv_std_logic_vector(9680, 16),
31057 => conv_std_logic_vector(9801, 16),
31058 => conv_std_logic_vector(9922, 16),
31059 => conv_std_logic_vector(10043, 16),
31060 => conv_std_logic_vector(10164, 16),
31061 => conv_std_logic_vector(10285, 16),
31062 => conv_std_logic_vector(10406, 16),
31063 => conv_std_logic_vector(10527, 16),
31064 => conv_std_logic_vector(10648, 16),
31065 => conv_std_logic_vector(10769, 16),
31066 => conv_std_logic_vector(10890, 16),
31067 => conv_std_logic_vector(11011, 16),
31068 => conv_std_logic_vector(11132, 16),
31069 => conv_std_logic_vector(11253, 16),
31070 => conv_std_logic_vector(11374, 16),
31071 => conv_std_logic_vector(11495, 16),
31072 => conv_std_logic_vector(11616, 16),
31073 => conv_std_logic_vector(11737, 16),
31074 => conv_std_logic_vector(11858, 16),
31075 => conv_std_logic_vector(11979, 16),
31076 => conv_std_logic_vector(12100, 16),
31077 => conv_std_logic_vector(12221, 16),
31078 => conv_std_logic_vector(12342, 16),
31079 => conv_std_logic_vector(12463, 16),
31080 => conv_std_logic_vector(12584, 16),
31081 => conv_std_logic_vector(12705, 16),
31082 => conv_std_logic_vector(12826, 16),
31083 => conv_std_logic_vector(12947, 16),
31084 => conv_std_logic_vector(13068, 16),
31085 => conv_std_logic_vector(13189, 16),
31086 => conv_std_logic_vector(13310, 16),
31087 => conv_std_logic_vector(13431, 16),
31088 => conv_std_logic_vector(13552, 16),
31089 => conv_std_logic_vector(13673, 16),
31090 => conv_std_logic_vector(13794, 16),
31091 => conv_std_logic_vector(13915, 16),
31092 => conv_std_logic_vector(14036, 16),
31093 => conv_std_logic_vector(14157, 16),
31094 => conv_std_logic_vector(14278, 16),
31095 => conv_std_logic_vector(14399, 16),
31096 => conv_std_logic_vector(14520, 16),
31097 => conv_std_logic_vector(14641, 16),
31098 => conv_std_logic_vector(14762, 16),
31099 => conv_std_logic_vector(14883, 16),
31100 => conv_std_logic_vector(15004, 16),
31101 => conv_std_logic_vector(15125, 16),
31102 => conv_std_logic_vector(15246, 16),
31103 => conv_std_logic_vector(15367, 16),
31104 => conv_std_logic_vector(15488, 16),
31105 => conv_std_logic_vector(15609, 16),
31106 => conv_std_logic_vector(15730, 16),
31107 => conv_std_logic_vector(15851, 16),
31108 => conv_std_logic_vector(15972, 16),
31109 => conv_std_logic_vector(16093, 16),
31110 => conv_std_logic_vector(16214, 16),
31111 => conv_std_logic_vector(16335, 16),
31112 => conv_std_logic_vector(16456, 16),
31113 => conv_std_logic_vector(16577, 16),
31114 => conv_std_logic_vector(16698, 16),
31115 => conv_std_logic_vector(16819, 16),
31116 => conv_std_logic_vector(16940, 16),
31117 => conv_std_logic_vector(17061, 16),
31118 => conv_std_logic_vector(17182, 16),
31119 => conv_std_logic_vector(17303, 16),
31120 => conv_std_logic_vector(17424, 16),
31121 => conv_std_logic_vector(17545, 16),
31122 => conv_std_logic_vector(17666, 16),
31123 => conv_std_logic_vector(17787, 16),
31124 => conv_std_logic_vector(17908, 16),
31125 => conv_std_logic_vector(18029, 16),
31126 => conv_std_logic_vector(18150, 16),
31127 => conv_std_logic_vector(18271, 16),
31128 => conv_std_logic_vector(18392, 16),
31129 => conv_std_logic_vector(18513, 16),
31130 => conv_std_logic_vector(18634, 16),
31131 => conv_std_logic_vector(18755, 16),
31132 => conv_std_logic_vector(18876, 16),
31133 => conv_std_logic_vector(18997, 16),
31134 => conv_std_logic_vector(19118, 16),
31135 => conv_std_logic_vector(19239, 16),
31136 => conv_std_logic_vector(19360, 16),
31137 => conv_std_logic_vector(19481, 16),
31138 => conv_std_logic_vector(19602, 16),
31139 => conv_std_logic_vector(19723, 16),
31140 => conv_std_logic_vector(19844, 16),
31141 => conv_std_logic_vector(19965, 16),
31142 => conv_std_logic_vector(20086, 16),
31143 => conv_std_logic_vector(20207, 16),
31144 => conv_std_logic_vector(20328, 16),
31145 => conv_std_logic_vector(20449, 16),
31146 => conv_std_logic_vector(20570, 16),
31147 => conv_std_logic_vector(20691, 16),
31148 => conv_std_logic_vector(20812, 16),
31149 => conv_std_logic_vector(20933, 16),
31150 => conv_std_logic_vector(21054, 16),
31151 => conv_std_logic_vector(21175, 16),
31152 => conv_std_logic_vector(21296, 16),
31153 => conv_std_logic_vector(21417, 16),
31154 => conv_std_logic_vector(21538, 16),
31155 => conv_std_logic_vector(21659, 16),
31156 => conv_std_logic_vector(21780, 16),
31157 => conv_std_logic_vector(21901, 16),
31158 => conv_std_logic_vector(22022, 16),
31159 => conv_std_logic_vector(22143, 16),
31160 => conv_std_logic_vector(22264, 16),
31161 => conv_std_logic_vector(22385, 16),
31162 => conv_std_logic_vector(22506, 16),
31163 => conv_std_logic_vector(22627, 16),
31164 => conv_std_logic_vector(22748, 16),
31165 => conv_std_logic_vector(22869, 16),
31166 => conv_std_logic_vector(22990, 16),
31167 => conv_std_logic_vector(23111, 16),
31168 => conv_std_logic_vector(23232, 16),
31169 => conv_std_logic_vector(23353, 16),
31170 => conv_std_logic_vector(23474, 16),
31171 => conv_std_logic_vector(23595, 16),
31172 => conv_std_logic_vector(23716, 16),
31173 => conv_std_logic_vector(23837, 16),
31174 => conv_std_logic_vector(23958, 16),
31175 => conv_std_logic_vector(24079, 16),
31176 => conv_std_logic_vector(24200, 16),
31177 => conv_std_logic_vector(24321, 16),
31178 => conv_std_logic_vector(24442, 16),
31179 => conv_std_logic_vector(24563, 16),
31180 => conv_std_logic_vector(24684, 16),
31181 => conv_std_logic_vector(24805, 16),
31182 => conv_std_logic_vector(24926, 16),
31183 => conv_std_logic_vector(25047, 16),
31184 => conv_std_logic_vector(25168, 16),
31185 => conv_std_logic_vector(25289, 16),
31186 => conv_std_logic_vector(25410, 16),
31187 => conv_std_logic_vector(25531, 16),
31188 => conv_std_logic_vector(25652, 16),
31189 => conv_std_logic_vector(25773, 16),
31190 => conv_std_logic_vector(25894, 16),
31191 => conv_std_logic_vector(26015, 16),
31192 => conv_std_logic_vector(26136, 16),
31193 => conv_std_logic_vector(26257, 16),
31194 => conv_std_logic_vector(26378, 16),
31195 => conv_std_logic_vector(26499, 16),
31196 => conv_std_logic_vector(26620, 16),
31197 => conv_std_logic_vector(26741, 16),
31198 => conv_std_logic_vector(26862, 16),
31199 => conv_std_logic_vector(26983, 16),
31200 => conv_std_logic_vector(27104, 16),
31201 => conv_std_logic_vector(27225, 16),
31202 => conv_std_logic_vector(27346, 16),
31203 => conv_std_logic_vector(27467, 16),
31204 => conv_std_logic_vector(27588, 16),
31205 => conv_std_logic_vector(27709, 16),
31206 => conv_std_logic_vector(27830, 16),
31207 => conv_std_logic_vector(27951, 16),
31208 => conv_std_logic_vector(28072, 16),
31209 => conv_std_logic_vector(28193, 16),
31210 => conv_std_logic_vector(28314, 16),
31211 => conv_std_logic_vector(28435, 16),
31212 => conv_std_logic_vector(28556, 16),
31213 => conv_std_logic_vector(28677, 16),
31214 => conv_std_logic_vector(28798, 16),
31215 => conv_std_logic_vector(28919, 16),
31216 => conv_std_logic_vector(29040, 16),
31217 => conv_std_logic_vector(29161, 16),
31218 => conv_std_logic_vector(29282, 16),
31219 => conv_std_logic_vector(29403, 16),
31220 => conv_std_logic_vector(29524, 16),
31221 => conv_std_logic_vector(29645, 16),
31222 => conv_std_logic_vector(29766, 16),
31223 => conv_std_logic_vector(29887, 16),
31224 => conv_std_logic_vector(30008, 16),
31225 => conv_std_logic_vector(30129, 16),
31226 => conv_std_logic_vector(30250, 16),
31227 => conv_std_logic_vector(30371, 16),
31228 => conv_std_logic_vector(30492, 16),
31229 => conv_std_logic_vector(30613, 16),
31230 => conv_std_logic_vector(30734, 16),
31231 => conv_std_logic_vector(30855, 16),
31232 => conv_std_logic_vector(0, 16),
31233 => conv_std_logic_vector(122, 16),
31234 => conv_std_logic_vector(244, 16),
31235 => conv_std_logic_vector(366, 16),
31236 => conv_std_logic_vector(488, 16),
31237 => conv_std_logic_vector(610, 16),
31238 => conv_std_logic_vector(732, 16),
31239 => conv_std_logic_vector(854, 16),
31240 => conv_std_logic_vector(976, 16),
31241 => conv_std_logic_vector(1098, 16),
31242 => conv_std_logic_vector(1220, 16),
31243 => conv_std_logic_vector(1342, 16),
31244 => conv_std_logic_vector(1464, 16),
31245 => conv_std_logic_vector(1586, 16),
31246 => conv_std_logic_vector(1708, 16),
31247 => conv_std_logic_vector(1830, 16),
31248 => conv_std_logic_vector(1952, 16),
31249 => conv_std_logic_vector(2074, 16),
31250 => conv_std_logic_vector(2196, 16),
31251 => conv_std_logic_vector(2318, 16),
31252 => conv_std_logic_vector(2440, 16),
31253 => conv_std_logic_vector(2562, 16),
31254 => conv_std_logic_vector(2684, 16),
31255 => conv_std_logic_vector(2806, 16),
31256 => conv_std_logic_vector(2928, 16),
31257 => conv_std_logic_vector(3050, 16),
31258 => conv_std_logic_vector(3172, 16),
31259 => conv_std_logic_vector(3294, 16),
31260 => conv_std_logic_vector(3416, 16),
31261 => conv_std_logic_vector(3538, 16),
31262 => conv_std_logic_vector(3660, 16),
31263 => conv_std_logic_vector(3782, 16),
31264 => conv_std_logic_vector(3904, 16),
31265 => conv_std_logic_vector(4026, 16),
31266 => conv_std_logic_vector(4148, 16),
31267 => conv_std_logic_vector(4270, 16),
31268 => conv_std_logic_vector(4392, 16),
31269 => conv_std_logic_vector(4514, 16),
31270 => conv_std_logic_vector(4636, 16),
31271 => conv_std_logic_vector(4758, 16),
31272 => conv_std_logic_vector(4880, 16),
31273 => conv_std_logic_vector(5002, 16),
31274 => conv_std_logic_vector(5124, 16),
31275 => conv_std_logic_vector(5246, 16),
31276 => conv_std_logic_vector(5368, 16),
31277 => conv_std_logic_vector(5490, 16),
31278 => conv_std_logic_vector(5612, 16),
31279 => conv_std_logic_vector(5734, 16),
31280 => conv_std_logic_vector(5856, 16),
31281 => conv_std_logic_vector(5978, 16),
31282 => conv_std_logic_vector(6100, 16),
31283 => conv_std_logic_vector(6222, 16),
31284 => conv_std_logic_vector(6344, 16),
31285 => conv_std_logic_vector(6466, 16),
31286 => conv_std_logic_vector(6588, 16),
31287 => conv_std_logic_vector(6710, 16),
31288 => conv_std_logic_vector(6832, 16),
31289 => conv_std_logic_vector(6954, 16),
31290 => conv_std_logic_vector(7076, 16),
31291 => conv_std_logic_vector(7198, 16),
31292 => conv_std_logic_vector(7320, 16),
31293 => conv_std_logic_vector(7442, 16),
31294 => conv_std_logic_vector(7564, 16),
31295 => conv_std_logic_vector(7686, 16),
31296 => conv_std_logic_vector(7808, 16),
31297 => conv_std_logic_vector(7930, 16),
31298 => conv_std_logic_vector(8052, 16),
31299 => conv_std_logic_vector(8174, 16),
31300 => conv_std_logic_vector(8296, 16),
31301 => conv_std_logic_vector(8418, 16),
31302 => conv_std_logic_vector(8540, 16),
31303 => conv_std_logic_vector(8662, 16),
31304 => conv_std_logic_vector(8784, 16),
31305 => conv_std_logic_vector(8906, 16),
31306 => conv_std_logic_vector(9028, 16),
31307 => conv_std_logic_vector(9150, 16),
31308 => conv_std_logic_vector(9272, 16),
31309 => conv_std_logic_vector(9394, 16),
31310 => conv_std_logic_vector(9516, 16),
31311 => conv_std_logic_vector(9638, 16),
31312 => conv_std_logic_vector(9760, 16),
31313 => conv_std_logic_vector(9882, 16),
31314 => conv_std_logic_vector(10004, 16),
31315 => conv_std_logic_vector(10126, 16),
31316 => conv_std_logic_vector(10248, 16),
31317 => conv_std_logic_vector(10370, 16),
31318 => conv_std_logic_vector(10492, 16),
31319 => conv_std_logic_vector(10614, 16),
31320 => conv_std_logic_vector(10736, 16),
31321 => conv_std_logic_vector(10858, 16),
31322 => conv_std_logic_vector(10980, 16),
31323 => conv_std_logic_vector(11102, 16),
31324 => conv_std_logic_vector(11224, 16),
31325 => conv_std_logic_vector(11346, 16),
31326 => conv_std_logic_vector(11468, 16),
31327 => conv_std_logic_vector(11590, 16),
31328 => conv_std_logic_vector(11712, 16),
31329 => conv_std_logic_vector(11834, 16),
31330 => conv_std_logic_vector(11956, 16),
31331 => conv_std_logic_vector(12078, 16),
31332 => conv_std_logic_vector(12200, 16),
31333 => conv_std_logic_vector(12322, 16),
31334 => conv_std_logic_vector(12444, 16),
31335 => conv_std_logic_vector(12566, 16),
31336 => conv_std_logic_vector(12688, 16),
31337 => conv_std_logic_vector(12810, 16),
31338 => conv_std_logic_vector(12932, 16),
31339 => conv_std_logic_vector(13054, 16),
31340 => conv_std_logic_vector(13176, 16),
31341 => conv_std_logic_vector(13298, 16),
31342 => conv_std_logic_vector(13420, 16),
31343 => conv_std_logic_vector(13542, 16),
31344 => conv_std_logic_vector(13664, 16),
31345 => conv_std_logic_vector(13786, 16),
31346 => conv_std_logic_vector(13908, 16),
31347 => conv_std_logic_vector(14030, 16),
31348 => conv_std_logic_vector(14152, 16),
31349 => conv_std_logic_vector(14274, 16),
31350 => conv_std_logic_vector(14396, 16),
31351 => conv_std_logic_vector(14518, 16),
31352 => conv_std_logic_vector(14640, 16),
31353 => conv_std_logic_vector(14762, 16),
31354 => conv_std_logic_vector(14884, 16),
31355 => conv_std_logic_vector(15006, 16),
31356 => conv_std_logic_vector(15128, 16),
31357 => conv_std_logic_vector(15250, 16),
31358 => conv_std_logic_vector(15372, 16),
31359 => conv_std_logic_vector(15494, 16),
31360 => conv_std_logic_vector(15616, 16),
31361 => conv_std_logic_vector(15738, 16),
31362 => conv_std_logic_vector(15860, 16),
31363 => conv_std_logic_vector(15982, 16),
31364 => conv_std_logic_vector(16104, 16),
31365 => conv_std_logic_vector(16226, 16),
31366 => conv_std_logic_vector(16348, 16),
31367 => conv_std_logic_vector(16470, 16),
31368 => conv_std_logic_vector(16592, 16),
31369 => conv_std_logic_vector(16714, 16),
31370 => conv_std_logic_vector(16836, 16),
31371 => conv_std_logic_vector(16958, 16),
31372 => conv_std_logic_vector(17080, 16),
31373 => conv_std_logic_vector(17202, 16),
31374 => conv_std_logic_vector(17324, 16),
31375 => conv_std_logic_vector(17446, 16),
31376 => conv_std_logic_vector(17568, 16),
31377 => conv_std_logic_vector(17690, 16),
31378 => conv_std_logic_vector(17812, 16),
31379 => conv_std_logic_vector(17934, 16),
31380 => conv_std_logic_vector(18056, 16),
31381 => conv_std_logic_vector(18178, 16),
31382 => conv_std_logic_vector(18300, 16),
31383 => conv_std_logic_vector(18422, 16),
31384 => conv_std_logic_vector(18544, 16),
31385 => conv_std_logic_vector(18666, 16),
31386 => conv_std_logic_vector(18788, 16),
31387 => conv_std_logic_vector(18910, 16),
31388 => conv_std_logic_vector(19032, 16),
31389 => conv_std_logic_vector(19154, 16),
31390 => conv_std_logic_vector(19276, 16),
31391 => conv_std_logic_vector(19398, 16),
31392 => conv_std_logic_vector(19520, 16),
31393 => conv_std_logic_vector(19642, 16),
31394 => conv_std_logic_vector(19764, 16),
31395 => conv_std_logic_vector(19886, 16),
31396 => conv_std_logic_vector(20008, 16),
31397 => conv_std_logic_vector(20130, 16),
31398 => conv_std_logic_vector(20252, 16),
31399 => conv_std_logic_vector(20374, 16),
31400 => conv_std_logic_vector(20496, 16),
31401 => conv_std_logic_vector(20618, 16),
31402 => conv_std_logic_vector(20740, 16),
31403 => conv_std_logic_vector(20862, 16),
31404 => conv_std_logic_vector(20984, 16),
31405 => conv_std_logic_vector(21106, 16),
31406 => conv_std_logic_vector(21228, 16),
31407 => conv_std_logic_vector(21350, 16),
31408 => conv_std_logic_vector(21472, 16),
31409 => conv_std_logic_vector(21594, 16),
31410 => conv_std_logic_vector(21716, 16),
31411 => conv_std_logic_vector(21838, 16),
31412 => conv_std_logic_vector(21960, 16),
31413 => conv_std_logic_vector(22082, 16),
31414 => conv_std_logic_vector(22204, 16),
31415 => conv_std_logic_vector(22326, 16),
31416 => conv_std_logic_vector(22448, 16),
31417 => conv_std_logic_vector(22570, 16),
31418 => conv_std_logic_vector(22692, 16),
31419 => conv_std_logic_vector(22814, 16),
31420 => conv_std_logic_vector(22936, 16),
31421 => conv_std_logic_vector(23058, 16),
31422 => conv_std_logic_vector(23180, 16),
31423 => conv_std_logic_vector(23302, 16),
31424 => conv_std_logic_vector(23424, 16),
31425 => conv_std_logic_vector(23546, 16),
31426 => conv_std_logic_vector(23668, 16),
31427 => conv_std_logic_vector(23790, 16),
31428 => conv_std_logic_vector(23912, 16),
31429 => conv_std_logic_vector(24034, 16),
31430 => conv_std_logic_vector(24156, 16),
31431 => conv_std_logic_vector(24278, 16),
31432 => conv_std_logic_vector(24400, 16),
31433 => conv_std_logic_vector(24522, 16),
31434 => conv_std_logic_vector(24644, 16),
31435 => conv_std_logic_vector(24766, 16),
31436 => conv_std_logic_vector(24888, 16),
31437 => conv_std_logic_vector(25010, 16),
31438 => conv_std_logic_vector(25132, 16),
31439 => conv_std_logic_vector(25254, 16),
31440 => conv_std_logic_vector(25376, 16),
31441 => conv_std_logic_vector(25498, 16),
31442 => conv_std_logic_vector(25620, 16),
31443 => conv_std_logic_vector(25742, 16),
31444 => conv_std_logic_vector(25864, 16),
31445 => conv_std_logic_vector(25986, 16),
31446 => conv_std_logic_vector(26108, 16),
31447 => conv_std_logic_vector(26230, 16),
31448 => conv_std_logic_vector(26352, 16),
31449 => conv_std_logic_vector(26474, 16),
31450 => conv_std_logic_vector(26596, 16),
31451 => conv_std_logic_vector(26718, 16),
31452 => conv_std_logic_vector(26840, 16),
31453 => conv_std_logic_vector(26962, 16),
31454 => conv_std_logic_vector(27084, 16),
31455 => conv_std_logic_vector(27206, 16),
31456 => conv_std_logic_vector(27328, 16),
31457 => conv_std_logic_vector(27450, 16),
31458 => conv_std_logic_vector(27572, 16),
31459 => conv_std_logic_vector(27694, 16),
31460 => conv_std_logic_vector(27816, 16),
31461 => conv_std_logic_vector(27938, 16),
31462 => conv_std_logic_vector(28060, 16),
31463 => conv_std_logic_vector(28182, 16),
31464 => conv_std_logic_vector(28304, 16),
31465 => conv_std_logic_vector(28426, 16),
31466 => conv_std_logic_vector(28548, 16),
31467 => conv_std_logic_vector(28670, 16),
31468 => conv_std_logic_vector(28792, 16),
31469 => conv_std_logic_vector(28914, 16),
31470 => conv_std_logic_vector(29036, 16),
31471 => conv_std_logic_vector(29158, 16),
31472 => conv_std_logic_vector(29280, 16),
31473 => conv_std_logic_vector(29402, 16),
31474 => conv_std_logic_vector(29524, 16),
31475 => conv_std_logic_vector(29646, 16),
31476 => conv_std_logic_vector(29768, 16),
31477 => conv_std_logic_vector(29890, 16),
31478 => conv_std_logic_vector(30012, 16),
31479 => conv_std_logic_vector(30134, 16),
31480 => conv_std_logic_vector(30256, 16),
31481 => conv_std_logic_vector(30378, 16),
31482 => conv_std_logic_vector(30500, 16),
31483 => conv_std_logic_vector(30622, 16),
31484 => conv_std_logic_vector(30744, 16),
31485 => conv_std_logic_vector(30866, 16),
31486 => conv_std_logic_vector(30988, 16),
31487 => conv_std_logic_vector(31110, 16),
31488 => conv_std_logic_vector(0, 16),
31489 => conv_std_logic_vector(123, 16),
31490 => conv_std_logic_vector(246, 16),
31491 => conv_std_logic_vector(369, 16),
31492 => conv_std_logic_vector(492, 16),
31493 => conv_std_logic_vector(615, 16),
31494 => conv_std_logic_vector(738, 16),
31495 => conv_std_logic_vector(861, 16),
31496 => conv_std_logic_vector(984, 16),
31497 => conv_std_logic_vector(1107, 16),
31498 => conv_std_logic_vector(1230, 16),
31499 => conv_std_logic_vector(1353, 16),
31500 => conv_std_logic_vector(1476, 16),
31501 => conv_std_logic_vector(1599, 16),
31502 => conv_std_logic_vector(1722, 16),
31503 => conv_std_logic_vector(1845, 16),
31504 => conv_std_logic_vector(1968, 16),
31505 => conv_std_logic_vector(2091, 16),
31506 => conv_std_logic_vector(2214, 16),
31507 => conv_std_logic_vector(2337, 16),
31508 => conv_std_logic_vector(2460, 16),
31509 => conv_std_logic_vector(2583, 16),
31510 => conv_std_logic_vector(2706, 16),
31511 => conv_std_logic_vector(2829, 16),
31512 => conv_std_logic_vector(2952, 16),
31513 => conv_std_logic_vector(3075, 16),
31514 => conv_std_logic_vector(3198, 16),
31515 => conv_std_logic_vector(3321, 16),
31516 => conv_std_logic_vector(3444, 16),
31517 => conv_std_logic_vector(3567, 16),
31518 => conv_std_logic_vector(3690, 16),
31519 => conv_std_logic_vector(3813, 16),
31520 => conv_std_logic_vector(3936, 16),
31521 => conv_std_logic_vector(4059, 16),
31522 => conv_std_logic_vector(4182, 16),
31523 => conv_std_logic_vector(4305, 16),
31524 => conv_std_logic_vector(4428, 16),
31525 => conv_std_logic_vector(4551, 16),
31526 => conv_std_logic_vector(4674, 16),
31527 => conv_std_logic_vector(4797, 16),
31528 => conv_std_logic_vector(4920, 16),
31529 => conv_std_logic_vector(5043, 16),
31530 => conv_std_logic_vector(5166, 16),
31531 => conv_std_logic_vector(5289, 16),
31532 => conv_std_logic_vector(5412, 16),
31533 => conv_std_logic_vector(5535, 16),
31534 => conv_std_logic_vector(5658, 16),
31535 => conv_std_logic_vector(5781, 16),
31536 => conv_std_logic_vector(5904, 16),
31537 => conv_std_logic_vector(6027, 16),
31538 => conv_std_logic_vector(6150, 16),
31539 => conv_std_logic_vector(6273, 16),
31540 => conv_std_logic_vector(6396, 16),
31541 => conv_std_logic_vector(6519, 16),
31542 => conv_std_logic_vector(6642, 16),
31543 => conv_std_logic_vector(6765, 16),
31544 => conv_std_logic_vector(6888, 16),
31545 => conv_std_logic_vector(7011, 16),
31546 => conv_std_logic_vector(7134, 16),
31547 => conv_std_logic_vector(7257, 16),
31548 => conv_std_logic_vector(7380, 16),
31549 => conv_std_logic_vector(7503, 16),
31550 => conv_std_logic_vector(7626, 16),
31551 => conv_std_logic_vector(7749, 16),
31552 => conv_std_logic_vector(7872, 16),
31553 => conv_std_logic_vector(7995, 16),
31554 => conv_std_logic_vector(8118, 16),
31555 => conv_std_logic_vector(8241, 16),
31556 => conv_std_logic_vector(8364, 16),
31557 => conv_std_logic_vector(8487, 16),
31558 => conv_std_logic_vector(8610, 16),
31559 => conv_std_logic_vector(8733, 16),
31560 => conv_std_logic_vector(8856, 16),
31561 => conv_std_logic_vector(8979, 16),
31562 => conv_std_logic_vector(9102, 16),
31563 => conv_std_logic_vector(9225, 16),
31564 => conv_std_logic_vector(9348, 16),
31565 => conv_std_logic_vector(9471, 16),
31566 => conv_std_logic_vector(9594, 16),
31567 => conv_std_logic_vector(9717, 16),
31568 => conv_std_logic_vector(9840, 16),
31569 => conv_std_logic_vector(9963, 16),
31570 => conv_std_logic_vector(10086, 16),
31571 => conv_std_logic_vector(10209, 16),
31572 => conv_std_logic_vector(10332, 16),
31573 => conv_std_logic_vector(10455, 16),
31574 => conv_std_logic_vector(10578, 16),
31575 => conv_std_logic_vector(10701, 16),
31576 => conv_std_logic_vector(10824, 16),
31577 => conv_std_logic_vector(10947, 16),
31578 => conv_std_logic_vector(11070, 16),
31579 => conv_std_logic_vector(11193, 16),
31580 => conv_std_logic_vector(11316, 16),
31581 => conv_std_logic_vector(11439, 16),
31582 => conv_std_logic_vector(11562, 16),
31583 => conv_std_logic_vector(11685, 16),
31584 => conv_std_logic_vector(11808, 16),
31585 => conv_std_logic_vector(11931, 16),
31586 => conv_std_logic_vector(12054, 16),
31587 => conv_std_logic_vector(12177, 16),
31588 => conv_std_logic_vector(12300, 16),
31589 => conv_std_logic_vector(12423, 16),
31590 => conv_std_logic_vector(12546, 16),
31591 => conv_std_logic_vector(12669, 16),
31592 => conv_std_logic_vector(12792, 16),
31593 => conv_std_logic_vector(12915, 16),
31594 => conv_std_logic_vector(13038, 16),
31595 => conv_std_logic_vector(13161, 16),
31596 => conv_std_logic_vector(13284, 16),
31597 => conv_std_logic_vector(13407, 16),
31598 => conv_std_logic_vector(13530, 16),
31599 => conv_std_logic_vector(13653, 16),
31600 => conv_std_logic_vector(13776, 16),
31601 => conv_std_logic_vector(13899, 16),
31602 => conv_std_logic_vector(14022, 16),
31603 => conv_std_logic_vector(14145, 16),
31604 => conv_std_logic_vector(14268, 16),
31605 => conv_std_logic_vector(14391, 16),
31606 => conv_std_logic_vector(14514, 16),
31607 => conv_std_logic_vector(14637, 16),
31608 => conv_std_logic_vector(14760, 16),
31609 => conv_std_logic_vector(14883, 16),
31610 => conv_std_logic_vector(15006, 16),
31611 => conv_std_logic_vector(15129, 16),
31612 => conv_std_logic_vector(15252, 16),
31613 => conv_std_logic_vector(15375, 16),
31614 => conv_std_logic_vector(15498, 16),
31615 => conv_std_logic_vector(15621, 16),
31616 => conv_std_logic_vector(15744, 16),
31617 => conv_std_logic_vector(15867, 16),
31618 => conv_std_logic_vector(15990, 16),
31619 => conv_std_logic_vector(16113, 16),
31620 => conv_std_logic_vector(16236, 16),
31621 => conv_std_logic_vector(16359, 16),
31622 => conv_std_logic_vector(16482, 16),
31623 => conv_std_logic_vector(16605, 16),
31624 => conv_std_logic_vector(16728, 16),
31625 => conv_std_logic_vector(16851, 16),
31626 => conv_std_logic_vector(16974, 16),
31627 => conv_std_logic_vector(17097, 16),
31628 => conv_std_logic_vector(17220, 16),
31629 => conv_std_logic_vector(17343, 16),
31630 => conv_std_logic_vector(17466, 16),
31631 => conv_std_logic_vector(17589, 16),
31632 => conv_std_logic_vector(17712, 16),
31633 => conv_std_logic_vector(17835, 16),
31634 => conv_std_logic_vector(17958, 16),
31635 => conv_std_logic_vector(18081, 16),
31636 => conv_std_logic_vector(18204, 16),
31637 => conv_std_logic_vector(18327, 16),
31638 => conv_std_logic_vector(18450, 16),
31639 => conv_std_logic_vector(18573, 16),
31640 => conv_std_logic_vector(18696, 16),
31641 => conv_std_logic_vector(18819, 16),
31642 => conv_std_logic_vector(18942, 16),
31643 => conv_std_logic_vector(19065, 16),
31644 => conv_std_logic_vector(19188, 16),
31645 => conv_std_logic_vector(19311, 16),
31646 => conv_std_logic_vector(19434, 16),
31647 => conv_std_logic_vector(19557, 16),
31648 => conv_std_logic_vector(19680, 16),
31649 => conv_std_logic_vector(19803, 16),
31650 => conv_std_logic_vector(19926, 16),
31651 => conv_std_logic_vector(20049, 16),
31652 => conv_std_logic_vector(20172, 16),
31653 => conv_std_logic_vector(20295, 16),
31654 => conv_std_logic_vector(20418, 16),
31655 => conv_std_logic_vector(20541, 16),
31656 => conv_std_logic_vector(20664, 16),
31657 => conv_std_logic_vector(20787, 16),
31658 => conv_std_logic_vector(20910, 16),
31659 => conv_std_logic_vector(21033, 16),
31660 => conv_std_logic_vector(21156, 16),
31661 => conv_std_logic_vector(21279, 16),
31662 => conv_std_logic_vector(21402, 16),
31663 => conv_std_logic_vector(21525, 16),
31664 => conv_std_logic_vector(21648, 16),
31665 => conv_std_logic_vector(21771, 16),
31666 => conv_std_logic_vector(21894, 16),
31667 => conv_std_logic_vector(22017, 16),
31668 => conv_std_logic_vector(22140, 16),
31669 => conv_std_logic_vector(22263, 16),
31670 => conv_std_logic_vector(22386, 16),
31671 => conv_std_logic_vector(22509, 16),
31672 => conv_std_logic_vector(22632, 16),
31673 => conv_std_logic_vector(22755, 16),
31674 => conv_std_logic_vector(22878, 16),
31675 => conv_std_logic_vector(23001, 16),
31676 => conv_std_logic_vector(23124, 16),
31677 => conv_std_logic_vector(23247, 16),
31678 => conv_std_logic_vector(23370, 16),
31679 => conv_std_logic_vector(23493, 16),
31680 => conv_std_logic_vector(23616, 16),
31681 => conv_std_logic_vector(23739, 16),
31682 => conv_std_logic_vector(23862, 16),
31683 => conv_std_logic_vector(23985, 16),
31684 => conv_std_logic_vector(24108, 16),
31685 => conv_std_logic_vector(24231, 16),
31686 => conv_std_logic_vector(24354, 16),
31687 => conv_std_logic_vector(24477, 16),
31688 => conv_std_logic_vector(24600, 16),
31689 => conv_std_logic_vector(24723, 16),
31690 => conv_std_logic_vector(24846, 16),
31691 => conv_std_logic_vector(24969, 16),
31692 => conv_std_logic_vector(25092, 16),
31693 => conv_std_logic_vector(25215, 16),
31694 => conv_std_logic_vector(25338, 16),
31695 => conv_std_logic_vector(25461, 16),
31696 => conv_std_logic_vector(25584, 16),
31697 => conv_std_logic_vector(25707, 16),
31698 => conv_std_logic_vector(25830, 16),
31699 => conv_std_logic_vector(25953, 16),
31700 => conv_std_logic_vector(26076, 16),
31701 => conv_std_logic_vector(26199, 16),
31702 => conv_std_logic_vector(26322, 16),
31703 => conv_std_logic_vector(26445, 16),
31704 => conv_std_logic_vector(26568, 16),
31705 => conv_std_logic_vector(26691, 16),
31706 => conv_std_logic_vector(26814, 16),
31707 => conv_std_logic_vector(26937, 16),
31708 => conv_std_logic_vector(27060, 16),
31709 => conv_std_logic_vector(27183, 16),
31710 => conv_std_logic_vector(27306, 16),
31711 => conv_std_logic_vector(27429, 16),
31712 => conv_std_logic_vector(27552, 16),
31713 => conv_std_logic_vector(27675, 16),
31714 => conv_std_logic_vector(27798, 16),
31715 => conv_std_logic_vector(27921, 16),
31716 => conv_std_logic_vector(28044, 16),
31717 => conv_std_logic_vector(28167, 16),
31718 => conv_std_logic_vector(28290, 16),
31719 => conv_std_logic_vector(28413, 16),
31720 => conv_std_logic_vector(28536, 16),
31721 => conv_std_logic_vector(28659, 16),
31722 => conv_std_logic_vector(28782, 16),
31723 => conv_std_logic_vector(28905, 16),
31724 => conv_std_logic_vector(29028, 16),
31725 => conv_std_logic_vector(29151, 16),
31726 => conv_std_logic_vector(29274, 16),
31727 => conv_std_logic_vector(29397, 16),
31728 => conv_std_logic_vector(29520, 16),
31729 => conv_std_logic_vector(29643, 16),
31730 => conv_std_logic_vector(29766, 16),
31731 => conv_std_logic_vector(29889, 16),
31732 => conv_std_logic_vector(30012, 16),
31733 => conv_std_logic_vector(30135, 16),
31734 => conv_std_logic_vector(30258, 16),
31735 => conv_std_logic_vector(30381, 16),
31736 => conv_std_logic_vector(30504, 16),
31737 => conv_std_logic_vector(30627, 16),
31738 => conv_std_logic_vector(30750, 16),
31739 => conv_std_logic_vector(30873, 16),
31740 => conv_std_logic_vector(30996, 16),
31741 => conv_std_logic_vector(31119, 16),
31742 => conv_std_logic_vector(31242, 16),
31743 => conv_std_logic_vector(31365, 16),
31744 => conv_std_logic_vector(0, 16),
31745 => conv_std_logic_vector(124, 16),
31746 => conv_std_logic_vector(248, 16),
31747 => conv_std_logic_vector(372, 16),
31748 => conv_std_logic_vector(496, 16),
31749 => conv_std_logic_vector(620, 16),
31750 => conv_std_logic_vector(744, 16),
31751 => conv_std_logic_vector(868, 16),
31752 => conv_std_logic_vector(992, 16),
31753 => conv_std_logic_vector(1116, 16),
31754 => conv_std_logic_vector(1240, 16),
31755 => conv_std_logic_vector(1364, 16),
31756 => conv_std_logic_vector(1488, 16),
31757 => conv_std_logic_vector(1612, 16),
31758 => conv_std_logic_vector(1736, 16),
31759 => conv_std_logic_vector(1860, 16),
31760 => conv_std_logic_vector(1984, 16),
31761 => conv_std_logic_vector(2108, 16),
31762 => conv_std_logic_vector(2232, 16),
31763 => conv_std_logic_vector(2356, 16),
31764 => conv_std_logic_vector(2480, 16),
31765 => conv_std_logic_vector(2604, 16),
31766 => conv_std_logic_vector(2728, 16),
31767 => conv_std_logic_vector(2852, 16),
31768 => conv_std_logic_vector(2976, 16),
31769 => conv_std_logic_vector(3100, 16),
31770 => conv_std_logic_vector(3224, 16),
31771 => conv_std_logic_vector(3348, 16),
31772 => conv_std_logic_vector(3472, 16),
31773 => conv_std_logic_vector(3596, 16),
31774 => conv_std_logic_vector(3720, 16),
31775 => conv_std_logic_vector(3844, 16),
31776 => conv_std_logic_vector(3968, 16),
31777 => conv_std_logic_vector(4092, 16),
31778 => conv_std_logic_vector(4216, 16),
31779 => conv_std_logic_vector(4340, 16),
31780 => conv_std_logic_vector(4464, 16),
31781 => conv_std_logic_vector(4588, 16),
31782 => conv_std_logic_vector(4712, 16),
31783 => conv_std_logic_vector(4836, 16),
31784 => conv_std_logic_vector(4960, 16),
31785 => conv_std_logic_vector(5084, 16),
31786 => conv_std_logic_vector(5208, 16),
31787 => conv_std_logic_vector(5332, 16),
31788 => conv_std_logic_vector(5456, 16),
31789 => conv_std_logic_vector(5580, 16),
31790 => conv_std_logic_vector(5704, 16),
31791 => conv_std_logic_vector(5828, 16),
31792 => conv_std_logic_vector(5952, 16),
31793 => conv_std_logic_vector(6076, 16),
31794 => conv_std_logic_vector(6200, 16),
31795 => conv_std_logic_vector(6324, 16),
31796 => conv_std_logic_vector(6448, 16),
31797 => conv_std_logic_vector(6572, 16),
31798 => conv_std_logic_vector(6696, 16),
31799 => conv_std_logic_vector(6820, 16),
31800 => conv_std_logic_vector(6944, 16),
31801 => conv_std_logic_vector(7068, 16),
31802 => conv_std_logic_vector(7192, 16),
31803 => conv_std_logic_vector(7316, 16),
31804 => conv_std_logic_vector(7440, 16),
31805 => conv_std_logic_vector(7564, 16),
31806 => conv_std_logic_vector(7688, 16),
31807 => conv_std_logic_vector(7812, 16),
31808 => conv_std_logic_vector(7936, 16),
31809 => conv_std_logic_vector(8060, 16),
31810 => conv_std_logic_vector(8184, 16),
31811 => conv_std_logic_vector(8308, 16),
31812 => conv_std_logic_vector(8432, 16),
31813 => conv_std_logic_vector(8556, 16),
31814 => conv_std_logic_vector(8680, 16),
31815 => conv_std_logic_vector(8804, 16),
31816 => conv_std_logic_vector(8928, 16),
31817 => conv_std_logic_vector(9052, 16),
31818 => conv_std_logic_vector(9176, 16),
31819 => conv_std_logic_vector(9300, 16),
31820 => conv_std_logic_vector(9424, 16),
31821 => conv_std_logic_vector(9548, 16),
31822 => conv_std_logic_vector(9672, 16),
31823 => conv_std_logic_vector(9796, 16),
31824 => conv_std_logic_vector(9920, 16),
31825 => conv_std_logic_vector(10044, 16),
31826 => conv_std_logic_vector(10168, 16),
31827 => conv_std_logic_vector(10292, 16),
31828 => conv_std_logic_vector(10416, 16),
31829 => conv_std_logic_vector(10540, 16),
31830 => conv_std_logic_vector(10664, 16),
31831 => conv_std_logic_vector(10788, 16),
31832 => conv_std_logic_vector(10912, 16),
31833 => conv_std_logic_vector(11036, 16),
31834 => conv_std_logic_vector(11160, 16),
31835 => conv_std_logic_vector(11284, 16),
31836 => conv_std_logic_vector(11408, 16),
31837 => conv_std_logic_vector(11532, 16),
31838 => conv_std_logic_vector(11656, 16),
31839 => conv_std_logic_vector(11780, 16),
31840 => conv_std_logic_vector(11904, 16),
31841 => conv_std_logic_vector(12028, 16),
31842 => conv_std_logic_vector(12152, 16),
31843 => conv_std_logic_vector(12276, 16),
31844 => conv_std_logic_vector(12400, 16),
31845 => conv_std_logic_vector(12524, 16),
31846 => conv_std_logic_vector(12648, 16),
31847 => conv_std_logic_vector(12772, 16),
31848 => conv_std_logic_vector(12896, 16),
31849 => conv_std_logic_vector(13020, 16),
31850 => conv_std_logic_vector(13144, 16),
31851 => conv_std_logic_vector(13268, 16),
31852 => conv_std_logic_vector(13392, 16),
31853 => conv_std_logic_vector(13516, 16),
31854 => conv_std_logic_vector(13640, 16),
31855 => conv_std_logic_vector(13764, 16),
31856 => conv_std_logic_vector(13888, 16),
31857 => conv_std_logic_vector(14012, 16),
31858 => conv_std_logic_vector(14136, 16),
31859 => conv_std_logic_vector(14260, 16),
31860 => conv_std_logic_vector(14384, 16),
31861 => conv_std_logic_vector(14508, 16),
31862 => conv_std_logic_vector(14632, 16),
31863 => conv_std_logic_vector(14756, 16),
31864 => conv_std_logic_vector(14880, 16),
31865 => conv_std_logic_vector(15004, 16),
31866 => conv_std_logic_vector(15128, 16),
31867 => conv_std_logic_vector(15252, 16),
31868 => conv_std_logic_vector(15376, 16),
31869 => conv_std_logic_vector(15500, 16),
31870 => conv_std_logic_vector(15624, 16),
31871 => conv_std_logic_vector(15748, 16),
31872 => conv_std_logic_vector(15872, 16),
31873 => conv_std_logic_vector(15996, 16),
31874 => conv_std_logic_vector(16120, 16),
31875 => conv_std_logic_vector(16244, 16),
31876 => conv_std_logic_vector(16368, 16),
31877 => conv_std_logic_vector(16492, 16),
31878 => conv_std_logic_vector(16616, 16),
31879 => conv_std_logic_vector(16740, 16),
31880 => conv_std_logic_vector(16864, 16),
31881 => conv_std_logic_vector(16988, 16),
31882 => conv_std_logic_vector(17112, 16),
31883 => conv_std_logic_vector(17236, 16),
31884 => conv_std_logic_vector(17360, 16),
31885 => conv_std_logic_vector(17484, 16),
31886 => conv_std_logic_vector(17608, 16),
31887 => conv_std_logic_vector(17732, 16),
31888 => conv_std_logic_vector(17856, 16),
31889 => conv_std_logic_vector(17980, 16),
31890 => conv_std_logic_vector(18104, 16),
31891 => conv_std_logic_vector(18228, 16),
31892 => conv_std_logic_vector(18352, 16),
31893 => conv_std_logic_vector(18476, 16),
31894 => conv_std_logic_vector(18600, 16),
31895 => conv_std_logic_vector(18724, 16),
31896 => conv_std_logic_vector(18848, 16),
31897 => conv_std_logic_vector(18972, 16),
31898 => conv_std_logic_vector(19096, 16),
31899 => conv_std_logic_vector(19220, 16),
31900 => conv_std_logic_vector(19344, 16),
31901 => conv_std_logic_vector(19468, 16),
31902 => conv_std_logic_vector(19592, 16),
31903 => conv_std_logic_vector(19716, 16),
31904 => conv_std_logic_vector(19840, 16),
31905 => conv_std_logic_vector(19964, 16),
31906 => conv_std_logic_vector(20088, 16),
31907 => conv_std_logic_vector(20212, 16),
31908 => conv_std_logic_vector(20336, 16),
31909 => conv_std_logic_vector(20460, 16),
31910 => conv_std_logic_vector(20584, 16),
31911 => conv_std_logic_vector(20708, 16),
31912 => conv_std_logic_vector(20832, 16),
31913 => conv_std_logic_vector(20956, 16),
31914 => conv_std_logic_vector(21080, 16),
31915 => conv_std_logic_vector(21204, 16),
31916 => conv_std_logic_vector(21328, 16),
31917 => conv_std_logic_vector(21452, 16),
31918 => conv_std_logic_vector(21576, 16),
31919 => conv_std_logic_vector(21700, 16),
31920 => conv_std_logic_vector(21824, 16),
31921 => conv_std_logic_vector(21948, 16),
31922 => conv_std_logic_vector(22072, 16),
31923 => conv_std_logic_vector(22196, 16),
31924 => conv_std_logic_vector(22320, 16),
31925 => conv_std_logic_vector(22444, 16),
31926 => conv_std_logic_vector(22568, 16),
31927 => conv_std_logic_vector(22692, 16),
31928 => conv_std_logic_vector(22816, 16),
31929 => conv_std_logic_vector(22940, 16),
31930 => conv_std_logic_vector(23064, 16),
31931 => conv_std_logic_vector(23188, 16),
31932 => conv_std_logic_vector(23312, 16),
31933 => conv_std_logic_vector(23436, 16),
31934 => conv_std_logic_vector(23560, 16),
31935 => conv_std_logic_vector(23684, 16),
31936 => conv_std_logic_vector(23808, 16),
31937 => conv_std_logic_vector(23932, 16),
31938 => conv_std_logic_vector(24056, 16),
31939 => conv_std_logic_vector(24180, 16),
31940 => conv_std_logic_vector(24304, 16),
31941 => conv_std_logic_vector(24428, 16),
31942 => conv_std_logic_vector(24552, 16),
31943 => conv_std_logic_vector(24676, 16),
31944 => conv_std_logic_vector(24800, 16),
31945 => conv_std_logic_vector(24924, 16),
31946 => conv_std_logic_vector(25048, 16),
31947 => conv_std_logic_vector(25172, 16),
31948 => conv_std_logic_vector(25296, 16),
31949 => conv_std_logic_vector(25420, 16),
31950 => conv_std_logic_vector(25544, 16),
31951 => conv_std_logic_vector(25668, 16),
31952 => conv_std_logic_vector(25792, 16),
31953 => conv_std_logic_vector(25916, 16),
31954 => conv_std_logic_vector(26040, 16),
31955 => conv_std_logic_vector(26164, 16),
31956 => conv_std_logic_vector(26288, 16),
31957 => conv_std_logic_vector(26412, 16),
31958 => conv_std_logic_vector(26536, 16),
31959 => conv_std_logic_vector(26660, 16),
31960 => conv_std_logic_vector(26784, 16),
31961 => conv_std_logic_vector(26908, 16),
31962 => conv_std_logic_vector(27032, 16),
31963 => conv_std_logic_vector(27156, 16),
31964 => conv_std_logic_vector(27280, 16),
31965 => conv_std_logic_vector(27404, 16),
31966 => conv_std_logic_vector(27528, 16),
31967 => conv_std_logic_vector(27652, 16),
31968 => conv_std_logic_vector(27776, 16),
31969 => conv_std_logic_vector(27900, 16),
31970 => conv_std_logic_vector(28024, 16),
31971 => conv_std_logic_vector(28148, 16),
31972 => conv_std_logic_vector(28272, 16),
31973 => conv_std_logic_vector(28396, 16),
31974 => conv_std_logic_vector(28520, 16),
31975 => conv_std_logic_vector(28644, 16),
31976 => conv_std_logic_vector(28768, 16),
31977 => conv_std_logic_vector(28892, 16),
31978 => conv_std_logic_vector(29016, 16),
31979 => conv_std_logic_vector(29140, 16),
31980 => conv_std_logic_vector(29264, 16),
31981 => conv_std_logic_vector(29388, 16),
31982 => conv_std_logic_vector(29512, 16),
31983 => conv_std_logic_vector(29636, 16),
31984 => conv_std_logic_vector(29760, 16),
31985 => conv_std_logic_vector(29884, 16),
31986 => conv_std_logic_vector(30008, 16),
31987 => conv_std_logic_vector(30132, 16),
31988 => conv_std_logic_vector(30256, 16),
31989 => conv_std_logic_vector(30380, 16),
31990 => conv_std_logic_vector(30504, 16),
31991 => conv_std_logic_vector(30628, 16),
31992 => conv_std_logic_vector(30752, 16),
31993 => conv_std_logic_vector(30876, 16),
31994 => conv_std_logic_vector(31000, 16),
31995 => conv_std_logic_vector(31124, 16),
31996 => conv_std_logic_vector(31248, 16),
31997 => conv_std_logic_vector(31372, 16),
31998 => conv_std_logic_vector(31496, 16),
31999 => conv_std_logic_vector(31620, 16),
32000 => conv_std_logic_vector(0, 16),
32001 => conv_std_logic_vector(125, 16),
32002 => conv_std_logic_vector(250, 16),
32003 => conv_std_logic_vector(375, 16),
32004 => conv_std_logic_vector(500, 16),
32005 => conv_std_logic_vector(625, 16),
32006 => conv_std_logic_vector(750, 16),
32007 => conv_std_logic_vector(875, 16),
32008 => conv_std_logic_vector(1000, 16),
32009 => conv_std_logic_vector(1125, 16),
32010 => conv_std_logic_vector(1250, 16),
32011 => conv_std_logic_vector(1375, 16),
32012 => conv_std_logic_vector(1500, 16),
32013 => conv_std_logic_vector(1625, 16),
32014 => conv_std_logic_vector(1750, 16),
32015 => conv_std_logic_vector(1875, 16),
32016 => conv_std_logic_vector(2000, 16),
32017 => conv_std_logic_vector(2125, 16),
32018 => conv_std_logic_vector(2250, 16),
32019 => conv_std_logic_vector(2375, 16),
32020 => conv_std_logic_vector(2500, 16),
32021 => conv_std_logic_vector(2625, 16),
32022 => conv_std_logic_vector(2750, 16),
32023 => conv_std_logic_vector(2875, 16),
32024 => conv_std_logic_vector(3000, 16),
32025 => conv_std_logic_vector(3125, 16),
32026 => conv_std_logic_vector(3250, 16),
32027 => conv_std_logic_vector(3375, 16),
32028 => conv_std_logic_vector(3500, 16),
32029 => conv_std_logic_vector(3625, 16),
32030 => conv_std_logic_vector(3750, 16),
32031 => conv_std_logic_vector(3875, 16),
32032 => conv_std_logic_vector(4000, 16),
32033 => conv_std_logic_vector(4125, 16),
32034 => conv_std_logic_vector(4250, 16),
32035 => conv_std_logic_vector(4375, 16),
32036 => conv_std_logic_vector(4500, 16),
32037 => conv_std_logic_vector(4625, 16),
32038 => conv_std_logic_vector(4750, 16),
32039 => conv_std_logic_vector(4875, 16),
32040 => conv_std_logic_vector(5000, 16),
32041 => conv_std_logic_vector(5125, 16),
32042 => conv_std_logic_vector(5250, 16),
32043 => conv_std_logic_vector(5375, 16),
32044 => conv_std_logic_vector(5500, 16),
32045 => conv_std_logic_vector(5625, 16),
32046 => conv_std_logic_vector(5750, 16),
32047 => conv_std_logic_vector(5875, 16),
32048 => conv_std_logic_vector(6000, 16),
32049 => conv_std_logic_vector(6125, 16),
32050 => conv_std_logic_vector(6250, 16),
32051 => conv_std_logic_vector(6375, 16),
32052 => conv_std_logic_vector(6500, 16),
32053 => conv_std_logic_vector(6625, 16),
32054 => conv_std_logic_vector(6750, 16),
32055 => conv_std_logic_vector(6875, 16),
32056 => conv_std_logic_vector(7000, 16),
32057 => conv_std_logic_vector(7125, 16),
32058 => conv_std_logic_vector(7250, 16),
32059 => conv_std_logic_vector(7375, 16),
32060 => conv_std_logic_vector(7500, 16),
32061 => conv_std_logic_vector(7625, 16),
32062 => conv_std_logic_vector(7750, 16),
32063 => conv_std_logic_vector(7875, 16),
32064 => conv_std_logic_vector(8000, 16),
32065 => conv_std_logic_vector(8125, 16),
32066 => conv_std_logic_vector(8250, 16),
32067 => conv_std_logic_vector(8375, 16),
32068 => conv_std_logic_vector(8500, 16),
32069 => conv_std_logic_vector(8625, 16),
32070 => conv_std_logic_vector(8750, 16),
32071 => conv_std_logic_vector(8875, 16),
32072 => conv_std_logic_vector(9000, 16),
32073 => conv_std_logic_vector(9125, 16),
32074 => conv_std_logic_vector(9250, 16),
32075 => conv_std_logic_vector(9375, 16),
32076 => conv_std_logic_vector(9500, 16),
32077 => conv_std_logic_vector(9625, 16),
32078 => conv_std_logic_vector(9750, 16),
32079 => conv_std_logic_vector(9875, 16),
32080 => conv_std_logic_vector(10000, 16),
32081 => conv_std_logic_vector(10125, 16),
32082 => conv_std_logic_vector(10250, 16),
32083 => conv_std_logic_vector(10375, 16),
32084 => conv_std_logic_vector(10500, 16),
32085 => conv_std_logic_vector(10625, 16),
32086 => conv_std_logic_vector(10750, 16),
32087 => conv_std_logic_vector(10875, 16),
32088 => conv_std_logic_vector(11000, 16),
32089 => conv_std_logic_vector(11125, 16),
32090 => conv_std_logic_vector(11250, 16),
32091 => conv_std_logic_vector(11375, 16),
32092 => conv_std_logic_vector(11500, 16),
32093 => conv_std_logic_vector(11625, 16),
32094 => conv_std_logic_vector(11750, 16),
32095 => conv_std_logic_vector(11875, 16),
32096 => conv_std_logic_vector(12000, 16),
32097 => conv_std_logic_vector(12125, 16),
32098 => conv_std_logic_vector(12250, 16),
32099 => conv_std_logic_vector(12375, 16),
32100 => conv_std_logic_vector(12500, 16),
32101 => conv_std_logic_vector(12625, 16),
32102 => conv_std_logic_vector(12750, 16),
32103 => conv_std_logic_vector(12875, 16),
32104 => conv_std_logic_vector(13000, 16),
32105 => conv_std_logic_vector(13125, 16),
32106 => conv_std_logic_vector(13250, 16),
32107 => conv_std_logic_vector(13375, 16),
32108 => conv_std_logic_vector(13500, 16),
32109 => conv_std_logic_vector(13625, 16),
32110 => conv_std_logic_vector(13750, 16),
32111 => conv_std_logic_vector(13875, 16),
32112 => conv_std_logic_vector(14000, 16),
32113 => conv_std_logic_vector(14125, 16),
32114 => conv_std_logic_vector(14250, 16),
32115 => conv_std_logic_vector(14375, 16),
32116 => conv_std_logic_vector(14500, 16),
32117 => conv_std_logic_vector(14625, 16),
32118 => conv_std_logic_vector(14750, 16),
32119 => conv_std_logic_vector(14875, 16),
32120 => conv_std_logic_vector(15000, 16),
32121 => conv_std_logic_vector(15125, 16),
32122 => conv_std_logic_vector(15250, 16),
32123 => conv_std_logic_vector(15375, 16),
32124 => conv_std_logic_vector(15500, 16),
32125 => conv_std_logic_vector(15625, 16),
32126 => conv_std_logic_vector(15750, 16),
32127 => conv_std_logic_vector(15875, 16),
32128 => conv_std_logic_vector(16000, 16),
32129 => conv_std_logic_vector(16125, 16),
32130 => conv_std_logic_vector(16250, 16),
32131 => conv_std_logic_vector(16375, 16),
32132 => conv_std_logic_vector(16500, 16),
32133 => conv_std_logic_vector(16625, 16),
32134 => conv_std_logic_vector(16750, 16),
32135 => conv_std_logic_vector(16875, 16),
32136 => conv_std_logic_vector(17000, 16),
32137 => conv_std_logic_vector(17125, 16),
32138 => conv_std_logic_vector(17250, 16),
32139 => conv_std_logic_vector(17375, 16),
32140 => conv_std_logic_vector(17500, 16),
32141 => conv_std_logic_vector(17625, 16),
32142 => conv_std_logic_vector(17750, 16),
32143 => conv_std_logic_vector(17875, 16),
32144 => conv_std_logic_vector(18000, 16),
32145 => conv_std_logic_vector(18125, 16),
32146 => conv_std_logic_vector(18250, 16),
32147 => conv_std_logic_vector(18375, 16),
32148 => conv_std_logic_vector(18500, 16),
32149 => conv_std_logic_vector(18625, 16),
32150 => conv_std_logic_vector(18750, 16),
32151 => conv_std_logic_vector(18875, 16),
32152 => conv_std_logic_vector(19000, 16),
32153 => conv_std_logic_vector(19125, 16),
32154 => conv_std_logic_vector(19250, 16),
32155 => conv_std_logic_vector(19375, 16),
32156 => conv_std_logic_vector(19500, 16),
32157 => conv_std_logic_vector(19625, 16),
32158 => conv_std_logic_vector(19750, 16),
32159 => conv_std_logic_vector(19875, 16),
32160 => conv_std_logic_vector(20000, 16),
32161 => conv_std_logic_vector(20125, 16),
32162 => conv_std_logic_vector(20250, 16),
32163 => conv_std_logic_vector(20375, 16),
32164 => conv_std_logic_vector(20500, 16),
32165 => conv_std_logic_vector(20625, 16),
32166 => conv_std_logic_vector(20750, 16),
32167 => conv_std_logic_vector(20875, 16),
32168 => conv_std_logic_vector(21000, 16),
32169 => conv_std_logic_vector(21125, 16),
32170 => conv_std_logic_vector(21250, 16),
32171 => conv_std_logic_vector(21375, 16),
32172 => conv_std_logic_vector(21500, 16),
32173 => conv_std_logic_vector(21625, 16),
32174 => conv_std_logic_vector(21750, 16),
32175 => conv_std_logic_vector(21875, 16),
32176 => conv_std_logic_vector(22000, 16),
32177 => conv_std_logic_vector(22125, 16),
32178 => conv_std_logic_vector(22250, 16),
32179 => conv_std_logic_vector(22375, 16),
32180 => conv_std_logic_vector(22500, 16),
32181 => conv_std_logic_vector(22625, 16),
32182 => conv_std_logic_vector(22750, 16),
32183 => conv_std_logic_vector(22875, 16),
32184 => conv_std_logic_vector(23000, 16),
32185 => conv_std_logic_vector(23125, 16),
32186 => conv_std_logic_vector(23250, 16),
32187 => conv_std_logic_vector(23375, 16),
32188 => conv_std_logic_vector(23500, 16),
32189 => conv_std_logic_vector(23625, 16),
32190 => conv_std_logic_vector(23750, 16),
32191 => conv_std_logic_vector(23875, 16),
32192 => conv_std_logic_vector(24000, 16),
32193 => conv_std_logic_vector(24125, 16),
32194 => conv_std_logic_vector(24250, 16),
32195 => conv_std_logic_vector(24375, 16),
32196 => conv_std_logic_vector(24500, 16),
32197 => conv_std_logic_vector(24625, 16),
32198 => conv_std_logic_vector(24750, 16),
32199 => conv_std_logic_vector(24875, 16),
32200 => conv_std_logic_vector(25000, 16),
32201 => conv_std_logic_vector(25125, 16),
32202 => conv_std_logic_vector(25250, 16),
32203 => conv_std_logic_vector(25375, 16),
32204 => conv_std_logic_vector(25500, 16),
32205 => conv_std_logic_vector(25625, 16),
32206 => conv_std_logic_vector(25750, 16),
32207 => conv_std_logic_vector(25875, 16),
32208 => conv_std_logic_vector(26000, 16),
32209 => conv_std_logic_vector(26125, 16),
32210 => conv_std_logic_vector(26250, 16),
32211 => conv_std_logic_vector(26375, 16),
32212 => conv_std_logic_vector(26500, 16),
32213 => conv_std_logic_vector(26625, 16),
32214 => conv_std_logic_vector(26750, 16),
32215 => conv_std_logic_vector(26875, 16),
32216 => conv_std_logic_vector(27000, 16),
32217 => conv_std_logic_vector(27125, 16),
32218 => conv_std_logic_vector(27250, 16),
32219 => conv_std_logic_vector(27375, 16),
32220 => conv_std_logic_vector(27500, 16),
32221 => conv_std_logic_vector(27625, 16),
32222 => conv_std_logic_vector(27750, 16),
32223 => conv_std_logic_vector(27875, 16),
32224 => conv_std_logic_vector(28000, 16),
32225 => conv_std_logic_vector(28125, 16),
32226 => conv_std_logic_vector(28250, 16),
32227 => conv_std_logic_vector(28375, 16),
32228 => conv_std_logic_vector(28500, 16),
32229 => conv_std_logic_vector(28625, 16),
32230 => conv_std_logic_vector(28750, 16),
32231 => conv_std_logic_vector(28875, 16),
32232 => conv_std_logic_vector(29000, 16),
32233 => conv_std_logic_vector(29125, 16),
32234 => conv_std_logic_vector(29250, 16),
32235 => conv_std_logic_vector(29375, 16),
32236 => conv_std_logic_vector(29500, 16),
32237 => conv_std_logic_vector(29625, 16),
32238 => conv_std_logic_vector(29750, 16),
32239 => conv_std_logic_vector(29875, 16),
32240 => conv_std_logic_vector(30000, 16),
32241 => conv_std_logic_vector(30125, 16),
32242 => conv_std_logic_vector(30250, 16),
32243 => conv_std_logic_vector(30375, 16),
32244 => conv_std_logic_vector(30500, 16),
32245 => conv_std_logic_vector(30625, 16),
32246 => conv_std_logic_vector(30750, 16),
32247 => conv_std_logic_vector(30875, 16),
32248 => conv_std_logic_vector(31000, 16),
32249 => conv_std_logic_vector(31125, 16),
32250 => conv_std_logic_vector(31250, 16),
32251 => conv_std_logic_vector(31375, 16),
32252 => conv_std_logic_vector(31500, 16),
32253 => conv_std_logic_vector(31625, 16),
32254 => conv_std_logic_vector(31750, 16),
32255 => conv_std_logic_vector(31875, 16),
32256 => conv_std_logic_vector(0, 16),
32257 => conv_std_logic_vector(126, 16),
32258 => conv_std_logic_vector(252, 16),
32259 => conv_std_logic_vector(378, 16),
32260 => conv_std_logic_vector(504, 16),
32261 => conv_std_logic_vector(630, 16),
32262 => conv_std_logic_vector(756, 16),
32263 => conv_std_logic_vector(882, 16),
32264 => conv_std_logic_vector(1008, 16),
32265 => conv_std_logic_vector(1134, 16),
32266 => conv_std_logic_vector(1260, 16),
32267 => conv_std_logic_vector(1386, 16),
32268 => conv_std_logic_vector(1512, 16),
32269 => conv_std_logic_vector(1638, 16),
32270 => conv_std_logic_vector(1764, 16),
32271 => conv_std_logic_vector(1890, 16),
32272 => conv_std_logic_vector(2016, 16),
32273 => conv_std_logic_vector(2142, 16),
32274 => conv_std_logic_vector(2268, 16),
32275 => conv_std_logic_vector(2394, 16),
32276 => conv_std_logic_vector(2520, 16),
32277 => conv_std_logic_vector(2646, 16),
32278 => conv_std_logic_vector(2772, 16),
32279 => conv_std_logic_vector(2898, 16),
32280 => conv_std_logic_vector(3024, 16),
32281 => conv_std_logic_vector(3150, 16),
32282 => conv_std_logic_vector(3276, 16),
32283 => conv_std_logic_vector(3402, 16),
32284 => conv_std_logic_vector(3528, 16),
32285 => conv_std_logic_vector(3654, 16),
32286 => conv_std_logic_vector(3780, 16),
32287 => conv_std_logic_vector(3906, 16),
32288 => conv_std_logic_vector(4032, 16),
32289 => conv_std_logic_vector(4158, 16),
32290 => conv_std_logic_vector(4284, 16),
32291 => conv_std_logic_vector(4410, 16),
32292 => conv_std_logic_vector(4536, 16),
32293 => conv_std_logic_vector(4662, 16),
32294 => conv_std_logic_vector(4788, 16),
32295 => conv_std_logic_vector(4914, 16),
32296 => conv_std_logic_vector(5040, 16),
32297 => conv_std_logic_vector(5166, 16),
32298 => conv_std_logic_vector(5292, 16),
32299 => conv_std_logic_vector(5418, 16),
32300 => conv_std_logic_vector(5544, 16),
32301 => conv_std_logic_vector(5670, 16),
32302 => conv_std_logic_vector(5796, 16),
32303 => conv_std_logic_vector(5922, 16),
32304 => conv_std_logic_vector(6048, 16),
32305 => conv_std_logic_vector(6174, 16),
32306 => conv_std_logic_vector(6300, 16),
32307 => conv_std_logic_vector(6426, 16),
32308 => conv_std_logic_vector(6552, 16),
32309 => conv_std_logic_vector(6678, 16),
32310 => conv_std_logic_vector(6804, 16),
32311 => conv_std_logic_vector(6930, 16),
32312 => conv_std_logic_vector(7056, 16),
32313 => conv_std_logic_vector(7182, 16),
32314 => conv_std_logic_vector(7308, 16),
32315 => conv_std_logic_vector(7434, 16),
32316 => conv_std_logic_vector(7560, 16),
32317 => conv_std_logic_vector(7686, 16),
32318 => conv_std_logic_vector(7812, 16),
32319 => conv_std_logic_vector(7938, 16),
32320 => conv_std_logic_vector(8064, 16),
32321 => conv_std_logic_vector(8190, 16),
32322 => conv_std_logic_vector(8316, 16),
32323 => conv_std_logic_vector(8442, 16),
32324 => conv_std_logic_vector(8568, 16),
32325 => conv_std_logic_vector(8694, 16),
32326 => conv_std_logic_vector(8820, 16),
32327 => conv_std_logic_vector(8946, 16),
32328 => conv_std_logic_vector(9072, 16),
32329 => conv_std_logic_vector(9198, 16),
32330 => conv_std_logic_vector(9324, 16),
32331 => conv_std_logic_vector(9450, 16),
32332 => conv_std_logic_vector(9576, 16),
32333 => conv_std_logic_vector(9702, 16),
32334 => conv_std_logic_vector(9828, 16),
32335 => conv_std_logic_vector(9954, 16),
32336 => conv_std_logic_vector(10080, 16),
32337 => conv_std_logic_vector(10206, 16),
32338 => conv_std_logic_vector(10332, 16),
32339 => conv_std_logic_vector(10458, 16),
32340 => conv_std_logic_vector(10584, 16),
32341 => conv_std_logic_vector(10710, 16),
32342 => conv_std_logic_vector(10836, 16),
32343 => conv_std_logic_vector(10962, 16),
32344 => conv_std_logic_vector(11088, 16),
32345 => conv_std_logic_vector(11214, 16),
32346 => conv_std_logic_vector(11340, 16),
32347 => conv_std_logic_vector(11466, 16),
32348 => conv_std_logic_vector(11592, 16),
32349 => conv_std_logic_vector(11718, 16),
32350 => conv_std_logic_vector(11844, 16),
32351 => conv_std_logic_vector(11970, 16),
32352 => conv_std_logic_vector(12096, 16),
32353 => conv_std_logic_vector(12222, 16),
32354 => conv_std_logic_vector(12348, 16),
32355 => conv_std_logic_vector(12474, 16),
32356 => conv_std_logic_vector(12600, 16),
32357 => conv_std_logic_vector(12726, 16),
32358 => conv_std_logic_vector(12852, 16),
32359 => conv_std_logic_vector(12978, 16),
32360 => conv_std_logic_vector(13104, 16),
32361 => conv_std_logic_vector(13230, 16),
32362 => conv_std_logic_vector(13356, 16),
32363 => conv_std_logic_vector(13482, 16),
32364 => conv_std_logic_vector(13608, 16),
32365 => conv_std_logic_vector(13734, 16),
32366 => conv_std_logic_vector(13860, 16),
32367 => conv_std_logic_vector(13986, 16),
32368 => conv_std_logic_vector(14112, 16),
32369 => conv_std_logic_vector(14238, 16),
32370 => conv_std_logic_vector(14364, 16),
32371 => conv_std_logic_vector(14490, 16),
32372 => conv_std_logic_vector(14616, 16),
32373 => conv_std_logic_vector(14742, 16),
32374 => conv_std_logic_vector(14868, 16),
32375 => conv_std_logic_vector(14994, 16),
32376 => conv_std_logic_vector(15120, 16),
32377 => conv_std_logic_vector(15246, 16),
32378 => conv_std_logic_vector(15372, 16),
32379 => conv_std_logic_vector(15498, 16),
32380 => conv_std_logic_vector(15624, 16),
32381 => conv_std_logic_vector(15750, 16),
32382 => conv_std_logic_vector(15876, 16),
32383 => conv_std_logic_vector(16002, 16),
32384 => conv_std_logic_vector(16128, 16),
32385 => conv_std_logic_vector(16254, 16),
32386 => conv_std_logic_vector(16380, 16),
32387 => conv_std_logic_vector(16506, 16),
32388 => conv_std_logic_vector(16632, 16),
32389 => conv_std_logic_vector(16758, 16),
32390 => conv_std_logic_vector(16884, 16),
32391 => conv_std_logic_vector(17010, 16),
32392 => conv_std_logic_vector(17136, 16),
32393 => conv_std_logic_vector(17262, 16),
32394 => conv_std_logic_vector(17388, 16),
32395 => conv_std_logic_vector(17514, 16),
32396 => conv_std_logic_vector(17640, 16),
32397 => conv_std_logic_vector(17766, 16),
32398 => conv_std_logic_vector(17892, 16),
32399 => conv_std_logic_vector(18018, 16),
32400 => conv_std_logic_vector(18144, 16),
32401 => conv_std_logic_vector(18270, 16),
32402 => conv_std_logic_vector(18396, 16),
32403 => conv_std_logic_vector(18522, 16),
32404 => conv_std_logic_vector(18648, 16),
32405 => conv_std_logic_vector(18774, 16),
32406 => conv_std_logic_vector(18900, 16),
32407 => conv_std_logic_vector(19026, 16),
32408 => conv_std_logic_vector(19152, 16),
32409 => conv_std_logic_vector(19278, 16),
32410 => conv_std_logic_vector(19404, 16),
32411 => conv_std_logic_vector(19530, 16),
32412 => conv_std_logic_vector(19656, 16),
32413 => conv_std_logic_vector(19782, 16),
32414 => conv_std_logic_vector(19908, 16),
32415 => conv_std_logic_vector(20034, 16),
32416 => conv_std_logic_vector(20160, 16),
32417 => conv_std_logic_vector(20286, 16),
32418 => conv_std_logic_vector(20412, 16),
32419 => conv_std_logic_vector(20538, 16),
32420 => conv_std_logic_vector(20664, 16),
32421 => conv_std_logic_vector(20790, 16),
32422 => conv_std_logic_vector(20916, 16),
32423 => conv_std_logic_vector(21042, 16),
32424 => conv_std_logic_vector(21168, 16),
32425 => conv_std_logic_vector(21294, 16),
32426 => conv_std_logic_vector(21420, 16),
32427 => conv_std_logic_vector(21546, 16),
32428 => conv_std_logic_vector(21672, 16),
32429 => conv_std_logic_vector(21798, 16),
32430 => conv_std_logic_vector(21924, 16),
32431 => conv_std_logic_vector(22050, 16),
32432 => conv_std_logic_vector(22176, 16),
32433 => conv_std_logic_vector(22302, 16),
32434 => conv_std_logic_vector(22428, 16),
32435 => conv_std_logic_vector(22554, 16),
32436 => conv_std_logic_vector(22680, 16),
32437 => conv_std_logic_vector(22806, 16),
32438 => conv_std_logic_vector(22932, 16),
32439 => conv_std_logic_vector(23058, 16),
32440 => conv_std_logic_vector(23184, 16),
32441 => conv_std_logic_vector(23310, 16),
32442 => conv_std_logic_vector(23436, 16),
32443 => conv_std_logic_vector(23562, 16),
32444 => conv_std_logic_vector(23688, 16),
32445 => conv_std_logic_vector(23814, 16),
32446 => conv_std_logic_vector(23940, 16),
32447 => conv_std_logic_vector(24066, 16),
32448 => conv_std_logic_vector(24192, 16),
32449 => conv_std_logic_vector(24318, 16),
32450 => conv_std_logic_vector(24444, 16),
32451 => conv_std_logic_vector(24570, 16),
32452 => conv_std_logic_vector(24696, 16),
32453 => conv_std_logic_vector(24822, 16),
32454 => conv_std_logic_vector(24948, 16),
32455 => conv_std_logic_vector(25074, 16),
32456 => conv_std_logic_vector(25200, 16),
32457 => conv_std_logic_vector(25326, 16),
32458 => conv_std_logic_vector(25452, 16),
32459 => conv_std_logic_vector(25578, 16),
32460 => conv_std_logic_vector(25704, 16),
32461 => conv_std_logic_vector(25830, 16),
32462 => conv_std_logic_vector(25956, 16),
32463 => conv_std_logic_vector(26082, 16),
32464 => conv_std_logic_vector(26208, 16),
32465 => conv_std_logic_vector(26334, 16),
32466 => conv_std_logic_vector(26460, 16),
32467 => conv_std_logic_vector(26586, 16),
32468 => conv_std_logic_vector(26712, 16),
32469 => conv_std_logic_vector(26838, 16),
32470 => conv_std_logic_vector(26964, 16),
32471 => conv_std_logic_vector(27090, 16),
32472 => conv_std_logic_vector(27216, 16),
32473 => conv_std_logic_vector(27342, 16),
32474 => conv_std_logic_vector(27468, 16),
32475 => conv_std_logic_vector(27594, 16),
32476 => conv_std_logic_vector(27720, 16),
32477 => conv_std_logic_vector(27846, 16),
32478 => conv_std_logic_vector(27972, 16),
32479 => conv_std_logic_vector(28098, 16),
32480 => conv_std_logic_vector(28224, 16),
32481 => conv_std_logic_vector(28350, 16),
32482 => conv_std_logic_vector(28476, 16),
32483 => conv_std_logic_vector(28602, 16),
32484 => conv_std_logic_vector(28728, 16),
32485 => conv_std_logic_vector(28854, 16),
32486 => conv_std_logic_vector(28980, 16),
32487 => conv_std_logic_vector(29106, 16),
32488 => conv_std_logic_vector(29232, 16),
32489 => conv_std_logic_vector(29358, 16),
32490 => conv_std_logic_vector(29484, 16),
32491 => conv_std_logic_vector(29610, 16),
32492 => conv_std_logic_vector(29736, 16),
32493 => conv_std_logic_vector(29862, 16),
32494 => conv_std_logic_vector(29988, 16),
32495 => conv_std_logic_vector(30114, 16),
32496 => conv_std_logic_vector(30240, 16),
32497 => conv_std_logic_vector(30366, 16),
32498 => conv_std_logic_vector(30492, 16),
32499 => conv_std_logic_vector(30618, 16),
32500 => conv_std_logic_vector(30744, 16),
32501 => conv_std_logic_vector(30870, 16),
32502 => conv_std_logic_vector(30996, 16),
32503 => conv_std_logic_vector(31122, 16),
32504 => conv_std_logic_vector(31248, 16),
32505 => conv_std_logic_vector(31374, 16),
32506 => conv_std_logic_vector(31500, 16),
32507 => conv_std_logic_vector(31626, 16),
32508 => conv_std_logic_vector(31752, 16),
32509 => conv_std_logic_vector(31878, 16),
32510 => conv_std_logic_vector(32004, 16),
32511 => conv_std_logic_vector(32130, 16),
32512 => conv_std_logic_vector(0, 16),
32513 => conv_std_logic_vector(127, 16),
32514 => conv_std_logic_vector(254, 16),
32515 => conv_std_logic_vector(381, 16),
32516 => conv_std_logic_vector(508, 16),
32517 => conv_std_logic_vector(635, 16),
32518 => conv_std_logic_vector(762, 16),
32519 => conv_std_logic_vector(889, 16),
32520 => conv_std_logic_vector(1016, 16),
32521 => conv_std_logic_vector(1143, 16),
32522 => conv_std_logic_vector(1270, 16),
32523 => conv_std_logic_vector(1397, 16),
32524 => conv_std_logic_vector(1524, 16),
32525 => conv_std_logic_vector(1651, 16),
32526 => conv_std_logic_vector(1778, 16),
32527 => conv_std_logic_vector(1905, 16),
32528 => conv_std_logic_vector(2032, 16),
32529 => conv_std_logic_vector(2159, 16),
32530 => conv_std_logic_vector(2286, 16),
32531 => conv_std_logic_vector(2413, 16),
32532 => conv_std_logic_vector(2540, 16),
32533 => conv_std_logic_vector(2667, 16),
32534 => conv_std_logic_vector(2794, 16),
32535 => conv_std_logic_vector(2921, 16),
32536 => conv_std_logic_vector(3048, 16),
32537 => conv_std_logic_vector(3175, 16),
32538 => conv_std_logic_vector(3302, 16),
32539 => conv_std_logic_vector(3429, 16),
32540 => conv_std_logic_vector(3556, 16),
32541 => conv_std_logic_vector(3683, 16),
32542 => conv_std_logic_vector(3810, 16),
32543 => conv_std_logic_vector(3937, 16),
32544 => conv_std_logic_vector(4064, 16),
32545 => conv_std_logic_vector(4191, 16),
32546 => conv_std_logic_vector(4318, 16),
32547 => conv_std_logic_vector(4445, 16),
32548 => conv_std_logic_vector(4572, 16),
32549 => conv_std_logic_vector(4699, 16),
32550 => conv_std_logic_vector(4826, 16),
32551 => conv_std_logic_vector(4953, 16),
32552 => conv_std_logic_vector(5080, 16),
32553 => conv_std_logic_vector(5207, 16),
32554 => conv_std_logic_vector(5334, 16),
32555 => conv_std_logic_vector(5461, 16),
32556 => conv_std_logic_vector(5588, 16),
32557 => conv_std_logic_vector(5715, 16),
32558 => conv_std_logic_vector(5842, 16),
32559 => conv_std_logic_vector(5969, 16),
32560 => conv_std_logic_vector(6096, 16),
32561 => conv_std_logic_vector(6223, 16),
32562 => conv_std_logic_vector(6350, 16),
32563 => conv_std_logic_vector(6477, 16),
32564 => conv_std_logic_vector(6604, 16),
32565 => conv_std_logic_vector(6731, 16),
32566 => conv_std_logic_vector(6858, 16),
32567 => conv_std_logic_vector(6985, 16),
32568 => conv_std_logic_vector(7112, 16),
32569 => conv_std_logic_vector(7239, 16),
32570 => conv_std_logic_vector(7366, 16),
32571 => conv_std_logic_vector(7493, 16),
32572 => conv_std_logic_vector(7620, 16),
32573 => conv_std_logic_vector(7747, 16),
32574 => conv_std_logic_vector(7874, 16),
32575 => conv_std_logic_vector(8001, 16),
32576 => conv_std_logic_vector(8128, 16),
32577 => conv_std_logic_vector(8255, 16),
32578 => conv_std_logic_vector(8382, 16),
32579 => conv_std_logic_vector(8509, 16),
32580 => conv_std_logic_vector(8636, 16),
32581 => conv_std_logic_vector(8763, 16),
32582 => conv_std_logic_vector(8890, 16),
32583 => conv_std_logic_vector(9017, 16),
32584 => conv_std_logic_vector(9144, 16),
32585 => conv_std_logic_vector(9271, 16),
32586 => conv_std_logic_vector(9398, 16),
32587 => conv_std_logic_vector(9525, 16),
32588 => conv_std_logic_vector(9652, 16),
32589 => conv_std_logic_vector(9779, 16),
32590 => conv_std_logic_vector(9906, 16),
32591 => conv_std_logic_vector(10033, 16),
32592 => conv_std_logic_vector(10160, 16),
32593 => conv_std_logic_vector(10287, 16),
32594 => conv_std_logic_vector(10414, 16),
32595 => conv_std_logic_vector(10541, 16),
32596 => conv_std_logic_vector(10668, 16),
32597 => conv_std_logic_vector(10795, 16),
32598 => conv_std_logic_vector(10922, 16),
32599 => conv_std_logic_vector(11049, 16),
32600 => conv_std_logic_vector(11176, 16),
32601 => conv_std_logic_vector(11303, 16),
32602 => conv_std_logic_vector(11430, 16),
32603 => conv_std_logic_vector(11557, 16),
32604 => conv_std_logic_vector(11684, 16),
32605 => conv_std_logic_vector(11811, 16),
32606 => conv_std_logic_vector(11938, 16),
32607 => conv_std_logic_vector(12065, 16),
32608 => conv_std_logic_vector(12192, 16),
32609 => conv_std_logic_vector(12319, 16),
32610 => conv_std_logic_vector(12446, 16),
32611 => conv_std_logic_vector(12573, 16),
32612 => conv_std_logic_vector(12700, 16),
32613 => conv_std_logic_vector(12827, 16),
32614 => conv_std_logic_vector(12954, 16),
32615 => conv_std_logic_vector(13081, 16),
32616 => conv_std_logic_vector(13208, 16),
32617 => conv_std_logic_vector(13335, 16),
32618 => conv_std_logic_vector(13462, 16),
32619 => conv_std_logic_vector(13589, 16),
32620 => conv_std_logic_vector(13716, 16),
32621 => conv_std_logic_vector(13843, 16),
32622 => conv_std_logic_vector(13970, 16),
32623 => conv_std_logic_vector(14097, 16),
32624 => conv_std_logic_vector(14224, 16),
32625 => conv_std_logic_vector(14351, 16),
32626 => conv_std_logic_vector(14478, 16),
32627 => conv_std_logic_vector(14605, 16),
32628 => conv_std_logic_vector(14732, 16),
32629 => conv_std_logic_vector(14859, 16),
32630 => conv_std_logic_vector(14986, 16),
32631 => conv_std_logic_vector(15113, 16),
32632 => conv_std_logic_vector(15240, 16),
32633 => conv_std_logic_vector(15367, 16),
32634 => conv_std_logic_vector(15494, 16),
32635 => conv_std_logic_vector(15621, 16),
32636 => conv_std_logic_vector(15748, 16),
32637 => conv_std_logic_vector(15875, 16),
32638 => conv_std_logic_vector(16002, 16),
32639 => conv_std_logic_vector(16129, 16),
32640 => conv_std_logic_vector(16256, 16),
32641 => conv_std_logic_vector(16383, 16),
32642 => conv_std_logic_vector(16510, 16),
32643 => conv_std_logic_vector(16637, 16),
32644 => conv_std_logic_vector(16764, 16),
32645 => conv_std_logic_vector(16891, 16),
32646 => conv_std_logic_vector(17018, 16),
32647 => conv_std_logic_vector(17145, 16),
32648 => conv_std_logic_vector(17272, 16),
32649 => conv_std_logic_vector(17399, 16),
32650 => conv_std_logic_vector(17526, 16),
32651 => conv_std_logic_vector(17653, 16),
32652 => conv_std_logic_vector(17780, 16),
32653 => conv_std_logic_vector(17907, 16),
32654 => conv_std_logic_vector(18034, 16),
32655 => conv_std_logic_vector(18161, 16),
32656 => conv_std_logic_vector(18288, 16),
32657 => conv_std_logic_vector(18415, 16),
32658 => conv_std_logic_vector(18542, 16),
32659 => conv_std_logic_vector(18669, 16),
32660 => conv_std_logic_vector(18796, 16),
32661 => conv_std_logic_vector(18923, 16),
32662 => conv_std_logic_vector(19050, 16),
32663 => conv_std_logic_vector(19177, 16),
32664 => conv_std_logic_vector(19304, 16),
32665 => conv_std_logic_vector(19431, 16),
32666 => conv_std_logic_vector(19558, 16),
32667 => conv_std_logic_vector(19685, 16),
32668 => conv_std_logic_vector(19812, 16),
32669 => conv_std_logic_vector(19939, 16),
32670 => conv_std_logic_vector(20066, 16),
32671 => conv_std_logic_vector(20193, 16),
32672 => conv_std_logic_vector(20320, 16),
32673 => conv_std_logic_vector(20447, 16),
32674 => conv_std_logic_vector(20574, 16),
32675 => conv_std_logic_vector(20701, 16),
32676 => conv_std_logic_vector(20828, 16),
32677 => conv_std_logic_vector(20955, 16),
32678 => conv_std_logic_vector(21082, 16),
32679 => conv_std_logic_vector(21209, 16),
32680 => conv_std_logic_vector(21336, 16),
32681 => conv_std_logic_vector(21463, 16),
32682 => conv_std_logic_vector(21590, 16),
32683 => conv_std_logic_vector(21717, 16),
32684 => conv_std_logic_vector(21844, 16),
32685 => conv_std_logic_vector(21971, 16),
32686 => conv_std_logic_vector(22098, 16),
32687 => conv_std_logic_vector(22225, 16),
32688 => conv_std_logic_vector(22352, 16),
32689 => conv_std_logic_vector(22479, 16),
32690 => conv_std_logic_vector(22606, 16),
32691 => conv_std_logic_vector(22733, 16),
32692 => conv_std_logic_vector(22860, 16),
32693 => conv_std_logic_vector(22987, 16),
32694 => conv_std_logic_vector(23114, 16),
32695 => conv_std_logic_vector(23241, 16),
32696 => conv_std_logic_vector(23368, 16),
32697 => conv_std_logic_vector(23495, 16),
32698 => conv_std_logic_vector(23622, 16),
32699 => conv_std_logic_vector(23749, 16),
32700 => conv_std_logic_vector(23876, 16),
32701 => conv_std_logic_vector(24003, 16),
32702 => conv_std_logic_vector(24130, 16),
32703 => conv_std_logic_vector(24257, 16),
32704 => conv_std_logic_vector(24384, 16),
32705 => conv_std_logic_vector(24511, 16),
32706 => conv_std_logic_vector(24638, 16),
32707 => conv_std_logic_vector(24765, 16),
32708 => conv_std_logic_vector(24892, 16),
32709 => conv_std_logic_vector(25019, 16),
32710 => conv_std_logic_vector(25146, 16),
32711 => conv_std_logic_vector(25273, 16),
32712 => conv_std_logic_vector(25400, 16),
32713 => conv_std_logic_vector(25527, 16),
32714 => conv_std_logic_vector(25654, 16),
32715 => conv_std_logic_vector(25781, 16),
32716 => conv_std_logic_vector(25908, 16),
32717 => conv_std_logic_vector(26035, 16),
32718 => conv_std_logic_vector(26162, 16),
32719 => conv_std_logic_vector(26289, 16),
32720 => conv_std_logic_vector(26416, 16),
32721 => conv_std_logic_vector(26543, 16),
32722 => conv_std_logic_vector(26670, 16),
32723 => conv_std_logic_vector(26797, 16),
32724 => conv_std_logic_vector(26924, 16),
32725 => conv_std_logic_vector(27051, 16),
32726 => conv_std_logic_vector(27178, 16),
32727 => conv_std_logic_vector(27305, 16),
32728 => conv_std_logic_vector(27432, 16),
32729 => conv_std_logic_vector(27559, 16),
32730 => conv_std_logic_vector(27686, 16),
32731 => conv_std_logic_vector(27813, 16),
32732 => conv_std_logic_vector(27940, 16),
32733 => conv_std_logic_vector(28067, 16),
32734 => conv_std_logic_vector(28194, 16),
32735 => conv_std_logic_vector(28321, 16),
32736 => conv_std_logic_vector(28448, 16),
32737 => conv_std_logic_vector(28575, 16),
32738 => conv_std_logic_vector(28702, 16),
32739 => conv_std_logic_vector(28829, 16),
32740 => conv_std_logic_vector(28956, 16),
32741 => conv_std_logic_vector(29083, 16),
32742 => conv_std_logic_vector(29210, 16),
32743 => conv_std_logic_vector(29337, 16),
32744 => conv_std_logic_vector(29464, 16),
32745 => conv_std_logic_vector(29591, 16),
32746 => conv_std_logic_vector(29718, 16),
32747 => conv_std_logic_vector(29845, 16),
32748 => conv_std_logic_vector(29972, 16),
32749 => conv_std_logic_vector(30099, 16),
32750 => conv_std_logic_vector(30226, 16),
32751 => conv_std_logic_vector(30353, 16),
32752 => conv_std_logic_vector(30480, 16),
32753 => conv_std_logic_vector(30607, 16),
32754 => conv_std_logic_vector(30734, 16),
32755 => conv_std_logic_vector(30861, 16),
32756 => conv_std_logic_vector(30988, 16),
32757 => conv_std_logic_vector(31115, 16),
32758 => conv_std_logic_vector(31242, 16),
32759 => conv_std_logic_vector(31369, 16),
32760 => conv_std_logic_vector(31496, 16),
32761 => conv_std_logic_vector(31623, 16),
32762 => conv_std_logic_vector(31750, 16),
32763 => conv_std_logic_vector(31877, 16),
32764 => conv_std_logic_vector(32004, 16),
32765 => conv_std_logic_vector(32131, 16),
32766 => conv_std_logic_vector(32258, 16),
32767 => conv_std_logic_vector(32385, 16),
32768 => conv_std_logic_vector(0, 16),
32769 => conv_std_logic_vector(128, 16),
32770 => conv_std_logic_vector(256, 16),
32771 => conv_std_logic_vector(384, 16),
32772 => conv_std_logic_vector(512, 16),
32773 => conv_std_logic_vector(640, 16),
32774 => conv_std_logic_vector(768, 16),
32775 => conv_std_logic_vector(896, 16),
32776 => conv_std_logic_vector(1024, 16),
32777 => conv_std_logic_vector(1152, 16),
32778 => conv_std_logic_vector(1280, 16),
32779 => conv_std_logic_vector(1408, 16),
32780 => conv_std_logic_vector(1536, 16),
32781 => conv_std_logic_vector(1664, 16),
32782 => conv_std_logic_vector(1792, 16),
32783 => conv_std_logic_vector(1920, 16),
32784 => conv_std_logic_vector(2048, 16),
32785 => conv_std_logic_vector(2176, 16),
32786 => conv_std_logic_vector(2304, 16),
32787 => conv_std_logic_vector(2432, 16),
32788 => conv_std_logic_vector(2560, 16),
32789 => conv_std_logic_vector(2688, 16),
32790 => conv_std_logic_vector(2816, 16),
32791 => conv_std_logic_vector(2944, 16),
32792 => conv_std_logic_vector(3072, 16),
32793 => conv_std_logic_vector(3200, 16),
32794 => conv_std_logic_vector(3328, 16),
32795 => conv_std_logic_vector(3456, 16),
32796 => conv_std_logic_vector(3584, 16),
32797 => conv_std_logic_vector(3712, 16),
32798 => conv_std_logic_vector(3840, 16),
32799 => conv_std_logic_vector(3968, 16),
32800 => conv_std_logic_vector(4096, 16),
32801 => conv_std_logic_vector(4224, 16),
32802 => conv_std_logic_vector(4352, 16),
32803 => conv_std_logic_vector(4480, 16),
32804 => conv_std_logic_vector(4608, 16),
32805 => conv_std_logic_vector(4736, 16),
32806 => conv_std_logic_vector(4864, 16),
32807 => conv_std_logic_vector(4992, 16),
32808 => conv_std_logic_vector(5120, 16),
32809 => conv_std_logic_vector(5248, 16),
32810 => conv_std_logic_vector(5376, 16),
32811 => conv_std_logic_vector(5504, 16),
32812 => conv_std_logic_vector(5632, 16),
32813 => conv_std_logic_vector(5760, 16),
32814 => conv_std_logic_vector(5888, 16),
32815 => conv_std_logic_vector(6016, 16),
32816 => conv_std_logic_vector(6144, 16),
32817 => conv_std_logic_vector(6272, 16),
32818 => conv_std_logic_vector(6400, 16),
32819 => conv_std_logic_vector(6528, 16),
32820 => conv_std_logic_vector(6656, 16),
32821 => conv_std_logic_vector(6784, 16),
32822 => conv_std_logic_vector(6912, 16),
32823 => conv_std_logic_vector(7040, 16),
32824 => conv_std_logic_vector(7168, 16),
32825 => conv_std_logic_vector(7296, 16),
32826 => conv_std_logic_vector(7424, 16),
32827 => conv_std_logic_vector(7552, 16),
32828 => conv_std_logic_vector(7680, 16),
32829 => conv_std_logic_vector(7808, 16),
32830 => conv_std_logic_vector(7936, 16),
32831 => conv_std_logic_vector(8064, 16),
32832 => conv_std_logic_vector(8192, 16),
32833 => conv_std_logic_vector(8320, 16),
32834 => conv_std_logic_vector(8448, 16),
32835 => conv_std_logic_vector(8576, 16),
32836 => conv_std_logic_vector(8704, 16),
32837 => conv_std_logic_vector(8832, 16),
32838 => conv_std_logic_vector(8960, 16),
32839 => conv_std_logic_vector(9088, 16),
32840 => conv_std_logic_vector(9216, 16),
32841 => conv_std_logic_vector(9344, 16),
32842 => conv_std_logic_vector(9472, 16),
32843 => conv_std_logic_vector(9600, 16),
32844 => conv_std_logic_vector(9728, 16),
32845 => conv_std_logic_vector(9856, 16),
32846 => conv_std_logic_vector(9984, 16),
32847 => conv_std_logic_vector(10112, 16),
32848 => conv_std_logic_vector(10240, 16),
32849 => conv_std_logic_vector(10368, 16),
32850 => conv_std_logic_vector(10496, 16),
32851 => conv_std_logic_vector(10624, 16),
32852 => conv_std_logic_vector(10752, 16),
32853 => conv_std_logic_vector(10880, 16),
32854 => conv_std_logic_vector(11008, 16),
32855 => conv_std_logic_vector(11136, 16),
32856 => conv_std_logic_vector(11264, 16),
32857 => conv_std_logic_vector(11392, 16),
32858 => conv_std_logic_vector(11520, 16),
32859 => conv_std_logic_vector(11648, 16),
32860 => conv_std_logic_vector(11776, 16),
32861 => conv_std_logic_vector(11904, 16),
32862 => conv_std_logic_vector(12032, 16),
32863 => conv_std_logic_vector(12160, 16),
32864 => conv_std_logic_vector(12288, 16),
32865 => conv_std_logic_vector(12416, 16),
32866 => conv_std_logic_vector(12544, 16),
32867 => conv_std_logic_vector(12672, 16),
32868 => conv_std_logic_vector(12800, 16),
32869 => conv_std_logic_vector(12928, 16),
32870 => conv_std_logic_vector(13056, 16),
32871 => conv_std_logic_vector(13184, 16),
32872 => conv_std_logic_vector(13312, 16),
32873 => conv_std_logic_vector(13440, 16),
32874 => conv_std_logic_vector(13568, 16),
32875 => conv_std_logic_vector(13696, 16),
32876 => conv_std_logic_vector(13824, 16),
32877 => conv_std_logic_vector(13952, 16),
32878 => conv_std_logic_vector(14080, 16),
32879 => conv_std_logic_vector(14208, 16),
32880 => conv_std_logic_vector(14336, 16),
32881 => conv_std_logic_vector(14464, 16),
32882 => conv_std_logic_vector(14592, 16),
32883 => conv_std_logic_vector(14720, 16),
32884 => conv_std_logic_vector(14848, 16),
32885 => conv_std_logic_vector(14976, 16),
32886 => conv_std_logic_vector(15104, 16),
32887 => conv_std_logic_vector(15232, 16),
32888 => conv_std_logic_vector(15360, 16),
32889 => conv_std_logic_vector(15488, 16),
32890 => conv_std_logic_vector(15616, 16),
32891 => conv_std_logic_vector(15744, 16),
32892 => conv_std_logic_vector(15872, 16),
32893 => conv_std_logic_vector(16000, 16),
32894 => conv_std_logic_vector(16128, 16),
32895 => conv_std_logic_vector(16256, 16),
32896 => conv_std_logic_vector(16384, 16),
32897 => conv_std_logic_vector(16512, 16),
32898 => conv_std_logic_vector(16640, 16),
32899 => conv_std_logic_vector(16768, 16),
32900 => conv_std_logic_vector(16896, 16),
32901 => conv_std_logic_vector(17024, 16),
32902 => conv_std_logic_vector(17152, 16),
32903 => conv_std_logic_vector(17280, 16),
32904 => conv_std_logic_vector(17408, 16),
32905 => conv_std_logic_vector(17536, 16),
32906 => conv_std_logic_vector(17664, 16),
32907 => conv_std_logic_vector(17792, 16),
32908 => conv_std_logic_vector(17920, 16),
32909 => conv_std_logic_vector(18048, 16),
32910 => conv_std_logic_vector(18176, 16),
32911 => conv_std_logic_vector(18304, 16),
32912 => conv_std_logic_vector(18432, 16),
32913 => conv_std_logic_vector(18560, 16),
32914 => conv_std_logic_vector(18688, 16),
32915 => conv_std_logic_vector(18816, 16),
32916 => conv_std_logic_vector(18944, 16),
32917 => conv_std_logic_vector(19072, 16),
32918 => conv_std_logic_vector(19200, 16),
32919 => conv_std_logic_vector(19328, 16),
32920 => conv_std_logic_vector(19456, 16),
32921 => conv_std_logic_vector(19584, 16),
32922 => conv_std_logic_vector(19712, 16),
32923 => conv_std_logic_vector(19840, 16),
32924 => conv_std_logic_vector(19968, 16),
32925 => conv_std_logic_vector(20096, 16),
32926 => conv_std_logic_vector(20224, 16),
32927 => conv_std_logic_vector(20352, 16),
32928 => conv_std_logic_vector(20480, 16),
32929 => conv_std_logic_vector(20608, 16),
32930 => conv_std_logic_vector(20736, 16),
32931 => conv_std_logic_vector(20864, 16),
32932 => conv_std_logic_vector(20992, 16),
32933 => conv_std_logic_vector(21120, 16),
32934 => conv_std_logic_vector(21248, 16),
32935 => conv_std_logic_vector(21376, 16),
32936 => conv_std_logic_vector(21504, 16),
32937 => conv_std_logic_vector(21632, 16),
32938 => conv_std_logic_vector(21760, 16),
32939 => conv_std_logic_vector(21888, 16),
32940 => conv_std_logic_vector(22016, 16),
32941 => conv_std_logic_vector(22144, 16),
32942 => conv_std_logic_vector(22272, 16),
32943 => conv_std_logic_vector(22400, 16),
32944 => conv_std_logic_vector(22528, 16),
32945 => conv_std_logic_vector(22656, 16),
32946 => conv_std_logic_vector(22784, 16),
32947 => conv_std_logic_vector(22912, 16),
32948 => conv_std_logic_vector(23040, 16),
32949 => conv_std_logic_vector(23168, 16),
32950 => conv_std_logic_vector(23296, 16),
32951 => conv_std_logic_vector(23424, 16),
32952 => conv_std_logic_vector(23552, 16),
32953 => conv_std_logic_vector(23680, 16),
32954 => conv_std_logic_vector(23808, 16),
32955 => conv_std_logic_vector(23936, 16),
32956 => conv_std_logic_vector(24064, 16),
32957 => conv_std_logic_vector(24192, 16),
32958 => conv_std_logic_vector(24320, 16),
32959 => conv_std_logic_vector(24448, 16),
32960 => conv_std_logic_vector(24576, 16),
32961 => conv_std_logic_vector(24704, 16),
32962 => conv_std_logic_vector(24832, 16),
32963 => conv_std_logic_vector(24960, 16),
32964 => conv_std_logic_vector(25088, 16),
32965 => conv_std_logic_vector(25216, 16),
32966 => conv_std_logic_vector(25344, 16),
32967 => conv_std_logic_vector(25472, 16),
32968 => conv_std_logic_vector(25600, 16),
32969 => conv_std_logic_vector(25728, 16),
32970 => conv_std_logic_vector(25856, 16),
32971 => conv_std_logic_vector(25984, 16),
32972 => conv_std_logic_vector(26112, 16),
32973 => conv_std_logic_vector(26240, 16),
32974 => conv_std_logic_vector(26368, 16),
32975 => conv_std_logic_vector(26496, 16),
32976 => conv_std_logic_vector(26624, 16),
32977 => conv_std_logic_vector(26752, 16),
32978 => conv_std_logic_vector(26880, 16),
32979 => conv_std_logic_vector(27008, 16),
32980 => conv_std_logic_vector(27136, 16),
32981 => conv_std_logic_vector(27264, 16),
32982 => conv_std_logic_vector(27392, 16),
32983 => conv_std_logic_vector(27520, 16),
32984 => conv_std_logic_vector(27648, 16),
32985 => conv_std_logic_vector(27776, 16),
32986 => conv_std_logic_vector(27904, 16),
32987 => conv_std_logic_vector(28032, 16),
32988 => conv_std_logic_vector(28160, 16),
32989 => conv_std_logic_vector(28288, 16),
32990 => conv_std_logic_vector(28416, 16),
32991 => conv_std_logic_vector(28544, 16),
32992 => conv_std_logic_vector(28672, 16),
32993 => conv_std_logic_vector(28800, 16),
32994 => conv_std_logic_vector(28928, 16),
32995 => conv_std_logic_vector(29056, 16),
32996 => conv_std_logic_vector(29184, 16),
32997 => conv_std_logic_vector(29312, 16),
32998 => conv_std_logic_vector(29440, 16),
32999 => conv_std_logic_vector(29568, 16),
33000 => conv_std_logic_vector(29696, 16),
33001 => conv_std_logic_vector(29824, 16),
33002 => conv_std_logic_vector(29952, 16),
33003 => conv_std_logic_vector(30080, 16),
33004 => conv_std_logic_vector(30208, 16),
33005 => conv_std_logic_vector(30336, 16),
33006 => conv_std_logic_vector(30464, 16),
33007 => conv_std_logic_vector(30592, 16),
33008 => conv_std_logic_vector(30720, 16),
33009 => conv_std_logic_vector(30848, 16),
33010 => conv_std_logic_vector(30976, 16),
33011 => conv_std_logic_vector(31104, 16),
33012 => conv_std_logic_vector(31232, 16),
33013 => conv_std_logic_vector(31360, 16),
33014 => conv_std_logic_vector(31488, 16),
33015 => conv_std_logic_vector(31616, 16),
33016 => conv_std_logic_vector(31744, 16),
33017 => conv_std_logic_vector(31872, 16),
33018 => conv_std_logic_vector(32000, 16),
33019 => conv_std_logic_vector(32128, 16),
33020 => conv_std_logic_vector(32256, 16),
33021 => conv_std_logic_vector(32384, 16),
33022 => conv_std_logic_vector(32512, 16),
33023 => conv_std_logic_vector(32640, 16),
33024 => conv_std_logic_vector(0, 16),
33025 => conv_std_logic_vector(129, 16),
33026 => conv_std_logic_vector(258, 16),
33027 => conv_std_logic_vector(387, 16),
33028 => conv_std_logic_vector(516, 16),
33029 => conv_std_logic_vector(645, 16),
33030 => conv_std_logic_vector(774, 16),
33031 => conv_std_logic_vector(903, 16),
33032 => conv_std_logic_vector(1032, 16),
33033 => conv_std_logic_vector(1161, 16),
33034 => conv_std_logic_vector(1290, 16),
33035 => conv_std_logic_vector(1419, 16),
33036 => conv_std_logic_vector(1548, 16),
33037 => conv_std_logic_vector(1677, 16),
33038 => conv_std_logic_vector(1806, 16),
33039 => conv_std_logic_vector(1935, 16),
33040 => conv_std_logic_vector(2064, 16),
33041 => conv_std_logic_vector(2193, 16),
33042 => conv_std_logic_vector(2322, 16),
33043 => conv_std_logic_vector(2451, 16),
33044 => conv_std_logic_vector(2580, 16),
33045 => conv_std_logic_vector(2709, 16),
33046 => conv_std_logic_vector(2838, 16),
33047 => conv_std_logic_vector(2967, 16),
33048 => conv_std_logic_vector(3096, 16),
33049 => conv_std_logic_vector(3225, 16),
33050 => conv_std_logic_vector(3354, 16),
33051 => conv_std_logic_vector(3483, 16),
33052 => conv_std_logic_vector(3612, 16),
33053 => conv_std_logic_vector(3741, 16),
33054 => conv_std_logic_vector(3870, 16),
33055 => conv_std_logic_vector(3999, 16),
33056 => conv_std_logic_vector(4128, 16),
33057 => conv_std_logic_vector(4257, 16),
33058 => conv_std_logic_vector(4386, 16),
33059 => conv_std_logic_vector(4515, 16),
33060 => conv_std_logic_vector(4644, 16),
33061 => conv_std_logic_vector(4773, 16),
33062 => conv_std_logic_vector(4902, 16),
33063 => conv_std_logic_vector(5031, 16),
33064 => conv_std_logic_vector(5160, 16),
33065 => conv_std_logic_vector(5289, 16),
33066 => conv_std_logic_vector(5418, 16),
33067 => conv_std_logic_vector(5547, 16),
33068 => conv_std_logic_vector(5676, 16),
33069 => conv_std_logic_vector(5805, 16),
33070 => conv_std_logic_vector(5934, 16),
33071 => conv_std_logic_vector(6063, 16),
33072 => conv_std_logic_vector(6192, 16),
33073 => conv_std_logic_vector(6321, 16),
33074 => conv_std_logic_vector(6450, 16),
33075 => conv_std_logic_vector(6579, 16),
33076 => conv_std_logic_vector(6708, 16),
33077 => conv_std_logic_vector(6837, 16),
33078 => conv_std_logic_vector(6966, 16),
33079 => conv_std_logic_vector(7095, 16),
33080 => conv_std_logic_vector(7224, 16),
33081 => conv_std_logic_vector(7353, 16),
33082 => conv_std_logic_vector(7482, 16),
33083 => conv_std_logic_vector(7611, 16),
33084 => conv_std_logic_vector(7740, 16),
33085 => conv_std_logic_vector(7869, 16),
33086 => conv_std_logic_vector(7998, 16),
33087 => conv_std_logic_vector(8127, 16),
33088 => conv_std_logic_vector(8256, 16),
33089 => conv_std_logic_vector(8385, 16),
33090 => conv_std_logic_vector(8514, 16),
33091 => conv_std_logic_vector(8643, 16),
33092 => conv_std_logic_vector(8772, 16),
33093 => conv_std_logic_vector(8901, 16),
33094 => conv_std_logic_vector(9030, 16),
33095 => conv_std_logic_vector(9159, 16),
33096 => conv_std_logic_vector(9288, 16),
33097 => conv_std_logic_vector(9417, 16),
33098 => conv_std_logic_vector(9546, 16),
33099 => conv_std_logic_vector(9675, 16),
33100 => conv_std_logic_vector(9804, 16),
33101 => conv_std_logic_vector(9933, 16),
33102 => conv_std_logic_vector(10062, 16),
33103 => conv_std_logic_vector(10191, 16),
33104 => conv_std_logic_vector(10320, 16),
33105 => conv_std_logic_vector(10449, 16),
33106 => conv_std_logic_vector(10578, 16),
33107 => conv_std_logic_vector(10707, 16),
33108 => conv_std_logic_vector(10836, 16),
33109 => conv_std_logic_vector(10965, 16),
33110 => conv_std_logic_vector(11094, 16),
33111 => conv_std_logic_vector(11223, 16),
33112 => conv_std_logic_vector(11352, 16),
33113 => conv_std_logic_vector(11481, 16),
33114 => conv_std_logic_vector(11610, 16),
33115 => conv_std_logic_vector(11739, 16),
33116 => conv_std_logic_vector(11868, 16),
33117 => conv_std_logic_vector(11997, 16),
33118 => conv_std_logic_vector(12126, 16),
33119 => conv_std_logic_vector(12255, 16),
33120 => conv_std_logic_vector(12384, 16),
33121 => conv_std_logic_vector(12513, 16),
33122 => conv_std_logic_vector(12642, 16),
33123 => conv_std_logic_vector(12771, 16),
33124 => conv_std_logic_vector(12900, 16),
33125 => conv_std_logic_vector(13029, 16),
33126 => conv_std_logic_vector(13158, 16),
33127 => conv_std_logic_vector(13287, 16),
33128 => conv_std_logic_vector(13416, 16),
33129 => conv_std_logic_vector(13545, 16),
33130 => conv_std_logic_vector(13674, 16),
33131 => conv_std_logic_vector(13803, 16),
33132 => conv_std_logic_vector(13932, 16),
33133 => conv_std_logic_vector(14061, 16),
33134 => conv_std_logic_vector(14190, 16),
33135 => conv_std_logic_vector(14319, 16),
33136 => conv_std_logic_vector(14448, 16),
33137 => conv_std_logic_vector(14577, 16),
33138 => conv_std_logic_vector(14706, 16),
33139 => conv_std_logic_vector(14835, 16),
33140 => conv_std_logic_vector(14964, 16),
33141 => conv_std_logic_vector(15093, 16),
33142 => conv_std_logic_vector(15222, 16),
33143 => conv_std_logic_vector(15351, 16),
33144 => conv_std_logic_vector(15480, 16),
33145 => conv_std_logic_vector(15609, 16),
33146 => conv_std_logic_vector(15738, 16),
33147 => conv_std_logic_vector(15867, 16),
33148 => conv_std_logic_vector(15996, 16),
33149 => conv_std_logic_vector(16125, 16),
33150 => conv_std_logic_vector(16254, 16),
33151 => conv_std_logic_vector(16383, 16),
33152 => conv_std_logic_vector(16512, 16),
33153 => conv_std_logic_vector(16641, 16),
33154 => conv_std_logic_vector(16770, 16),
33155 => conv_std_logic_vector(16899, 16),
33156 => conv_std_logic_vector(17028, 16),
33157 => conv_std_logic_vector(17157, 16),
33158 => conv_std_logic_vector(17286, 16),
33159 => conv_std_logic_vector(17415, 16),
33160 => conv_std_logic_vector(17544, 16),
33161 => conv_std_logic_vector(17673, 16),
33162 => conv_std_logic_vector(17802, 16),
33163 => conv_std_logic_vector(17931, 16),
33164 => conv_std_logic_vector(18060, 16),
33165 => conv_std_logic_vector(18189, 16),
33166 => conv_std_logic_vector(18318, 16),
33167 => conv_std_logic_vector(18447, 16),
33168 => conv_std_logic_vector(18576, 16),
33169 => conv_std_logic_vector(18705, 16),
33170 => conv_std_logic_vector(18834, 16),
33171 => conv_std_logic_vector(18963, 16),
33172 => conv_std_logic_vector(19092, 16),
33173 => conv_std_logic_vector(19221, 16),
33174 => conv_std_logic_vector(19350, 16),
33175 => conv_std_logic_vector(19479, 16),
33176 => conv_std_logic_vector(19608, 16),
33177 => conv_std_logic_vector(19737, 16),
33178 => conv_std_logic_vector(19866, 16),
33179 => conv_std_logic_vector(19995, 16),
33180 => conv_std_logic_vector(20124, 16),
33181 => conv_std_logic_vector(20253, 16),
33182 => conv_std_logic_vector(20382, 16),
33183 => conv_std_logic_vector(20511, 16),
33184 => conv_std_logic_vector(20640, 16),
33185 => conv_std_logic_vector(20769, 16),
33186 => conv_std_logic_vector(20898, 16),
33187 => conv_std_logic_vector(21027, 16),
33188 => conv_std_logic_vector(21156, 16),
33189 => conv_std_logic_vector(21285, 16),
33190 => conv_std_logic_vector(21414, 16),
33191 => conv_std_logic_vector(21543, 16),
33192 => conv_std_logic_vector(21672, 16),
33193 => conv_std_logic_vector(21801, 16),
33194 => conv_std_logic_vector(21930, 16),
33195 => conv_std_logic_vector(22059, 16),
33196 => conv_std_logic_vector(22188, 16),
33197 => conv_std_logic_vector(22317, 16),
33198 => conv_std_logic_vector(22446, 16),
33199 => conv_std_logic_vector(22575, 16),
33200 => conv_std_logic_vector(22704, 16),
33201 => conv_std_logic_vector(22833, 16),
33202 => conv_std_logic_vector(22962, 16),
33203 => conv_std_logic_vector(23091, 16),
33204 => conv_std_logic_vector(23220, 16),
33205 => conv_std_logic_vector(23349, 16),
33206 => conv_std_logic_vector(23478, 16),
33207 => conv_std_logic_vector(23607, 16),
33208 => conv_std_logic_vector(23736, 16),
33209 => conv_std_logic_vector(23865, 16),
33210 => conv_std_logic_vector(23994, 16),
33211 => conv_std_logic_vector(24123, 16),
33212 => conv_std_logic_vector(24252, 16),
33213 => conv_std_logic_vector(24381, 16),
33214 => conv_std_logic_vector(24510, 16),
33215 => conv_std_logic_vector(24639, 16),
33216 => conv_std_logic_vector(24768, 16),
33217 => conv_std_logic_vector(24897, 16),
33218 => conv_std_logic_vector(25026, 16),
33219 => conv_std_logic_vector(25155, 16),
33220 => conv_std_logic_vector(25284, 16),
33221 => conv_std_logic_vector(25413, 16),
33222 => conv_std_logic_vector(25542, 16),
33223 => conv_std_logic_vector(25671, 16),
33224 => conv_std_logic_vector(25800, 16),
33225 => conv_std_logic_vector(25929, 16),
33226 => conv_std_logic_vector(26058, 16),
33227 => conv_std_logic_vector(26187, 16),
33228 => conv_std_logic_vector(26316, 16),
33229 => conv_std_logic_vector(26445, 16),
33230 => conv_std_logic_vector(26574, 16),
33231 => conv_std_logic_vector(26703, 16),
33232 => conv_std_logic_vector(26832, 16),
33233 => conv_std_logic_vector(26961, 16),
33234 => conv_std_logic_vector(27090, 16),
33235 => conv_std_logic_vector(27219, 16),
33236 => conv_std_logic_vector(27348, 16),
33237 => conv_std_logic_vector(27477, 16),
33238 => conv_std_logic_vector(27606, 16),
33239 => conv_std_logic_vector(27735, 16),
33240 => conv_std_logic_vector(27864, 16),
33241 => conv_std_logic_vector(27993, 16),
33242 => conv_std_logic_vector(28122, 16),
33243 => conv_std_logic_vector(28251, 16),
33244 => conv_std_logic_vector(28380, 16),
33245 => conv_std_logic_vector(28509, 16),
33246 => conv_std_logic_vector(28638, 16),
33247 => conv_std_logic_vector(28767, 16),
33248 => conv_std_logic_vector(28896, 16),
33249 => conv_std_logic_vector(29025, 16),
33250 => conv_std_logic_vector(29154, 16),
33251 => conv_std_logic_vector(29283, 16),
33252 => conv_std_logic_vector(29412, 16),
33253 => conv_std_logic_vector(29541, 16),
33254 => conv_std_logic_vector(29670, 16),
33255 => conv_std_logic_vector(29799, 16),
33256 => conv_std_logic_vector(29928, 16),
33257 => conv_std_logic_vector(30057, 16),
33258 => conv_std_logic_vector(30186, 16),
33259 => conv_std_logic_vector(30315, 16),
33260 => conv_std_logic_vector(30444, 16),
33261 => conv_std_logic_vector(30573, 16),
33262 => conv_std_logic_vector(30702, 16),
33263 => conv_std_logic_vector(30831, 16),
33264 => conv_std_logic_vector(30960, 16),
33265 => conv_std_logic_vector(31089, 16),
33266 => conv_std_logic_vector(31218, 16),
33267 => conv_std_logic_vector(31347, 16),
33268 => conv_std_logic_vector(31476, 16),
33269 => conv_std_logic_vector(31605, 16),
33270 => conv_std_logic_vector(31734, 16),
33271 => conv_std_logic_vector(31863, 16),
33272 => conv_std_logic_vector(31992, 16),
33273 => conv_std_logic_vector(32121, 16),
33274 => conv_std_logic_vector(32250, 16),
33275 => conv_std_logic_vector(32379, 16),
33276 => conv_std_logic_vector(32508, 16),
33277 => conv_std_logic_vector(32637, 16),
33278 => conv_std_logic_vector(32766, 16),
33279 => conv_std_logic_vector(32895, 16),
33280 => conv_std_logic_vector(0, 16),
33281 => conv_std_logic_vector(130, 16),
33282 => conv_std_logic_vector(260, 16),
33283 => conv_std_logic_vector(390, 16),
33284 => conv_std_logic_vector(520, 16),
33285 => conv_std_logic_vector(650, 16),
33286 => conv_std_logic_vector(780, 16),
33287 => conv_std_logic_vector(910, 16),
33288 => conv_std_logic_vector(1040, 16),
33289 => conv_std_logic_vector(1170, 16),
33290 => conv_std_logic_vector(1300, 16),
33291 => conv_std_logic_vector(1430, 16),
33292 => conv_std_logic_vector(1560, 16),
33293 => conv_std_logic_vector(1690, 16),
33294 => conv_std_logic_vector(1820, 16),
33295 => conv_std_logic_vector(1950, 16),
33296 => conv_std_logic_vector(2080, 16),
33297 => conv_std_logic_vector(2210, 16),
33298 => conv_std_logic_vector(2340, 16),
33299 => conv_std_logic_vector(2470, 16),
33300 => conv_std_logic_vector(2600, 16),
33301 => conv_std_logic_vector(2730, 16),
33302 => conv_std_logic_vector(2860, 16),
33303 => conv_std_logic_vector(2990, 16),
33304 => conv_std_logic_vector(3120, 16),
33305 => conv_std_logic_vector(3250, 16),
33306 => conv_std_logic_vector(3380, 16),
33307 => conv_std_logic_vector(3510, 16),
33308 => conv_std_logic_vector(3640, 16),
33309 => conv_std_logic_vector(3770, 16),
33310 => conv_std_logic_vector(3900, 16),
33311 => conv_std_logic_vector(4030, 16),
33312 => conv_std_logic_vector(4160, 16),
33313 => conv_std_logic_vector(4290, 16),
33314 => conv_std_logic_vector(4420, 16),
33315 => conv_std_logic_vector(4550, 16),
33316 => conv_std_logic_vector(4680, 16),
33317 => conv_std_logic_vector(4810, 16),
33318 => conv_std_logic_vector(4940, 16),
33319 => conv_std_logic_vector(5070, 16),
33320 => conv_std_logic_vector(5200, 16),
33321 => conv_std_logic_vector(5330, 16),
33322 => conv_std_logic_vector(5460, 16),
33323 => conv_std_logic_vector(5590, 16),
33324 => conv_std_logic_vector(5720, 16),
33325 => conv_std_logic_vector(5850, 16),
33326 => conv_std_logic_vector(5980, 16),
33327 => conv_std_logic_vector(6110, 16),
33328 => conv_std_logic_vector(6240, 16),
33329 => conv_std_logic_vector(6370, 16),
33330 => conv_std_logic_vector(6500, 16),
33331 => conv_std_logic_vector(6630, 16),
33332 => conv_std_logic_vector(6760, 16),
33333 => conv_std_logic_vector(6890, 16),
33334 => conv_std_logic_vector(7020, 16),
33335 => conv_std_logic_vector(7150, 16),
33336 => conv_std_logic_vector(7280, 16),
33337 => conv_std_logic_vector(7410, 16),
33338 => conv_std_logic_vector(7540, 16),
33339 => conv_std_logic_vector(7670, 16),
33340 => conv_std_logic_vector(7800, 16),
33341 => conv_std_logic_vector(7930, 16),
33342 => conv_std_logic_vector(8060, 16),
33343 => conv_std_logic_vector(8190, 16),
33344 => conv_std_logic_vector(8320, 16),
33345 => conv_std_logic_vector(8450, 16),
33346 => conv_std_logic_vector(8580, 16),
33347 => conv_std_logic_vector(8710, 16),
33348 => conv_std_logic_vector(8840, 16),
33349 => conv_std_logic_vector(8970, 16),
33350 => conv_std_logic_vector(9100, 16),
33351 => conv_std_logic_vector(9230, 16),
33352 => conv_std_logic_vector(9360, 16),
33353 => conv_std_logic_vector(9490, 16),
33354 => conv_std_logic_vector(9620, 16),
33355 => conv_std_logic_vector(9750, 16),
33356 => conv_std_logic_vector(9880, 16),
33357 => conv_std_logic_vector(10010, 16),
33358 => conv_std_logic_vector(10140, 16),
33359 => conv_std_logic_vector(10270, 16),
33360 => conv_std_logic_vector(10400, 16),
33361 => conv_std_logic_vector(10530, 16),
33362 => conv_std_logic_vector(10660, 16),
33363 => conv_std_logic_vector(10790, 16),
33364 => conv_std_logic_vector(10920, 16),
33365 => conv_std_logic_vector(11050, 16),
33366 => conv_std_logic_vector(11180, 16),
33367 => conv_std_logic_vector(11310, 16),
33368 => conv_std_logic_vector(11440, 16),
33369 => conv_std_logic_vector(11570, 16),
33370 => conv_std_logic_vector(11700, 16),
33371 => conv_std_logic_vector(11830, 16),
33372 => conv_std_logic_vector(11960, 16),
33373 => conv_std_logic_vector(12090, 16),
33374 => conv_std_logic_vector(12220, 16),
33375 => conv_std_logic_vector(12350, 16),
33376 => conv_std_logic_vector(12480, 16),
33377 => conv_std_logic_vector(12610, 16),
33378 => conv_std_logic_vector(12740, 16),
33379 => conv_std_logic_vector(12870, 16),
33380 => conv_std_logic_vector(13000, 16),
33381 => conv_std_logic_vector(13130, 16),
33382 => conv_std_logic_vector(13260, 16),
33383 => conv_std_logic_vector(13390, 16),
33384 => conv_std_logic_vector(13520, 16),
33385 => conv_std_logic_vector(13650, 16),
33386 => conv_std_logic_vector(13780, 16),
33387 => conv_std_logic_vector(13910, 16),
33388 => conv_std_logic_vector(14040, 16),
33389 => conv_std_logic_vector(14170, 16),
33390 => conv_std_logic_vector(14300, 16),
33391 => conv_std_logic_vector(14430, 16),
33392 => conv_std_logic_vector(14560, 16),
33393 => conv_std_logic_vector(14690, 16),
33394 => conv_std_logic_vector(14820, 16),
33395 => conv_std_logic_vector(14950, 16),
33396 => conv_std_logic_vector(15080, 16),
33397 => conv_std_logic_vector(15210, 16),
33398 => conv_std_logic_vector(15340, 16),
33399 => conv_std_logic_vector(15470, 16),
33400 => conv_std_logic_vector(15600, 16),
33401 => conv_std_logic_vector(15730, 16),
33402 => conv_std_logic_vector(15860, 16),
33403 => conv_std_logic_vector(15990, 16),
33404 => conv_std_logic_vector(16120, 16),
33405 => conv_std_logic_vector(16250, 16),
33406 => conv_std_logic_vector(16380, 16),
33407 => conv_std_logic_vector(16510, 16),
33408 => conv_std_logic_vector(16640, 16),
33409 => conv_std_logic_vector(16770, 16),
33410 => conv_std_logic_vector(16900, 16),
33411 => conv_std_logic_vector(17030, 16),
33412 => conv_std_logic_vector(17160, 16),
33413 => conv_std_logic_vector(17290, 16),
33414 => conv_std_logic_vector(17420, 16),
33415 => conv_std_logic_vector(17550, 16),
33416 => conv_std_logic_vector(17680, 16),
33417 => conv_std_logic_vector(17810, 16),
33418 => conv_std_logic_vector(17940, 16),
33419 => conv_std_logic_vector(18070, 16),
33420 => conv_std_logic_vector(18200, 16),
33421 => conv_std_logic_vector(18330, 16),
33422 => conv_std_logic_vector(18460, 16),
33423 => conv_std_logic_vector(18590, 16),
33424 => conv_std_logic_vector(18720, 16),
33425 => conv_std_logic_vector(18850, 16),
33426 => conv_std_logic_vector(18980, 16),
33427 => conv_std_logic_vector(19110, 16),
33428 => conv_std_logic_vector(19240, 16),
33429 => conv_std_logic_vector(19370, 16),
33430 => conv_std_logic_vector(19500, 16),
33431 => conv_std_logic_vector(19630, 16),
33432 => conv_std_logic_vector(19760, 16),
33433 => conv_std_logic_vector(19890, 16),
33434 => conv_std_logic_vector(20020, 16),
33435 => conv_std_logic_vector(20150, 16),
33436 => conv_std_logic_vector(20280, 16),
33437 => conv_std_logic_vector(20410, 16),
33438 => conv_std_logic_vector(20540, 16),
33439 => conv_std_logic_vector(20670, 16),
33440 => conv_std_logic_vector(20800, 16),
33441 => conv_std_logic_vector(20930, 16),
33442 => conv_std_logic_vector(21060, 16),
33443 => conv_std_logic_vector(21190, 16),
33444 => conv_std_logic_vector(21320, 16),
33445 => conv_std_logic_vector(21450, 16),
33446 => conv_std_logic_vector(21580, 16),
33447 => conv_std_logic_vector(21710, 16),
33448 => conv_std_logic_vector(21840, 16),
33449 => conv_std_logic_vector(21970, 16),
33450 => conv_std_logic_vector(22100, 16),
33451 => conv_std_logic_vector(22230, 16),
33452 => conv_std_logic_vector(22360, 16),
33453 => conv_std_logic_vector(22490, 16),
33454 => conv_std_logic_vector(22620, 16),
33455 => conv_std_logic_vector(22750, 16),
33456 => conv_std_logic_vector(22880, 16),
33457 => conv_std_logic_vector(23010, 16),
33458 => conv_std_logic_vector(23140, 16),
33459 => conv_std_logic_vector(23270, 16),
33460 => conv_std_logic_vector(23400, 16),
33461 => conv_std_logic_vector(23530, 16),
33462 => conv_std_logic_vector(23660, 16),
33463 => conv_std_logic_vector(23790, 16),
33464 => conv_std_logic_vector(23920, 16),
33465 => conv_std_logic_vector(24050, 16),
33466 => conv_std_logic_vector(24180, 16),
33467 => conv_std_logic_vector(24310, 16),
33468 => conv_std_logic_vector(24440, 16),
33469 => conv_std_logic_vector(24570, 16),
33470 => conv_std_logic_vector(24700, 16),
33471 => conv_std_logic_vector(24830, 16),
33472 => conv_std_logic_vector(24960, 16),
33473 => conv_std_logic_vector(25090, 16),
33474 => conv_std_logic_vector(25220, 16),
33475 => conv_std_logic_vector(25350, 16),
33476 => conv_std_logic_vector(25480, 16),
33477 => conv_std_logic_vector(25610, 16),
33478 => conv_std_logic_vector(25740, 16),
33479 => conv_std_logic_vector(25870, 16),
33480 => conv_std_logic_vector(26000, 16),
33481 => conv_std_logic_vector(26130, 16),
33482 => conv_std_logic_vector(26260, 16),
33483 => conv_std_logic_vector(26390, 16),
33484 => conv_std_logic_vector(26520, 16),
33485 => conv_std_logic_vector(26650, 16),
33486 => conv_std_logic_vector(26780, 16),
33487 => conv_std_logic_vector(26910, 16),
33488 => conv_std_logic_vector(27040, 16),
33489 => conv_std_logic_vector(27170, 16),
33490 => conv_std_logic_vector(27300, 16),
33491 => conv_std_logic_vector(27430, 16),
33492 => conv_std_logic_vector(27560, 16),
33493 => conv_std_logic_vector(27690, 16),
33494 => conv_std_logic_vector(27820, 16),
33495 => conv_std_logic_vector(27950, 16),
33496 => conv_std_logic_vector(28080, 16),
33497 => conv_std_logic_vector(28210, 16),
33498 => conv_std_logic_vector(28340, 16),
33499 => conv_std_logic_vector(28470, 16),
33500 => conv_std_logic_vector(28600, 16),
33501 => conv_std_logic_vector(28730, 16),
33502 => conv_std_logic_vector(28860, 16),
33503 => conv_std_logic_vector(28990, 16),
33504 => conv_std_logic_vector(29120, 16),
33505 => conv_std_logic_vector(29250, 16),
33506 => conv_std_logic_vector(29380, 16),
33507 => conv_std_logic_vector(29510, 16),
33508 => conv_std_logic_vector(29640, 16),
33509 => conv_std_logic_vector(29770, 16),
33510 => conv_std_logic_vector(29900, 16),
33511 => conv_std_logic_vector(30030, 16),
33512 => conv_std_logic_vector(30160, 16),
33513 => conv_std_logic_vector(30290, 16),
33514 => conv_std_logic_vector(30420, 16),
33515 => conv_std_logic_vector(30550, 16),
33516 => conv_std_logic_vector(30680, 16),
33517 => conv_std_logic_vector(30810, 16),
33518 => conv_std_logic_vector(30940, 16),
33519 => conv_std_logic_vector(31070, 16),
33520 => conv_std_logic_vector(31200, 16),
33521 => conv_std_logic_vector(31330, 16),
33522 => conv_std_logic_vector(31460, 16),
33523 => conv_std_logic_vector(31590, 16),
33524 => conv_std_logic_vector(31720, 16),
33525 => conv_std_logic_vector(31850, 16),
33526 => conv_std_logic_vector(31980, 16),
33527 => conv_std_logic_vector(32110, 16),
33528 => conv_std_logic_vector(32240, 16),
33529 => conv_std_logic_vector(32370, 16),
33530 => conv_std_logic_vector(32500, 16),
33531 => conv_std_logic_vector(32630, 16),
33532 => conv_std_logic_vector(32760, 16),
33533 => conv_std_logic_vector(32890, 16),
33534 => conv_std_logic_vector(33020, 16),
33535 => conv_std_logic_vector(33150, 16),
33536 => conv_std_logic_vector(0, 16),
33537 => conv_std_logic_vector(131, 16),
33538 => conv_std_logic_vector(262, 16),
33539 => conv_std_logic_vector(393, 16),
33540 => conv_std_logic_vector(524, 16),
33541 => conv_std_logic_vector(655, 16),
33542 => conv_std_logic_vector(786, 16),
33543 => conv_std_logic_vector(917, 16),
33544 => conv_std_logic_vector(1048, 16),
33545 => conv_std_logic_vector(1179, 16),
33546 => conv_std_logic_vector(1310, 16),
33547 => conv_std_logic_vector(1441, 16),
33548 => conv_std_logic_vector(1572, 16),
33549 => conv_std_logic_vector(1703, 16),
33550 => conv_std_logic_vector(1834, 16),
33551 => conv_std_logic_vector(1965, 16),
33552 => conv_std_logic_vector(2096, 16),
33553 => conv_std_logic_vector(2227, 16),
33554 => conv_std_logic_vector(2358, 16),
33555 => conv_std_logic_vector(2489, 16),
33556 => conv_std_logic_vector(2620, 16),
33557 => conv_std_logic_vector(2751, 16),
33558 => conv_std_logic_vector(2882, 16),
33559 => conv_std_logic_vector(3013, 16),
33560 => conv_std_logic_vector(3144, 16),
33561 => conv_std_logic_vector(3275, 16),
33562 => conv_std_logic_vector(3406, 16),
33563 => conv_std_logic_vector(3537, 16),
33564 => conv_std_logic_vector(3668, 16),
33565 => conv_std_logic_vector(3799, 16),
33566 => conv_std_logic_vector(3930, 16),
33567 => conv_std_logic_vector(4061, 16),
33568 => conv_std_logic_vector(4192, 16),
33569 => conv_std_logic_vector(4323, 16),
33570 => conv_std_logic_vector(4454, 16),
33571 => conv_std_logic_vector(4585, 16),
33572 => conv_std_logic_vector(4716, 16),
33573 => conv_std_logic_vector(4847, 16),
33574 => conv_std_logic_vector(4978, 16),
33575 => conv_std_logic_vector(5109, 16),
33576 => conv_std_logic_vector(5240, 16),
33577 => conv_std_logic_vector(5371, 16),
33578 => conv_std_logic_vector(5502, 16),
33579 => conv_std_logic_vector(5633, 16),
33580 => conv_std_logic_vector(5764, 16),
33581 => conv_std_logic_vector(5895, 16),
33582 => conv_std_logic_vector(6026, 16),
33583 => conv_std_logic_vector(6157, 16),
33584 => conv_std_logic_vector(6288, 16),
33585 => conv_std_logic_vector(6419, 16),
33586 => conv_std_logic_vector(6550, 16),
33587 => conv_std_logic_vector(6681, 16),
33588 => conv_std_logic_vector(6812, 16),
33589 => conv_std_logic_vector(6943, 16),
33590 => conv_std_logic_vector(7074, 16),
33591 => conv_std_logic_vector(7205, 16),
33592 => conv_std_logic_vector(7336, 16),
33593 => conv_std_logic_vector(7467, 16),
33594 => conv_std_logic_vector(7598, 16),
33595 => conv_std_logic_vector(7729, 16),
33596 => conv_std_logic_vector(7860, 16),
33597 => conv_std_logic_vector(7991, 16),
33598 => conv_std_logic_vector(8122, 16),
33599 => conv_std_logic_vector(8253, 16),
33600 => conv_std_logic_vector(8384, 16),
33601 => conv_std_logic_vector(8515, 16),
33602 => conv_std_logic_vector(8646, 16),
33603 => conv_std_logic_vector(8777, 16),
33604 => conv_std_logic_vector(8908, 16),
33605 => conv_std_logic_vector(9039, 16),
33606 => conv_std_logic_vector(9170, 16),
33607 => conv_std_logic_vector(9301, 16),
33608 => conv_std_logic_vector(9432, 16),
33609 => conv_std_logic_vector(9563, 16),
33610 => conv_std_logic_vector(9694, 16),
33611 => conv_std_logic_vector(9825, 16),
33612 => conv_std_logic_vector(9956, 16),
33613 => conv_std_logic_vector(10087, 16),
33614 => conv_std_logic_vector(10218, 16),
33615 => conv_std_logic_vector(10349, 16),
33616 => conv_std_logic_vector(10480, 16),
33617 => conv_std_logic_vector(10611, 16),
33618 => conv_std_logic_vector(10742, 16),
33619 => conv_std_logic_vector(10873, 16),
33620 => conv_std_logic_vector(11004, 16),
33621 => conv_std_logic_vector(11135, 16),
33622 => conv_std_logic_vector(11266, 16),
33623 => conv_std_logic_vector(11397, 16),
33624 => conv_std_logic_vector(11528, 16),
33625 => conv_std_logic_vector(11659, 16),
33626 => conv_std_logic_vector(11790, 16),
33627 => conv_std_logic_vector(11921, 16),
33628 => conv_std_logic_vector(12052, 16),
33629 => conv_std_logic_vector(12183, 16),
33630 => conv_std_logic_vector(12314, 16),
33631 => conv_std_logic_vector(12445, 16),
33632 => conv_std_logic_vector(12576, 16),
33633 => conv_std_logic_vector(12707, 16),
33634 => conv_std_logic_vector(12838, 16),
33635 => conv_std_logic_vector(12969, 16),
33636 => conv_std_logic_vector(13100, 16),
33637 => conv_std_logic_vector(13231, 16),
33638 => conv_std_logic_vector(13362, 16),
33639 => conv_std_logic_vector(13493, 16),
33640 => conv_std_logic_vector(13624, 16),
33641 => conv_std_logic_vector(13755, 16),
33642 => conv_std_logic_vector(13886, 16),
33643 => conv_std_logic_vector(14017, 16),
33644 => conv_std_logic_vector(14148, 16),
33645 => conv_std_logic_vector(14279, 16),
33646 => conv_std_logic_vector(14410, 16),
33647 => conv_std_logic_vector(14541, 16),
33648 => conv_std_logic_vector(14672, 16),
33649 => conv_std_logic_vector(14803, 16),
33650 => conv_std_logic_vector(14934, 16),
33651 => conv_std_logic_vector(15065, 16),
33652 => conv_std_logic_vector(15196, 16),
33653 => conv_std_logic_vector(15327, 16),
33654 => conv_std_logic_vector(15458, 16),
33655 => conv_std_logic_vector(15589, 16),
33656 => conv_std_logic_vector(15720, 16),
33657 => conv_std_logic_vector(15851, 16),
33658 => conv_std_logic_vector(15982, 16),
33659 => conv_std_logic_vector(16113, 16),
33660 => conv_std_logic_vector(16244, 16),
33661 => conv_std_logic_vector(16375, 16),
33662 => conv_std_logic_vector(16506, 16),
33663 => conv_std_logic_vector(16637, 16),
33664 => conv_std_logic_vector(16768, 16),
33665 => conv_std_logic_vector(16899, 16),
33666 => conv_std_logic_vector(17030, 16),
33667 => conv_std_logic_vector(17161, 16),
33668 => conv_std_logic_vector(17292, 16),
33669 => conv_std_logic_vector(17423, 16),
33670 => conv_std_logic_vector(17554, 16),
33671 => conv_std_logic_vector(17685, 16),
33672 => conv_std_logic_vector(17816, 16),
33673 => conv_std_logic_vector(17947, 16),
33674 => conv_std_logic_vector(18078, 16),
33675 => conv_std_logic_vector(18209, 16),
33676 => conv_std_logic_vector(18340, 16),
33677 => conv_std_logic_vector(18471, 16),
33678 => conv_std_logic_vector(18602, 16),
33679 => conv_std_logic_vector(18733, 16),
33680 => conv_std_logic_vector(18864, 16),
33681 => conv_std_logic_vector(18995, 16),
33682 => conv_std_logic_vector(19126, 16),
33683 => conv_std_logic_vector(19257, 16),
33684 => conv_std_logic_vector(19388, 16),
33685 => conv_std_logic_vector(19519, 16),
33686 => conv_std_logic_vector(19650, 16),
33687 => conv_std_logic_vector(19781, 16),
33688 => conv_std_logic_vector(19912, 16),
33689 => conv_std_logic_vector(20043, 16),
33690 => conv_std_logic_vector(20174, 16),
33691 => conv_std_logic_vector(20305, 16),
33692 => conv_std_logic_vector(20436, 16),
33693 => conv_std_logic_vector(20567, 16),
33694 => conv_std_logic_vector(20698, 16),
33695 => conv_std_logic_vector(20829, 16),
33696 => conv_std_logic_vector(20960, 16),
33697 => conv_std_logic_vector(21091, 16),
33698 => conv_std_logic_vector(21222, 16),
33699 => conv_std_logic_vector(21353, 16),
33700 => conv_std_logic_vector(21484, 16),
33701 => conv_std_logic_vector(21615, 16),
33702 => conv_std_logic_vector(21746, 16),
33703 => conv_std_logic_vector(21877, 16),
33704 => conv_std_logic_vector(22008, 16),
33705 => conv_std_logic_vector(22139, 16),
33706 => conv_std_logic_vector(22270, 16),
33707 => conv_std_logic_vector(22401, 16),
33708 => conv_std_logic_vector(22532, 16),
33709 => conv_std_logic_vector(22663, 16),
33710 => conv_std_logic_vector(22794, 16),
33711 => conv_std_logic_vector(22925, 16),
33712 => conv_std_logic_vector(23056, 16),
33713 => conv_std_logic_vector(23187, 16),
33714 => conv_std_logic_vector(23318, 16),
33715 => conv_std_logic_vector(23449, 16),
33716 => conv_std_logic_vector(23580, 16),
33717 => conv_std_logic_vector(23711, 16),
33718 => conv_std_logic_vector(23842, 16),
33719 => conv_std_logic_vector(23973, 16),
33720 => conv_std_logic_vector(24104, 16),
33721 => conv_std_logic_vector(24235, 16),
33722 => conv_std_logic_vector(24366, 16),
33723 => conv_std_logic_vector(24497, 16),
33724 => conv_std_logic_vector(24628, 16),
33725 => conv_std_logic_vector(24759, 16),
33726 => conv_std_logic_vector(24890, 16),
33727 => conv_std_logic_vector(25021, 16),
33728 => conv_std_logic_vector(25152, 16),
33729 => conv_std_logic_vector(25283, 16),
33730 => conv_std_logic_vector(25414, 16),
33731 => conv_std_logic_vector(25545, 16),
33732 => conv_std_logic_vector(25676, 16),
33733 => conv_std_logic_vector(25807, 16),
33734 => conv_std_logic_vector(25938, 16),
33735 => conv_std_logic_vector(26069, 16),
33736 => conv_std_logic_vector(26200, 16),
33737 => conv_std_logic_vector(26331, 16),
33738 => conv_std_logic_vector(26462, 16),
33739 => conv_std_logic_vector(26593, 16),
33740 => conv_std_logic_vector(26724, 16),
33741 => conv_std_logic_vector(26855, 16),
33742 => conv_std_logic_vector(26986, 16),
33743 => conv_std_logic_vector(27117, 16),
33744 => conv_std_logic_vector(27248, 16),
33745 => conv_std_logic_vector(27379, 16),
33746 => conv_std_logic_vector(27510, 16),
33747 => conv_std_logic_vector(27641, 16),
33748 => conv_std_logic_vector(27772, 16),
33749 => conv_std_logic_vector(27903, 16),
33750 => conv_std_logic_vector(28034, 16),
33751 => conv_std_logic_vector(28165, 16),
33752 => conv_std_logic_vector(28296, 16),
33753 => conv_std_logic_vector(28427, 16),
33754 => conv_std_logic_vector(28558, 16),
33755 => conv_std_logic_vector(28689, 16),
33756 => conv_std_logic_vector(28820, 16),
33757 => conv_std_logic_vector(28951, 16),
33758 => conv_std_logic_vector(29082, 16),
33759 => conv_std_logic_vector(29213, 16),
33760 => conv_std_logic_vector(29344, 16),
33761 => conv_std_logic_vector(29475, 16),
33762 => conv_std_logic_vector(29606, 16),
33763 => conv_std_logic_vector(29737, 16),
33764 => conv_std_logic_vector(29868, 16),
33765 => conv_std_logic_vector(29999, 16),
33766 => conv_std_logic_vector(30130, 16),
33767 => conv_std_logic_vector(30261, 16),
33768 => conv_std_logic_vector(30392, 16),
33769 => conv_std_logic_vector(30523, 16),
33770 => conv_std_logic_vector(30654, 16),
33771 => conv_std_logic_vector(30785, 16),
33772 => conv_std_logic_vector(30916, 16),
33773 => conv_std_logic_vector(31047, 16),
33774 => conv_std_logic_vector(31178, 16),
33775 => conv_std_logic_vector(31309, 16),
33776 => conv_std_logic_vector(31440, 16),
33777 => conv_std_logic_vector(31571, 16),
33778 => conv_std_logic_vector(31702, 16),
33779 => conv_std_logic_vector(31833, 16),
33780 => conv_std_logic_vector(31964, 16),
33781 => conv_std_logic_vector(32095, 16),
33782 => conv_std_logic_vector(32226, 16),
33783 => conv_std_logic_vector(32357, 16),
33784 => conv_std_logic_vector(32488, 16),
33785 => conv_std_logic_vector(32619, 16),
33786 => conv_std_logic_vector(32750, 16),
33787 => conv_std_logic_vector(32881, 16),
33788 => conv_std_logic_vector(33012, 16),
33789 => conv_std_logic_vector(33143, 16),
33790 => conv_std_logic_vector(33274, 16),
33791 => conv_std_logic_vector(33405, 16),
33792 => conv_std_logic_vector(0, 16),
33793 => conv_std_logic_vector(132, 16),
33794 => conv_std_logic_vector(264, 16),
33795 => conv_std_logic_vector(396, 16),
33796 => conv_std_logic_vector(528, 16),
33797 => conv_std_logic_vector(660, 16),
33798 => conv_std_logic_vector(792, 16),
33799 => conv_std_logic_vector(924, 16),
33800 => conv_std_logic_vector(1056, 16),
33801 => conv_std_logic_vector(1188, 16),
33802 => conv_std_logic_vector(1320, 16),
33803 => conv_std_logic_vector(1452, 16),
33804 => conv_std_logic_vector(1584, 16),
33805 => conv_std_logic_vector(1716, 16),
33806 => conv_std_logic_vector(1848, 16),
33807 => conv_std_logic_vector(1980, 16),
33808 => conv_std_logic_vector(2112, 16),
33809 => conv_std_logic_vector(2244, 16),
33810 => conv_std_logic_vector(2376, 16),
33811 => conv_std_logic_vector(2508, 16),
33812 => conv_std_logic_vector(2640, 16),
33813 => conv_std_logic_vector(2772, 16),
33814 => conv_std_logic_vector(2904, 16),
33815 => conv_std_logic_vector(3036, 16),
33816 => conv_std_logic_vector(3168, 16),
33817 => conv_std_logic_vector(3300, 16),
33818 => conv_std_logic_vector(3432, 16),
33819 => conv_std_logic_vector(3564, 16),
33820 => conv_std_logic_vector(3696, 16),
33821 => conv_std_logic_vector(3828, 16),
33822 => conv_std_logic_vector(3960, 16),
33823 => conv_std_logic_vector(4092, 16),
33824 => conv_std_logic_vector(4224, 16),
33825 => conv_std_logic_vector(4356, 16),
33826 => conv_std_logic_vector(4488, 16),
33827 => conv_std_logic_vector(4620, 16),
33828 => conv_std_logic_vector(4752, 16),
33829 => conv_std_logic_vector(4884, 16),
33830 => conv_std_logic_vector(5016, 16),
33831 => conv_std_logic_vector(5148, 16),
33832 => conv_std_logic_vector(5280, 16),
33833 => conv_std_logic_vector(5412, 16),
33834 => conv_std_logic_vector(5544, 16),
33835 => conv_std_logic_vector(5676, 16),
33836 => conv_std_logic_vector(5808, 16),
33837 => conv_std_logic_vector(5940, 16),
33838 => conv_std_logic_vector(6072, 16),
33839 => conv_std_logic_vector(6204, 16),
33840 => conv_std_logic_vector(6336, 16),
33841 => conv_std_logic_vector(6468, 16),
33842 => conv_std_logic_vector(6600, 16),
33843 => conv_std_logic_vector(6732, 16),
33844 => conv_std_logic_vector(6864, 16),
33845 => conv_std_logic_vector(6996, 16),
33846 => conv_std_logic_vector(7128, 16),
33847 => conv_std_logic_vector(7260, 16),
33848 => conv_std_logic_vector(7392, 16),
33849 => conv_std_logic_vector(7524, 16),
33850 => conv_std_logic_vector(7656, 16),
33851 => conv_std_logic_vector(7788, 16),
33852 => conv_std_logic_vector(7920, 16),
33853 => conv_std_logic_vector(8052, 16),
33854 => conv_std_logic_vector(8184, 16),
33855 => conv_std_logic_vector(8316, 16),
33856 => conv_std_logic_vector(8448, 16),
33857 => conv_std_logic_vector(8580, 16),
33858 => conv_std_logic_vector(8712, 16),
33859 => conv_std_logic_vector(8844, 16),
33860 => conv_std_logic_vector(8976, 16),
33861 => conv_std_logic_vector(9108, 16),
33862 => conv_std_logic_vector(9240, 16),
33863 => conv_std_logic_vector(9372, 16),
33864 => conv_std_logic_vector(9504, 16),
33865 => conv_std_logic_vector(9636, 16),
33866 => conv_std_logic_vector(9768, 16),
33867 => conv_std_logic_vector(9900, 16),
33868 => conv_std_logic_vector(10032, 16),
33869 => conv_std_logic_vector(10164, 16),
33870 => conv_std_logic_vector(10296, 16),
33871 => conv_std_logic_vector(10428, 16),
33872 => conv_std_logic_vector(10560, 16),
33873 => conv_std_logic_vector(10692, 16),
33874 => conv_std_logic_vector(10824, 16),
33875 => conv_std_logic_vector(10956, 16),
33876 => conv_std_logic_vector(11088, 16),
33877 => conv_std_logic_vector(11220, 16),
33878 => conv_std_logic_vector(11352, 16),
33879 => conv_std_logic_vector(11484, 16),
33880 => conv_std_logic_vector(11616, 16),
33881 => conv_std_logic_vector(11748, 16),
33882 => conv_std_logic_vector(11880, 16),
33883 => conv_std_logic_vector(12012, 16),
33884 => conv_std_logic_vector(12144, 16),
33885 => conv_std_logic_vector(12276, 16),
33886 => conv_std_logic_vector(12408, 16),
33887 => conv_std_logic_vector(12540, 16),
33888 => conv_std_logic_vector(12672, 16),
33889 => conv_std_logic_vector(12804, 16),
33890 => conv_std_logic_vector(12936, 16),
33891 => conv_std_logic_vector(13068, 16),
33892 => conv_std_logic_vector(13200, 16),
33893 => conv_std_logic_vector(13332, 16),
33894 => conv_std_logic_vector(13464, 16),
33895 => conv_std_logic_vector(13596, 16),
33896 => conv_std_logic_vector(13728, 16),
33897 => conv_std_logic_vector(13860, 16),
33898 => conv_std_logic_vector(13992, 16),
33899 => conv_std_logic_vector(14124, 16),
33900 => conv_std_logic_vector(14256, 16),
33901 => conv_std_logic_vector(14388, 16),
33902 => conv_std_logic_vector(14520, 16),
33903 => conv_std_logic_vector(14652, 16),
33904 => conv_std_logic_vector(14784, 16),
33905 => conv_std_logic_vector(14916, 16),
33906 => conv_std_logic_vector(15048, 16),
33907 => conv_std_logic_vector(15180, 16),
33908 => conv_std_logic_vector(15312, 16),
33909 => conv_std_logic_vector(15444, 16),
33910 => conv_std_logic_vector(15576, 16),
33911 => conv_std_logic_vector(15708, 16),
33912 => conv_std_logic_vector(15840, 16),
33913 => conv_std_logic_vector(15972, 16),
33914 => conv_std_logic_vector(16104, 16),
33915 => conv_std_logic_vector(16236, 16),
33916 => conv_std_logic_vector(16368, 16),
33917 => conv_std_logic_vector(16500, 16),
33918 => conv_std_logic_vector(16632, 16),
33919 => conv_std_logic_vector(16764, 16),
33920 => conv_std_logic_vector(16896, 16),
33921 => conv_std_logic_vector(17028, 16),
33922 => conv_std_logic_vector(17160, 16),
33923 => conv_std_logic_vector(17292, 16),
33924 => conv_std_logic_vector(17424, 16),
33925 => conv_std_logic_vector(17556, 16),
33926 => conv_std_logic_vector(17688, 16),
33927 => conv_std_logic_vector(17820, 16),
33928 => conv_std_logic_vector(17952, 16),
33929 => conv_std_logic_vector(18084, 16),
33930 => conv_std_logic_vector(18216, 16),
33931 => conv_std_logic_vector(18348, 16),
33932 => conv_std_logic_vector(18480, 16),
33933 => conv_std_logic_vector(18612, 16),
33934 => conv_std_logic_vector(18744, 16),
33935 => conv_std_logic_vector(18876, 16),
33936 => conv_std_logic_vector(19008, 16),
33937 => conv_std_logic_vector(19140, 16),
33938 => conv_std_logic_vector(19272, 16),
33939 => conv_std_logic_vector(19404, 16),
33940 => conv_std_logic_vector(19536, 16),
33941 => conv_std_logic_vector(19668, 16),
33942 => conv_std_logic_vector(19800, 16),
33943 => conv_std_logic_vector(19932, 16),
33944 => conv_std_logic_vector(20064, 16),
33945 => conv_std_logic_vector(20196, 16),
33946 => conv_std_logic_vector(20328, 16),
33947 => conv_std_logic_vector(20460, 16),
33948 => conv_std_logic_vector(20592, 16),
33949 => conv_std_logic_vector(20724, 16),
33950 => conv_std_logic_vector(20856, 16),
33951 => conv_std_logic_vector(20988, 16),
33952 => conv_std_logic_vector(21120, 16),
33953 => conv_std_logic_vector(21252, 16),
33954 => conv_std_logic_vector(21384, 16),
33955 => conv_std_logic_vector(21516, 16),
33956 => conv_std_logic_vector(21648, 16),
33957 => conv_std_logic_vector(21780, 16),
33958 => conv_std_logic_vector(21912, 16),
33959 => conv_std_logic_vector(22044, 16),
33960 => conv_std_logic_vector(22176, 16),
33961 => conv_std_logic_vector(22308, 16),
33962 => conv_std_logic_vector(22440, 16),
33963 => conv_std_logic_vector(22572, 16),
33964 => conv_std_logic_vector(22704, 16),
33965 => conv_std_logic_vector(22836, 16),
33966 => conv_std_logic_vector(22968, 16),
33967 => conv_std_logic_vector(23100, 16),
33968 => conv_std_logic_vector(23232, 16),
33969 => conv_std_logic_vector(23364, 16),
33970 => conv_std_logic_vector(23496, 16),
33971 => conv_std_logic_vector(23628, 16),
33972 => conv_std_logic_vector(23760, 16),
33973 => conv_std_logic_vector(23892, 16),
33974 => conv_std_logic_vector(24024, 16),
33975 => conv_std_logic_vector(24156, 16),
33976 => conv_std_logic_vector(24288, 16),
33977 => conv_std_logic_vector(24420, 16),
33978 => conv_std_logic_vector(24552, 16),
33979 => conv_std_logic_vector(24684, 16),
33980 => conv_std_logic_vector(24816, 16),
33981 => conv_std_logic_vector(24948, 16),
33982 => conv_std_logic_vector(25080, 16),
33983 => conv_std_logic_vector(25212, 16),
33984 => conv_std_logic_vector(25344, 16),
33985 => conv_std_logic_vector(25476, 16),
33986 => conv_std_logic_vector(25608, 16),
33987 => conv_std_logic_vector(25740, 16),
33988 => conv_std_logic_vector(25872, 16),
33989 => conv_std_logic_vector(26004, 16),
33990 => conv_std_logic_vector(26136, 16),
33991 => conv_std_logic_vector(26268, 16),
33992 => conv_std_logic_vector(26400, 16),
33993 => conv_std_logic_vector(26532, 16),
33994 => conv_std_logic_vector(26664, 16),
33995 => conv_std_logic_vector(26796, 16),
33996 => conv_std_logic_vector(26928, 16),
33997 => conv_std_logic_vector(27060, 16),
33998 => conv_std_logic_vector(27192, 16),
33999 => conv_std_logic_vector(27324, 16),
34000 => conv_std_logic_vector(27456, 16),
34001 => conv_std_logic_vector(27588, 16),
34002 => conv_std_logic_vector(27720, 16),
34003 => conv_std_logic_vector(27852, 16),
34004 => conv_std_logic_vector(27984, 16),
34005 => conv_std_logic_vector(28116, 16),
34006 => conv_std_logic_vector(28248, 16),
34007 => conv_std_logic_vector(28380, 16),
34008 => conv_std_logic_vector(28512, 16),
34009 => conv_std_logic_vector(28644, 16),
34010 => conv_std_logic_vector(28776, 16),
34011 => conv_std_logic_vector(28908, 16),
34012 => conv_std_logic_vector(29040, 16),
34013 => conv_std_logic_vector(29172, 16),
34014 => conv_std_logic_vector(29304, 16),
34015 => conv_std_logic_vector(29436, 16),
34016 => conv_std_logic_vector(29568, 16),
34017 => conv_std_logic_vector(29700, 16),
34018 => conv_std_logic_vector(29832, 16),
34019 => conv_std_logic_vector(29964, 16),
34020 => conv_std_logic_vector(30096, 16),
34021 => conv_std_logic_vector(30228, 16),
34022 => conv_std_logic_vector(30360, 16),
34023 => conv_std_logic_vector(30492, 16),
34024 => conv_std_logic_vector(30624, 16),
34025 => conv_std_logic_vector(30756, 16),
34026 => conv_std_logic_vector(30888, 16),
34027 => conv_std_logic_vector(31020, 16),
34028 => conv_std_logic_vector(31152, 16),
34029 => conv_std_logic_vector(31284, 16),
34030 => conv_std_logic_vector(31416, 16),
34031 => conv_std_logic_vector(31548, 16),
34032 => conv_std_logic_vector(31680, 16),
34033 => conv_std_logic_vector(31812, 16),
34034 => conv_std_logic_vector(31944, 16),
34035 => conv_std_logic_vector(32076, 16),
34036 => conv_std_logic_vector(32208, 16),
34037 => conv_std_logic_vector(32340, 16),
34038 => conv_std_logic_vector(32472, 16),
34039 => conv_std_logic_vector(32604, 16),
34040 => conv_std_logic_vector(32736, 16),
34041 => conv_std_logic_vector(32868, 16),
34042 => conv_std_logic_vector(33000, 16),
34043 => conv_std_logic_vector(33132, 16),
34044 => conv_std_logic_vector(33264, 16),
34045 => conv_std_logic_vector(33396, 16),
34046 => conv_std_logic_vector(33528, 16),
34047 => conv_std_logic_vector(33660, 16),
34048 => conv_std_logic_vector(0, 16),
34049 => conv_std_logic_vector(133, 16),
34050 => conv_std_logic_vector(266, 16),
34051 => conv_std_logic_vector(399, 16),
34052 => conv_std_logic_vector(532, 16),
34053 => conv_std_logic_vector(665, 16),
34054 => conv_std_logic_vector(798, 16),
34055 => conv_std_logic_vector(931, 16),
34056 => conv_std_logic_vector(1064, 16),
34057 => conv_std_logic_vector(1197, 16),
34058 => conv_std_logic_vector(1330, 16),
34059 => conv_std_logic_vector(1463, 16),
34060 => conv_std_logic_vector(1596, 16),
34061 => conv_std_logic_vector(1729, 16),
34062 => conv_std_logic_vector(1862, 16),
34063 => conv_std_logic_vector(1995, 16),
34064 => conv_std_logic_vector(2128, 16),
34065 => conv_std_logic_vector(2261, 16),
34066 => conv_std_logic_vector(2394, 16),
34067 => conv_std_logic_vector(2527, 16),
34068 => conv_std_logic_vector(2660, 16),
34069 => conv_std_logic_vector(2793, 16),
34070 => conv_std_logic_vector(2926, 16),
34071 => conv_std_logic_vector(3059, 16),
34072 => conv_std_logic_vector(3192, 16),
34073 => conv_std_logic_vector(3325, 16),
34074 => conv_std_logic_vector(3458, 16),
34075 => conv_std_logic_vector(3591, 16),
34076 => conv_std_logic_vector(3724, 16),
34077 => conv_std_logic_vector(3857, 16),
34078 => conv_std_logic_vector(3990, 16),
34079 => conv_std_logic_vector(4123, 16),
34080 => conv_std_logic_vector(4256, 16),
34081 => conv_std_logic_vector(4389, 16),
34082 => conv_std_logic_vector(4522, 16),
34083 => conv_std_logic_vector(4655, 16),
34084 => conv_std_logic_vector(4788, 16),
34085 => conv_std_logic_vector(4921, 16),
34086 => conv_std_logic_vector(5054, 16),
34087 => conv_std_logic_vector(5187, 16),
34088 => conv_std_logic_vector(5320, 16),
34089 => conv_std_logic_vector(5453, 16),
34090 => conv_std_logic_vector(5586, 16),
34091 => conv_std_logic_vector(5719, 16),
34092 => conv_std_logic_vector(5852, 16),
34093 => conv_std_logic_vector(5985, 16),
34094 => conv_std_logic_vector(6118, 16),
34095 => conv_std_logic_vector(6251, 16),
34096 => conv_std_logic_vector(6384, 16),
34097 => conv_std_logic_vector(6517, 16),
34098 => conv_std_logic_vector(6650, 16),
34099 => conv_std_logic_vector(6783, 16),
34100 => conv_std_logic_vector(6916, 16),
34101 => conv_std_logic_vector(7049, 16),
34102 => conv_std_logic_vector(7182, 16),
34103 => conv_std_logic_vector(7315, 16),
34104 => conv_std_logic_vector(7448, 16),
34105 => conv_std_logic_vector(7581, 16),
34106 => conv_std_logic_vector(7714, 16),
34107 => conv_std_logic_vector(7847, 16),
34108 => conv_std_logic_vector(7980, 16),
34109 => conv_std_logic_vector(8113, 16),
34110 => conv_std_logic_vector(8246, 16),
34111 => conv_std_logic_vector(8379, 16),
34112 => conv_std_logic_vector(8512, 16),
34113 => conv_std_logic_vector(8645, 16),
34114 => conv_std_logic_vector(8778, 16),
34115 => conv_std_logic_vector(8911, 16),
34116 => conv_std_logic_vector(9044, 16),
34117 => conv_std_logic_vector(9177, 16),
34118 => conv_std_logic_vector(9310, 16),
34119 => conv_std_logic_vector(9443, 16),
34120 => conv_std_logic_vector(9576, 16),
34121 => conv_std_logic_vector(9709, 16),
34122 => conv_std_logic_vector(9842, 16),
34123 => conv_std_logic_vector(9975, 16),
34124 => conv_std_logic_vector(10108, 16),
34125 => conv_std_logic_vector(10241, 16),
34126 => conv_std_logic_vector(10374, 16),
34127 => conv_std_logic_vector(10507, 16),
34128 => conv_std_logic_vector(10640, 16),
34129 => conv_std_logic_vector(10773, 16),
34130 => conv_std_logic_vector(10906, 16),
34131 => conv_std_logic_vector(11039, 16),
34132 => conv_std_logic_vector(11172, 16),
34133 => conv_std_logic_vector(11305, 16),
34134 => conv_std_logic_vector(11438, 16),
34135 => conv_std_logic_vector(11571, 16),
34136 => conv_std_logic_vector(11704, 16),
34137 => conv_std_logic_vector(11837, 16),
34138 => conv_std_logic_vector(11970, 16),
34139 => conv_std_logic_vector(12103, 16),
34140 => conv_std_logic_vector(12236, 16),
34141 => conv_std_logic_vector(12369, 16),
34142 => conv_std_logic_vector(12502, 16),
34143 => conv_std_logic_vector(12635, 16),
34144 => conv_std_logic_vector(12768, 16),
34145 => conv_std_logic_vector(12901, 16),
34146 => conv_std_logic_vector(13034, 16),
34147 => conv_std_logic_vector(13167, 16),
34148 => conv_std_logic_vector(13300, 16),
34149 => conv_std_logic_vector(13433, 16),
34150 => conv_std_logic_vector(13566, 16),
34151 => conv_std_logic_vector(13699, 16),
34152 => conv_std_logic_vector(13832, 16),
34153 => conv_std_logic_vector(13965, 16),
34154 => conv_std_logic_vector(14098, 16),
34155 => conv_std_logic_vector(14231, 16),
34156 => conv_std_logic_vector(14364, 16),
34157 => conv_std_logic_vector(14497, 16),
34158 => conv_std_logic_vector(14630, 16),
34159 => conv_std_logic_vector(14763, 16),
34160 => conv_std_logic_vector(14896, 16),
34161 => conv_std_logic_vector(15029, 16),
34162 => conv_std_logic_vector(15162, 16),
34163 => conv_std_logic_vector(15295, 16),
34164 => conv_std_logic_vector(15428, 16),
34165 => conv_std_logic_vector(15561, 16),
34166 => conv_std_logic_vector(15694, 16),
34167 => conv_std_logic_vector(15827, 16),
34168 => conv_std_logic_vector(15960, 16),
34169 => conv_std_logic_vector(16093, 16),
34170 => conv_std_logic_vector(16226, 16),
34171 => conv_std_logic_vector(16359, 16),
34172 => conv_std_logic_vector(16492, 16),
34173 => conv_std_logic_vector(16625, 16),
34174 => conv_std_logic_vector(16758, 16),
34175 => conv_std_logic_vector(16891, 16),
34176 => conv_std_logic_vector(17024, 16),
34177 => conv_std_logic_vector(17157, 16),
34178 => conv_std_logic_vector(17290, 16),
34179 => conv_std_logic_vector(17423, 16),
34180 => conv_std_logic_vector(17556, 16),
34181 => conv_std_logic_vector(17689, 16),
34182 => conv_std_logic_vector(17822, 16),
34183 => conv_std_logic_vector(17955, 16),
34184 => conv_std_logic_vector(18088, 16),
34185 => conv_std_logic_vector(18221, 16),
34186 => conv_std_logic_vector(18354, 16),
34187 => conv_std_logic_vector(18487, 16),
34188 => conv_std_logic_vector(18620, 16),
34189 => conv_std_logic_vector(18753, 16),
34190 => conv_std_logic_vector(18886, 16),
34191 => conv_std_logic_vector(19019, 16),
34192 => conv_std_logic_vector(19152, 16),
34193 => conv_std_logic_vector(19285, 16),
34194 => conv_std_logic_vector(19418, 16),
34195 => conv_std_logic_vector(19551, 16),
34196 => conv_std_logic_vector(19684, 16),
34197 => conv_std_logic_vector(19817, 16),
34198 => conv_std_logic_vector(19950, 16),
34199 => conv_std_logic_vector(20083, 16),
34200 => conv_std_logic_vector(20216, 16),
34201 => conv_std_logic_vector(20349, 16),
34202 => conv_std_logic_vector(20482, 16),
34203 => conv_std_logic_vector(20615, 16),
34204 => conv_std_logic_vector(20748, 16),
34205 => conv_std_logic_vector(20881, 16),
34206 => conv_std_logic_vector(21014, 16),
34207 => conv_std_logic_vector(21147, 16),
34208 => conv_std_logic_vector(21280, 16),
34209 => conv_std_logic_vector(21413, 16),
34210 => conv_std_logic_vector(21546, 16),
34211 => conv_std_logic_vector(21679, 16),
34212 => conv_std_logic_vector(21812, 16),
34213 => conv_std_logic_vector(21945, 16),
34214 => conv_std_logic_vector(22078, 16),
34215 => conv_std_logic_vector(22211, 16),
34216 => conv_std_logic_vector(22344, 16),
34217 => conv_std_logic_vector(22477, 16),
34218 => conv_std_logic_vector(22610, 16),
34219 => conv_std_logic_vector(22743, 16),
34220 => conv_std_logic_vector(22876, 16),
34221 => conv_std_logic_vector(23009, 16),
34222 => conv_std_logic_vector(23142, 16),
34223 => conv_std_logic_vector(23275, 16),
34224 => conv_std_logic_vector(23408, 16),
34225 => conv_std_logic_vector(23541, 16),
34226 => conv_std_logic_vector(23674, 16),
34227 => conv_std_logic_vector(23807, 16),
34228 => conv_std_logic_vector(23940, 16),
34229 => conv_std_logic_vector(24073, 16),
34230 => conv_std_logic_vector(24206, 16),
34231 => conv_std_logic_vector(24339, 16),
34232 => conv_std_logic_vector(24472, 16),
34233 => conv_std_logic_vector(24605, 16),
34234 => conv_std_logic_vector(24738, 16),
34235 => conv_std_logic_vector(24871, 16),
34236 => conv_std_logic_vector(25004, 16),
34237 => conv_std_logic_vector(25137, 16),
34238 => conv_std_logic_vector(25270, 16),
34239 => conv_std_logic_vector(25403, 16),
34240 => conv_std_logic_vector(25536, 16),
34241 => conv_std_logic_vector(25669, 16),
34242 => conv_std_logic_vector(25802, 16),
34243 => conv_std_logic_vector(25935, 16),
34244 => conv_std_logic_vector(26068, 16),
34245 => conv_std_logic_vector(26201, 16),
34246 => conv_std_logic_vector(26334, 16),
34247 => conv_std_logic_vector(26467, 16),
34248 => conv_std_logic_vector(26600, 16),
34249 => conv_std_logic_vector(26733, 16),
34250 => conv_std_logic_vector(26866, 16),
34251 => conv_std_logic_vector(26999, 16),
34252 => conv_std_logic_vector(27132, 16),
34253 => conv_std_logic_vector(27265, 16),
34254 => conv_std_logic_vector(27398, 16),
34255 => conv_std_logic_vector(27531, 16),
34256 => conv_std_logic_vector(27664, 16),
34257 => conv_std_logic_vector(27797, 16),
34258 => conv_std_logic_vector(27930, 16),
34259 => conv_std_logic_vector(28063, 16),
34260 => conv_std_logic_vector(28196, 16),
34261 => conv_std_logic_vector(28329, 16),
34262 => conv_std_logic_vector(28462, 16),
34263 => conv_std_logic_vector(28595, 16),
34264 => conv_std_logic_vector(28728, 16),
34265 => conv_std_logic_vector(28861, 16),
34266 => conv_std_logic_vector(28994, 16),
34267 => conv_std_logic_vector(29127, 16),
34268 => conv_std_logic_vector(29260, 16),
34269 => conv_std_logic_vector(29393, 16),
34270 => conv_std_logic_vector(29526, 16),
34271 => conv_std_logic_vector(29659, 16),
34272 => conv_std_logic_vector(29792, 16),
34273 => conv_std_logic_vector(29925, 16),
34274 => conv_std_logic_vector(30058, 16),
34275 => conv_std_logic_vector(30191, 16),
34276 => conv_std_logic_vector(30324, 16),
34277 => conv_std_logic_vector(30457, 16),
34278 => conv_std_logic_vector(30590, 16),
34279 => conv_std_logic_vector(30723, 16),
34280 => conv_std_logic_vector(30856, 16),
34281 => conv_std_logic_vector(30989, 16),
34282 => conv_std_logic_vector(31122, 16),
34283 => conv_std_logic_vector(31255, 16),
34284 => conv_std_logic_vector(31388, 16),
34285 => conv_std_logic_vector(31521, 16),
34286 => conv_std_logic_vector(31654, 16),
34287 => conv_std_logic_vector(31787, 16),
34288 => conv_std_logic_vector(31920, 16),
34289 => conv_std_logic_vector(32053, 16),
34290 => conv_std_logic_vector(32186, 16),
34291 => conv_std_logic_vector(32319, 16),
34292 => conv_std_logic_vector(32452, 16),
34293 => conv_std_logic_vector(32585, 16),
34294 => conv_std_logic_vector(32718, 16),
34295 => conv_std_logic_vector(32851, 16),
34296 => conv_std_logic_vector(32984, 16),
34297 => conv_std_logic_vector(33117, 16),
34298 => conv_std_logic_vector(33250, 16),
34299 => conv_std_logic_vector(33383, 16),
34300 => conv_std_logic_vector(33516, 16),
34301 => conv_std_logic_vector(33649, 16),
34302 => conv_std_logic_vector(33782, 16),
34303 => conv_std_logic_vector(33915, 16),
34304 => conv_std_logic_vector(0, 16),
34305 => conv_std_logic_vector(134, 16),
34306 => conv_std_logic_vector(268, 16),
34307 => conv_std_logic_vector(402, 16),
34308 => conv_std_logic_vector(536, 16),
34309 => conv_std_logic_vector(670, 16),
34310 => conv_std_logic_vector(804, 16),
34311 => conv_std_logic_vector(938, 16),
34312 => conv_std_logic_vector(1072, 16),
34313 => conv_std_logic_vector(1206, 16),
34314 => conv_std_logic_vector(1340, 16),
34315 => conv_std_logic_vector(1474, 16),
34316 => conv_std_logic_vector(1608, 16),
34317 => conv_std_logic_vector(1742, 16),
34318 => conv_std_logic_vector(1876, 16),
34319 => conv_std_logic_vector(2010, 16),
34320 => conv_std_logic_vector(2144, 16),
34321 => conv_std_logic_vector(2278, 16),
34322 => conv_std_logic_vector(2412, 16),
34323 => conv_std_logic_vector(2546, 16),
34324 => conv_std_logic_vector(2680, 16),
34325 => conv_std_logic_vector(2814, 16),
34326 => conv_std_logic_vector(2948, 16),
34327 => conv_std_logic_vector(3082, 16),
34328 => conv_std_logic_vector(3216, 16),
34329 => conv_std_logic_vector(3350, 16),
34330 => conv_std_logic_vector(3484, 16),
34331 => conv_std_logic_vector(3618, 16),
34332 => conv_std_logic_vector(3752, 16),
34333 => conv_std_logic_vector(3886, 16),
34334 => conv_std_logic_vector(4020, 16),
34335 => conv_std_logic_vector(4154, 16),
34336 => conv_std_logic_vector(4288, 16),
34337 => conv_std_logic_vector(4422, 16),
34338 => conv_std_logic_vector(4556, 16),
34339 => conv_std_logic_vector(4690, 16),
34340 => conv_std_logic_vector(4824, 16),
34341 => conv_std_logic_vector(4958, 16),
34342 => conv_std_logic_vector(5092, 16),
34343 => conv_std_logic_vector(5226, 16),
34344 => conv_std_logic_vector(5360, 16),
34345 => conv_std_logic_vector(5494, 16),
34346 => conv_std_logic_vector(5628, 16),
34347 => conv_std_logic_vector(5762, 16),
34348 => conv_std_logic_vector(5896, 16),
34349 => conv_std_logic_vector(6030, 16),
34350 => conv_std_logic_vector(6164, 16),
34351 => conv_std_logic_vector(6298, 16),
34352 => conv_std_logic_vector(6432, 16),
34353 => conv_std_logic_vector(6566, 16),
34354 => conv_std_logic_vector(6700, 16),
34355 => conv_std_logic_vector(6834, 16),
34356 => conv_std_logic_vector(6968, 16),
34357 => conv_std_logic_vector(7102, 16),
34358 => conv_std_logic_vector(7236, 16),
34359 => conv_std_logic_vector(7370, 16),
34360 => conv_std_logic_vector(7504, 16),
34361 => conv_std_logic_vector(7638, 16),
34362 => conv_std_logic_vector(7772, 16),
34363 => conv_std_logic_vector(7906, 16),
34364 => conv_std_logic_vector(8040, 16),
34365 => conv_std_logic_vector(8174, 16),
34366 => conv_std_logic_vector(8308, 16),
34367 => conv_std_logic_vector(8442, 16),
34368 => conv_std_logic_vector(8576, 16),
34369 => conv_std_logic_vector(8710, 16),
34370 => conv_std_logic_vector(8844, 16),
34371 => conv_std_logic_vector(8978, 16),
34372 => conv_std_logic_vector(9112, 16),
34373 => conv_std_logic_vector(9246, 16),
34374 => conv_std_logic_vector(9380, 16),
34375 => conv_std_logic_vector(9514, 16),
34376 => conv_std_logic_vector(9648, 16),
34377 => conv_std_logic_vector(9782, 16),
34378 => conv_std_logic_vector(9916, 16),
34379 => conv_std_logic_vector(10050, 16),
34380 => conv_std_logic_vector(10184, 16),
34381 => conv_std_logic_vector(10318, 16),
34382 => conv_std_logic_vector(10452, 16),
34383 => conv_std_logic_vector(10586, 16),
34384 => conv_std_logic_vector(10720, 16),
34385 => conv_std_logic_vector(10854, 16),
34386 => conv_std_logic_vector(10988, 16),
34387 => conv_std_logic_vector(11122, 16),
34388 => conv_std_logic_vector(11256, 16),
34389 => conv_std_logic_vector(11390, 16),
34390 => conv_std_logic_vector(11524, 16),
34391 => conv_std_logic_vector(11658, 16),
34392 => conv_std_logic_vector(11792, 16),
34393 => conv_std_logic_vector(11926, 16),
34394 => conv_std_logic_vector(12060, 16),
34395 => conv_std_logic_vector(12194, 16),
34396 => conv_std_logic_vector(12328, 16),
34397 => conv_std_logic_vector(12462, 16),
34398 => conv_std_logic_vector(12596, 16),
34399 => conv_std_logic_vector(12730, 16),
34400 => conv_std_logic_vector(12864, 16),
34401 => conv_std_logic_vector(12998, 16),
34402 => conv_std_logic_vector(13132, 16),
34403 => conv_std_logic_vector(13266, 16),
34404 => conv_std_logic_vector(13400, 16),
34405 => conv_std_logic_vector(13534, 16),
34406 => conv_std_logic_vector(13668, 16),
34407 => conv_std_logic_vector(13802, 16),
34408 => conv_std_logic_vector(13936, 16),
34409 => conv_std_logic_vector(14070, 16),
34410 => conv_std_logic_vector(14204, 16),
34411 => conv_std_logic_vector(14338, 16),
34412 => conv_std_logic_vector(14472, 16),
34413 => conv_std_logic_vector(14606, 16),
34414 => conv_std_logic_vector(14740, 16),
34415 => conv_std_logic_vector(14874, 16),
34416 => conv_std_logic_vector(15008, 16),
34417 => conv_std_logic_vector(15142, 16),
34418 => conv_std_logic_vector(15276, 16),
34419 => conv_std_logic_vector(15410, 16),
34420 => conv_std_logic_vector(15544, 16),
34421 => conv_std_logic_vector(15678, 16),
34422 => conv_std_logic_vector(15812, 16),
34423 => conv_std_logic_vector(15946, 16),
34424 => conv_std_logic_vector(16080, 16),
34425 => conv_std_logic_vector(16214, 16),
34426 => conv_std_logic_vector(16348, 16),
34427 => conv_std_logic_vector(16482, 16),
34428 => conv_std_logic_vector(16616, 16),
34429 => conv_std_logic_vector(16750, 16),
34430 => conv_std_logic_vector(16884, 16),
34431 => conv_std_logic_vector(17018, 16),
34432 => conv_std_logic_vector(17152, 16),
34433 => conv_std_logic_vector(17286, 16),
34434 => conv_std_logic_vector(17420, 16),
34435 => conv_std_logic_vector(17554, 16),
34436 => conv_std_logic_vector(17688, 16),
34437 => conv_std_logic_vector(17822, 16),
34438 => conv_std_logic_vector(17956, 16),
34439 => conv_std_logic_vector(18090, 16),
34440 => conv_std_logic_vector(18224, 16),
34441 => conv_std_logic_vector(18358, 16),
34442 => conv_std_logic_vector(18492, 16),
34443 => conv_std_logic_vector(18626, 16),
34444 => conv_std_logic_vector(18760, 16),
34445 => conv_std_logic_vector(18894, 16),
34446 => conv_std_logic_vector(19028, 16),
34447 => conv_std_logic_vector(19162, 16),
34448 => conv_std_logic_vector(19296, 16),
34449 => conv_std_logic_vector(19430, 16),
34450 => conv_std_logic_vector(19564, 16),
34451 => conv_std_logic_vector(19698, 16),
34452 => conv_std_logic_vector(19832, 16),
34453 => conv_std_logic_vector(19966, 16),
34454 => conv_std_logic_vector(20100, 16),
34455 => conv_std_logic_vector(20234, 16),
34456 => conv_std_logic_vector(20368, 16),
34457 => conv_std_logic_vector(20502, 16),
34458 => conv_std_logic_vector(20636, 16),
34459 => conv_std_logic_vector(20770, 16),
34460 => conv_std_logic_vector(20904, 16),
34461 => conv_std_logic_vector(21038, 16),
34462 => conv_std_logic_vector(21172, 16),
34463 => conv_std_logic_vector(21306, 16),
34464 => conv_std_logic_vector(21440, 16),
34465 => conv_std_logic_vector(21574, 16),
34466 => conv_std_logic_vector(21708, 16),
34467 => conv_std_logic_vector(21842, 16),
34468 => conv_std_logic_vector(21976, 16),
34469 => conv_std_logic_vector(22110, 16),
34470 => conv_std_logic_vector(22244, 16),
34471 => conv_std_logic_vector(22378, 16),
34472 => conv_std_logic_vector(22512, 16),
34473 => conv_std_logic_vector(22646, 16),
34474 => conv_std_logic_vector(22780, 16),
34475 => conv_std_logic_vector(22914, 16),
34476 => conv_std_logic_vector(23048, 16),
34477 => conv_std_logic_vector(23182, 16),
34478 => conv_std_logic_vector(23316, 16),
34479 => conv_std_logic_vector(23450, 16),
34480 => conv_std_logic_vector(23584, 16),
34481 => conv_std_logic_vector(23718, 16),
34482 => conv_std_logic_vector(23852, 16),
34483 => conv_std_logic_vector(23986, 16),
34484 => conv_std_logic_vector(24120, 16),
34485 => conv_std_logic_vector(24254, 16),
34486 => conv_std_logic_vector(24388, 16),
34487 => conv_std_logic_vector(24522, 16),
34488 => conv_std_logic_vector(24656, 16),
34489 => conv_std_logic_vector(24790, 16),
34490 => conv_std_logic_vector(24924, 16),
34491 => conv_std_logic_vector(25058, 16),
34492 => conv_std_logic_vector(25192, 16),
34493 => conv_std_logic_vector(25326, 16),
34494 => conv_std_logic_vector(25460, 16),
34495 => conv_std_logic_vector(25594, 16),
34496 => conv_std_logic_vector(25728, 16),
34497 => conv_std_logic_vector(25862, 16),
34498 => conv_std_logic_vector(25996, 16),
34499 => conv_std_logic_vector(26130, 16),
34500 => conv_std_logic_vector(26264, 16),
34501 => conv_std_logic_vector(26398, 16),
34502 => conv_std_logic_vector(26532, 16),
34503 => conv_std_logic_vector(26666, 16),
34504 => conv_std_logic_vector(26800, 16),
34505 => conv_std_logic_vector(26934, 16),
34506 => conv_std_logic_vector(27068, 16),
34507 => conv_std_logic_vector(27202, 16),
34508 => conv_std_logic_vector(27336, 16),
34509 => conv_std_logic_vector(27470, 16),
34510 => conv_std_logic_vector(27604, 16),
34511 => conv_std_logic_vector(27738, 16),
34512 => conv_std_logic_vector(27872, 16),
34513 => conv_std_logic_vector(28006, 16),
34514 => conv_std_logic_vector(28140, 16),
34515 => conv_std_logic_vector(28274, 16),
34516 => conv_std_logic_vector(28408, 16),
34517 => conv_std_logic_vector(28542, 16),
34518 => conv_std_logic_vector(28676, 16),
34519 => conv_std_logic_vector(28810, 16),
34520 => conv_std_logic_vector(28944, 16),
34521 => conv_std_logic_vector(29078, 16),
34522 => conv_std_logic_vector(29212, 16),
34523 => conv_std_logic_vector(29346, 16),
34524 => conv_std_logic_vector(29480, 16),
34525 => conv_std_logic_vector(29614, 16),
34526 => conv_std_logic_vector(29748, 16),
34527 => conv_std_logic_vector(29882, 16),
34528 => conv_std_logic_vector(30016, 16),
34529 => conv_std_logic_vector(30150, 16),
34530 => conv_std_logic_vector(30284, 16),
34531 => conv_std_logic_vector(30418, 16),
34532 => conv_std_logic_vector(30552, 16),
34533 => conv_std_logic_vector(30686, 16),
34534 => conv_std_logic_vector(30820, 16),
34535 => conv_std_logic_vector(30954, 16),
34536 => conv_std_logic_vector(31088, 16),
34537 => conv_std_logic_vector(31222, 16),
34538 => conv_std_logic_vector(31356, 16),
34539 => conv_std_logic_vector(31490, 16),
34540 => conv_std_logic_vector(31624, 16),
34541 => conv_std_logic_vector(31758, 16),
34542 => conv_std_logic_vector(31892, 16),
34543 => conv_std_logic_vector(32026, 16),
34544 => conv_std_logic_vector(32160, 16),
34545 => conv_std_logic_vector(32294, 16),
34546 => conv_std_logic_vector(32428, 16),
34547 => conv_std_logic_vector(32562, 16),
34548 => conv_std_logic_vector(32696, 16),
34549 => conv_std_logic_vector(32830, 16),
34550 => conv_std_logic_vector(32964, 16),
34551 => conv_std_logic_vector(33098, 16),
34552 => conv_std_logic_vector(33232, 16),
34553 => conv_std_logic_vector(33366, 16),
34554 => conv_std_logic_vector(33500, 16),
34555 => conv_std_logic_vector(33634, 16),
34556 => conv_std_logic_vector(33768, 16),
34557 => conv_std_logic_vector(33902, 16),
34558 => conv_std_logic_vector(34036, 16),
34559 => conv_std_logic_vector(34170, 16),
34560 => conv_std_logic_vector(0, 16),
34561 => conv_std_logic_vector(135, 16),
34562 => conv_std_logic_vector(270, 16),
34563 => conv_std_logic_vector(405, 16),
34564 => conv_std_logic_vector(540, 16),
34565 => conv_std_logic_vector(675, 16),
34566 => conv_std_logic_vector(810, 16),
34567 => conv_std_logic_vector(945, 16),
34568 => conv_std_logic_vector(1080, 16),
34569 => conv_std_logic_vector(1215, 16),
34570 => conv_std_logic_vector(1350, 16),
34571 => conv_std_logic_vector(1485, 16),
34572 => conv_std_logic_vector(1620, 16),
34573 => conv_std_logic_vector(1755, 16),
34574 => conv_std_logic_vector(1890, 16),
34575 => conv_std_logic_vector(2025, 16),
34576 => conv_std_logic_vector(2160, 16),
34577 => conv_std_logic_vector(2295, 16),
34578 => conv_std_logic_vector(2430, 16),
34579 => conv_std_logic_vector(2565, 16),
34580 => conv_std_logic_vector(2700, 16),
34581 => conv_std_logic_vector(2835, 16),
34582 => conv_std_logic_vector(2970, 16),
34583 => conv_std_logic_vector(3105, 16),
34584 => conv_std_logic_vector(3240, 16),
34585 => conv_std_logic_vector(3375, 16),
34586 => conv_std_logic_vector(3510, 16),
34587 => conv_std_logic_vector(3645, 16),
34588 => conv_std_logic_vector(3780, 16),
34589 => conv_std_logic_vector(3915, 16),
34590 => conv_std_logic_vector(4050, 16),
34591 => conv_std_logic_vector(4185, 16),
34592 => conv_std_logic_vector(4320, 16),
34593 => conv_std_logic_vector(4455, 16),
34594 => conv_std_logic_vector(4590, 16),
34595 => conv_std_logic_vector(4725, 16),
34596 => conv_std_logic_vector(4860, 16),
34597 => conv_std_logic_vector(4995, 16),
34598 => conv_std_logic_vector(5130, 16),
34599 => conv_std_logic_vector(5265, 16),
34600 => conv_std_logic_vector(5400, 16),
34601 => conv_std_logic_vector(5535, 16),
34602 => conv_std_logic_vector(5670, 16),
34603 => conv_std_logic_vector(5805, 16),
34604 => conv_std_logic_vector(5940, 16),
34605 => conv_std_logic_vector(6075, 16),
34606 => conv_std_logic_vector(6210, 16),
34607 => conv_std_logic_vector(6345, 16),
34608 => conv_std_logic_vector(6480, 16),
34609 => conv_std_logic_vector(6615, 16),
34610 => conv_std_logic_vector(6750, 16),
34611 => conv_std_logic_vector(6885, 16),
34612 => conv_std_logic_vector(7020, 16),
34613 => conv_std_logic_vector(7155, 16),
34614 => conv_std_logic_vector(7290, 16),
34615 => conv_std_logic_vector(7425, 16),
34616 => conv_std_logic_vector(7560, 16),
34617 => conv_std_logic_vector(7695, 16),
34618 => conv_std_logic_vector(7830, 16),
34619 => conv_std_logic_vector(7965, 16),
34620 => conv_std_logic_vector(8100, 16),
34621 => conv_std_logic_vector(8235, 16),
34622 => conv_std_logic_vector(8370, 16),
34623 => conv_std_logic_vector(8505, 16),
34624 => conv_std_logic_vector(8640, 16),
34625 => conv_std_logic_vector(8775, 16),
34626 => conv_std_logic_vector(8910, 16),
34627 => conv_std_logic_vector(9045, 16),
34628 => conv_std_logic_vector(9180, 16),
34629 => conv_std_logic_vector(9315, 16),
34630 => conv_std_logic_vector(9450, 16),
34631 => conv_std_logic_vector(9585, 16),
34632 => conv_std_logic_vector(9720, 16),
34633 => conv_std_logic_vector(9855, 16),
34634 => conv_std_logic_vector(9990, 16),
34635 => conv_std_logic_vector(10125, 16),
34636 => conv_std_logic_vector(10260, 16),
34637 => conv_std_logic_vector(10395, 16),
34638 => conv_std_logic_vector(10530, 16),
34639 => conv_std_logic_vector(10665, 16),
34640 => conv_std_logic_vector(10800, 16),
34641 => conv_std_logic_vector(10935, 16),
34642 => conv_std_logic_vector(11070, 16),
34643 => conv_std_logic_vector(11205, 16),
34644 => conv_std_logic_vector(11340, 16),
34645 => conv_std_logic_vector(11475, 16),
34646 => conv_std_logic_vector(11610, 16),
34647 => conv_std_logic_vector(11745, 16),
34648 => conv_std_logic_vector(11880, 16),
34649 => conv_std_logic_vector(12015, 16),
34650 => conv_std_logic_vector(12150, 16),
34651 => conv_std_logic_vector(12285, 16),
34652 => conv_std_logic_vector(12420, 16),
34653 => conv_std_logic_vector(12555, 16),
34654 => conv_std_logic_vector(12690, 16),
34655 => conv_std_logic_vector(12825, 16),
34656 => conv_std_logic_vector(12960, 16),
34657 => conv_std_logic_vector(13095, 16),
34658 => conv_std_logic_vector(13230, 16),
34659 => conv_std_logic_vector(13365, 16),
34660 => conv_std_logic_vector(13500, 16),
34661 => conv_std_logic_vector(13635, 16),
34662 => conv_std_logic_vector(13770, 16),
34663 => conv_std_logic_vector(13905, 16),
34664 => conv_std_logic_vector(14040, 16),
34665 => conv_std_logic_vector(14175, 16),
34666 => conv_std_logic_vector(14310, 16),
34667 => conv_std_logic_vector(14445, 16),
34668 => conv_std_logic_vector(14580, 16),
34669 => conv_std_logic_vector(14715, 16),
34670 => conv_std_logic_vector(14850, 16),
34671 => conv_std_logic_vector(14985, 16),
34672 => conv_std_logic_vector(15120, 16),
34673 => conv_std_logic_vector(15255, 16),
34674 => conv_std_logic_vector(15390, 16),
34675 => conv_std_logic_vector(15525, 16),
34676 => conv_std_logic_vector(15660, 16),
34677 => conv_std_logic_vector(15795, 16),
34678 => conv_std_logic_vector(15930, 16),
34679 => conv_std_logic_vector(16065, 16),
34680 => conv_std_logic_vector(16200, 16),
34681 => conv_std_logic_vector(16335, 16),
34682 => conv_std_logic_vector(16470, 16),
34683 => conv_std_logic_vector(16605, 16),
34684 => conv_std_logic_vector(16740, 16),
34685 => conv_std_logic_vector(16875, 16),
34686 => conv_std_logic_vector(17010, 16),
34687 => conv_std_logic_vector(17145, 16),
34688 => conv_std_logic_vector(17280, 16),
34689 => conv_std_logic_vector(17415, 16),
34690 => conv_std_logic_vector(17550, 16),
34691 => conv_std_logic_vector(17685, 16),
34692 => conv_std_logic_vector(17820, 16),
34693 => conv_std_logic_vector(17955, 16),
34694 => conv_std_logic_vector(18090, 16),
34695 => conv_std_logic_vector(18225, 16),
34696 => conv_std_logic_vector(18360, 16),
34697 => conv_std_logic_vector(18495, 16),
34698 => conv_std_logic_vector(18630, 16),
34699 => conv_std_logic_vector(18765, 16),
34700 => conv_std_logic_vector(18900, 16),
34701 => conv_std_logic_vector(19035, 16),
34702 => conv_std_logic_vector(19170, 16),
34703 => conv_std_logic_vector(19305, 16),
34704 => conv_std_logic_vector(19440, 16),
34705 => conv_std_logic_vector(19575, 16),
34706 => conv_std_logic_vector(19710, 16),
34707 => conv_std_logic_vector(19845, 16),
34708 => conv_std_logic_vector(19980, 16),
34709 => conv_std_logic_vector(20115, 16),
34710 => conv_std_logic_vector(20250, 16),
34711 => conv_std_logic_vector(20385, 16),
34712 => conv_std_logic_vector(20520, 16),
34713 => conv_std_logic_vector(20655, 16),
34714 => conv_std_logic_vector(20790, 16),
34715 => conv_std_logic_vector(20925, 16),
34716 => conv_std_logic_vector(21060, 16),
34717 => conv_std_logic_vector(21195, 16),
34718 => conv_std_logic_vector(21330, 16),
34719 => conv_std_logic_vector(21465, 16),
34720 => conv_std_logic_vector(21600, 16),
34721 => conv_std_logic_vector(21735, 16),
34722 => conv_std_logic_vector(21870, 16),
34723 => conv_std_logic_vector(22005, 16),
34724 => conv_std_logic_vector(22140, 16),
34725 => conv_std_logic_vector(22275, 16),
34726 => conv_std_logic_vector(22410, 16),
34727 => conv_std_logic_vector(22545, 16),
34728 => conv_std_logic_vector(22680, 16),
34729 => conv_std_logic_vector(22815, 16),
34730 => conv_std_logic_vector(22950, 16),
34731 => conv_std_logic_vector(23085, 16),
34732 => conv_std_logic_vector(23220, 16),
34733 => conv_std_logic_vector(23355, 16),
34734 => conv_std_logic_vector(23490, 16),
34735 => conv_std_logic_vector(23625, 16),
34736 => conv_std_logic_vector(23760, 16),
34737 => conv_std_logic_vector(23895, 16),
34738 => conv_std_logic_vector(24030, 16),
34739 => conv_std_logic_vector(24165, 16),
34740 => conv_std_logic_vector(24300, 16),
34741 => conv_std_logic_vector(24435, 16),
34742 => conv_std_logic_vector(24570, 16),
34743 => conv_std_logic_vector(24705, 16),
34744 => conv_std_logic_vector(24840, 16),
34745 => conv_std_logic_vector(24975, 16),
34746 => conv_std_logic_vector(25110, 16),
34747 => conv_std_logic_vector(25245, 16),
34748 => conv_std_logic_vector(25380, 16),
34749 => conv_std_logic_vector(25515, 16),
34750 => conv_std_logic_vector(25650, 16),
34751 => conv_std_logic_vector(25785, 16),
34752 => conv_std_logic_vector(25920, 16),
34753 => conv_std_logic_vector(26055, 16),
34754 => conv_std_logic_vector(26190, 16),
34755 => conv_std_logic_vector(26325, 16),
34756 => conv_std_logic_vector(26460, 16),
34757 => conv_std_logic_vector(26595, 16),
34758 => conv_std_logic_vector(26730, 16),
34759 => conv_std_logic_vector(26865, 16),
34760 => conv_std_logic_vector(27000, 16),
34761 => conv_std_logic_vector(27135, 16),
34762 => conv_std_logic_vector(27270, 16),
34763 => conv_std_logic_vector(27405, 16),
34764 => conv_std_logic_vector(27540, 16),
34765 => conv_std_logic_vector(27675, 16),
34766 => conv_std_logic_vector(27810, 16),
34767 => conv_std_logic_vector(27945, 16),
34768 => conv_std_logic_vector(28080, 16),
34769 => conv_std_logic_vector(28215, 16),
34770 => conv_std_logic_vector(28350, 16),
34771 => conv_std_logic_vector(28485, 16),
34772 => conv_std_logic_vector(28620, 16),
34773 => conv_std_logic_vector(28755, 16),
34774 => conv_std_logic_vector(28890, 16),
34775 => conv_std_logic_vector(29025, 16),
34776 => conv_std_logic_vector(29160, 16),
34777 => conv_std_logic_vector(29295, 16),
34778 => conv_std_logic_vector(29430, 16),
34779 => conv_std_logic_vector(29565, 16),
34780 => conv_std_logic_vector(29700, 16),
34781 => conv_std_logic_vector(29835, 16),
34782 => conv_std_logic_vector(29970, 16),
34783 => conv_std_logic_vector(30105, 16),
34784 => conv_std_logic_vector(30240, 16),
34785 => conv_std_logic_vector(30375, 16),
34786 => conv_std_logic_vector(30510, 16),
34787 => conv_std_logic_vector(30645, 16),
34788 => conv_std_logic_vector(30780, 16),
34789 => conv_std_logic_vector(30915, 16),
34790 => conv_std_logic_vector(31050, 16),
34791 => conv_std_logic_vector(31185, 16),
34792 => conv_std_logic_vector(31320, 16),
34793 => conv_std_logic_vector(31455, 16),
34794 => conv_std_logic_vector(31590, 16),
34795 => conv_std_logic_vector(31725, 16),
34796 => conv_std_logic_vector(31860, 16),
34797 => conv_std_logic_vector(31995, 16),
34798 => conv_std_logic_vector(32130, 16),
34799 => conv_std_logic_vector(32265, 16),
34800 => conv_std_logic_vector(32400, 16),
34801 => conv_std_logic_vector(32535, 16),
34802 => conv_std_logic_vector(32670, 16),
34803 => conv_std_logic_vector(32805, 16),
34804 => conv_std_logic_vector(32940, 16),
34805 => conv_std_logic_vector(33075, 16),
34806 => conv_std_logic_vector(33210, 16),
34807 => conv_std_logic_vector(33345, 16),
34808 => conv_std_logic_vector(33480, 16),
34809 => conv_std_logic_vector(33615, 16),
34810 => conv_std_logic_vector(33750, 16),
34811 => conv_std_logic_vector(33885, 16),
34812 => conv_std_logic_vector(34020, 16),
34813 => conv_std_logic_vector(34155, 16),
34814 => conv_std_logic_vector(34290, 16),
34815 => conv_std_logic_vector(34425, 16),
34816 => conv_std_logic_vector(0, 16),
34817 => conv_std_logic_vector(136, 16),
34818 => conv_std_logic_vector(272, 16),
34819 => conv_std_logic_vector(408, 16),
34820 => conv_std_logic_vector(544, 16),
34821 => conv_std_logic_vector(680, 16),
34822 => conv_std_logic_vector(816, 16),
34823 => conv_std_logic_vector(952, 16),
34824 => conv_std_logic_vector(1088, 16),
34825 => conv_std_logic_vector(1224, 16),
34826 => conv_std_logic_vector(1360, 16),
34827 => conv_std_logic_vector(1496, 16),
34828 => conv_std_logic_vector(1632, 16),
34829 => conv_std_logic_vector(1768, 16),
34830 => conv_std_logic_vector(1904, 16),
34831 => conv_std_logic_vector(2040, 16),
34832 => conv_std_logic_vector(2176, 16),
34833 => conv_std_logic_vector(2312, 16),
34834 => conv_std_logic_vector(2448, 16),
34835 => conv_std_logic_vector(2584, 16),
34836 => conv_std_logic_vector(2720, 16),
34837 => conv_std_logic_vector(2856, 16),
34838 => conv_std_logic_vector(2992, 16),
34839 => conv_std_logic_vector(3128, 16),
34840 => conv_std_logic_vector(3264, 16),
34841 => conv_std_logic_vector(3400, 16),
34842 => conv_std_logic_vector(3536, 16),
34843 => conv_std_logic_vector(3672, 16),
34844 => conv_std_logic_vector(3808, 16),
34845 => conv_std_logic_vector(3944, 16),
34846 => conv_std_logic_vector(4080, 16),
34847 => conv_std_logic_vector(4216, 16),
34848 => conv_std_logic_vector(4352, 16),
34849 => conv_std_logic_vector(4488, 16),
34850 => conv_std_logic_vector(4624, 16),
34851 => conv_std_logic_vector(4760, 16),
34852 => conv_std_logic_vector(4896, 16),
34853 => conv_std_logic_vector(5032, 16),
34854 => conv_std_logic_vector(5168, 16),
34855 => conv_std_logic_vector(5304, 16),
34856 => conv_std_logic_vector(5440, 16),
34857 => conv_std_logic_vector(5576, 16),
34858 => conv_std_logic_vector(5712, 16),
34859 => conv_std_logic_vector(5848, 16),
34860 => conv_std_logic_vector(5984, 16),
34861 => conv_std_logic_vector(6120, 16),
34862 => conv_std_logic_vector(6256, 16),
34863 => conv_std_logic_vector(6392, 16),
34864 => conv_std_logic_vector(6528, 16),
34865 => conv_std_logic_vector(6664, 16),
34866 => conv_std_logic_vector(6800, 16),
34867 => conv_std_logic_vector(6936, 16),
34868 => conv_std_logic_vector(7072, 16),
34869 => conv_std_logic_vector(7208, 16),
34870 => conv_std_logic_vector(7344, 16),
34871 => conv_std_logic_vector(7480, 16),
34872 => conv_std_logic_vector(7616, 16),
34873 => conv_std_logic_vector(7752, 16),
34874 => conv_std_logic_vector(7888, 16),
34875 => conv_std_logic_vector(8024, 16),
34876 => conv_std_logic_vector(8160, 16),
34877 => conv_std_logic_vector(8296, 16),
34878 => conv_std_logic_vector(8432, 16),
34879 => conv_std_logic_vector(8568, 16),
34880 => conv_std_logic_vector(8704, 16),
34881 => conv_std_logic_vector(8840, 16),
34882 => conv_std_logic_vector(8976, 16),
34883 => conv_std_logic_vector(9112, 16),
34884 => conv_std_logic_vector(9248, 16),
34885 => conv_std_logic_vector(9384, 16),
34886 => conv_std_logic_vector(9520, 16),
34887 => conv_std_logic_vector(9656, 16),
34888 => conv_std_logic_vector(9792, 16),
34889 => conv_std_logic_vector(9928, 16),
34890 => conv_std_logic_vector(10064, 16),
34891 => conv_std_logic_vector(10200, 16),
34892 => conv_std_logic_vector(10336, 16),
34893 => conv_std_logic_vector(10472, 16),
34894 => conv_std_logic_vector(10608, 16),
34895 => conv_std_logic_vector(10744, 16),
34896 => conv_std_logic_vector(10880, 16),
34897 => conv_std_logic_vector(11016, 16),
34898 => conv_std_logic_vector(11152, 16),
34899 => conv_std_logic_vector(11288, 16),
34900 => conv_std_logic_vector(11424, 16),
34901 => conv_std_logic_vector(11560, 16),
34902 => conv_std_logic_vector(11696, 16),
34903 => conv_std_logic_vector(11832, 16),
34904 => conv_std_logic_vector(11968, 16),
34905 => conv_std_logic_vector(12104, 16),
34906 => conv_std_logic_vector(12240, 16),
34907 => conv_std_logic_vector(12376, 16),
34908 => conv_std_logic_vector(12512, 16),
34909 => conv_std_logic_vector(12648, 16),
34910 => conv_std_logic_vector(12784, 16),
34911 => conv_std_logic_vector(12920, 16),
34912 => conv_std_logic_vector(13056, 16),
34913 => conv_std_logic_vector(13192, 16),
34914 => conv_std_logic_vector(13328, 16),
34915 => conv_std_logic_vector(13464, 16),
34916 => conv_std_logic_vector(13600, 16),
34917 => conv_std_logic_vector(13736, 16),
34918 => conv_std_logic_vector(13872, 16),
34919 => conv_std_logic_vector(14008, 16),
34920 => conv_std_logic_vector(14144, 16),
34921 => conv_std_logic_vector(14280, 16),
34922 => conv_std_logic_vector(14416, 16),
34923 => conv_std_logic_vector(14552, 16),
34924 => conv_std_logic_vector(14688, 16),
34925 => conv_std_logic_vector(14824, 16),
34926 => conv_std_logic_vector(14960, 16),
34927 => conv_std_logic_vector(15096, 16),
34928 => conv_std_logic_vector(15232, 16),
34929 => conv_std_logic_vector(15368, 16),
34930 => conv_std_logic_vector(15504, 16),
34931 => conv_std_logic_vector(15640, 16),
34932 => conv_std_logic_vector(15776, 16),
34933 => conv_std_logic_vector(15912, 16),
34934 => conv_std_logic_vector(16048, 16),
34935 => conv_std_logic_vector(16184, 16),
34936 => conv_std_logic_vector(16320, 16),
34937 => conv_std_logic_vector(16456, 16),
34938 => conv_std_logic_vector(16592, 16),
34939 => conv_std_logic_vector(16728, 16),
34940 => conv_std_logic_vector(16864, 16),
34941 => conv_std_logic_vector(17000, 16),
34942 => conv_std_logic_vector(17136, 16),
34943 => conv_std_logic_vector(17272, 16),
34944 => conv_std_logic_vector(17408, 16),
34945 => conv_std_logic_vector(17544, 16),
34946 => conv_std_logic_vector(17680, 16),
34947 => conv_std_logic_vector(17816, 16),
34948 => conv_std_logic_vector(17952, 16),
34949 => conv_std_logic_vector(18088, 16),
34950 => conv_std_logic_vector(18224, 16),
34951 => conv_std_logic_vector(18360, 16),
34952 => conv_std_logic_vector(18496, 16),
34953 => conv_std_logic_vector(18632, 16),
34954 => conv_std_logic_vector(18768, 16),
34955 => conv_std_logic_vector(18904, 16),
34956 => conv_std_logic_vector(19040, 16),
34957 => conv_std_logic_vector(19176, 16),
34958 => conv_std_logic_vector(19312, 16),
34959 => conv_std_logic_vector(19448, 16),
34960 => conv_std_logic_vector(19584, 16),
34961 => conv_std_logic_vector(19720, 16),
34962 => conv_std_logic_vector(19856, 16),
34963 => conv_std_logic_vector(19992, 16),
34964 => conv_std_logic_vector(20128, 16),
34965 => conv_std_logic_vector(20264, 16),
34966 => conv_std_logic_vector(20400, 16),
34967 => conv_std_logic_vector(20536, 16),
34968 => conv_std_logic_vector(20672, 16),
34969 => conv_std_logic_vector(20808, 16),
34970 => conv_std_logic_vector(20944, 16),
34971 => conv_std_logic_vector(21080, 16),
34972 => conv_std_logic_vector(21216, 16),
34973 => conv_std_logic_vector(21352, 16),
34974 => conv_std_logic_vector(21488, 16),
34975 => conv_std_logic_vector(21624, 16),
34976 => conv_std_logic_vector(21760, 16),
34977 => conv_std_logic_vector(21896, 16),
34978 => conv_std_logic_vector(22032, 16),
34979 => conv_std_logic_vector(22168, 16),
34980 => conv_std_logic_vector(22304, 16),
34981 => conv_std_logic_vector(22440, 16),
34982 => conv_std_logic_vector(22576, 16),
34983 => conv_std_logic_vector(22712, 16),
34984 => conv_std_logic_vector(22848, 16),
34985 => conv_std_logic_vector(22984, 16),
34986 => conv_std_logic_vector(23120, 16),
34987 => conv_std_logic_vector(23256, 16),
34988 => conv_std_logic_vector(23392, 16),
34989 => conv_std_logic_vector(23528, 16),
34990 => conv_std_logic_vector(23664, 16),
34991 => conv_std_logic_vector(23800, 16),
34992 => conv_std_logic_vector(23936, 16),
34993 => conv_std_logic_vector(24072, 16),
34994 => conv_std_logic_vector(24208, 16),
34995 => conv_std_logic_vector(24344, 16),
34996 => conv_std_logic_vector(24480, 16),
34997 => conv_std_logic_vector(24616, 16),
34998 => conv_std_logic_vector(24752, 16),
34999 => conv_std_logic_vector(24888, 16),
35000 => conv_std_logic_vector(25024, 16),
35001 => conv_std_logic_vector(25160, 16),
35002 => conv_std_logic_vector(25296, 16),
35003 => conv_std_logic_vector(25432, 16),
35004 => conv_std_logic_vector(25568, 16),
35005 => conv_std_logic_vector(25704, 16),
35006 => conv_std_logic_vector(25840, 16),
35007 => conv_std_logic_vector(25976, 16),
35008 => conv_std_logic_vector(26112, 16),
35009 => conv_std_logic_vector(26248, 16),
35010 => conv_std_logic_vector(26384, 16),
35011 => conv_std_logic_vector(26520, 16),
35012 => conv_std_logic_vector(26656, 16),
35013 => conv_std_logic_vector(26792, 16),
35014 => conv_std_logic_vector(26928, 16),
35015 => conv_std_logic_vector(27064, 16),
35016 => conv_std_logic_vector(27200, 16),
35017 => conv_std_logic_vector(27336, 16),
35018 => conv_std_logic_vector(27472, 16),
35019 => conv_std_logic_vector(27608, 16),
35020 => conv_std_logic_vector(27744, 16),
35021 => conv_std_logic_vector(27880, 16),
35022 => conv_std_logic_vector(28016, 16),
35023 => conv_std_logic_vector(28152, 16),
35024 => conv_std_logic_vector(28288, 16),
35025 => conv_std_logic_vector(28424, 16),
35026 => conv_std_logic_vector(28560, 16),
35027 => conv_std_logic_vector(28696, 16),
35028 => conv_std_logic_vector(28832, 16),
35029 => conv_std_logic_vector(28968, 16),
35030 => conv_std_logic_vector(29104, 16),
35031 => conv_std_logic_vector(29240, 16),
35032 => conv_std_logic_vector(29376, 16),
35033 => conv_std_logic_vector(29512, 16),
35034 => conv_std_logic_vector(29648, 16),
35035 => conv_std_logic_vector(29784, 16),
35036 => conv_std_logic_vector(29920, 16),
35037 => conv_std_logic_vector(30056, 16),
35038 => conv_std_logic_vector(30192, 16),
35039 => conv_std_logic_vector(30328, 16),
35040 => conv_std_logic_vector(30464, 16),
35041 => conv_std_logic_vector(30600, 16),
35042 => conv_std_logic_vector(30736, 16),
35043 => conv_std_logic_vector(30872, 16),
35044 => conv_std_logic_vector(31008, 16),
35045 => conv_std_logic_vector(31144, 16),
35046 => conv_std_logic_vector(31280, 16),
35047 => conv_std_logic_vector(31416, 16),
35048 => conv_std_logic_vector(31552, 16),
35049 => conv_std_logic_vector(31688, 16),
35050 => conv_std_logic_vector(31824, 16),
35051 => conv_std_logic_vector(31960, 16),
35052 => conv_std_logic_vector(32096, 16),
35053 => conv_std_logic_vector(32232, 16),
35054 => conv_std_logic_vector(32368, 16),
35055 => conv_std_logic_vector(32504, 16),
35056 => conv_std_logic_vector(32640, 16),
35057 => conv_std_logic_vector(32776, 16),
35058 => conv_std_logic_vector(32912, 16),
35059 => conv_std_logic_vector(33048, 16),
35060 => conv_std_logic_vector(33184, 16),
35061 => conv_std_logic_vector(33320, 16),
35062 => conv_std_logic_vector(33456, 16),
35063 => conv_std_logic_vector(33592, 16),
35064 => conv_std_logic_vector(33728, 16),
35065 => conv_std_logic_vector(33864, 16),
35066 => conv_std_logic_vector(34000, 16),
35067 => conv_std_logic_vector(34136, 16),
35068 => conv_std_logic_vector(34272, 16),
35069 => conv_std_logic_vector(34408, 16),
35070 => conv_std_logic_vector(34544, 16),
35071 => conv_std_logic_vector(34680, 16),
35072 => conv_std_logic_vector(0, 16),
35073 => conv_std_logic_vector(137, 16),
35074 => conv_std_logic_vector(274, 16),
35075 => conv_std_logic_vector(411, 16),
35076 => conv_std_logic_vector(548, 16),
35077 => conv_std_logic_vector(685, 16),
35078 => conv_std_logic_vector(822, 16),
35079 => conv_std_logic_vector(959, 16),
35080 => conv_std_logic_vector(1096, 16),
35081 => conv_std_logic_vector(1233, 16),
35082 => conv_std_logic_vector(1370, 16),
35083 => conv_std_logic_vector(1507, 16),
35084 => conv_std_logic_vector(1644, 16),
35085 => conv_std_logic_vector(1781, 16),
35086 => conv_std_logic_vector(1918, 16),
35087 => conv_std_logic_vector(2055, 16),
35088 => conv_std_logic_vector(2192, 16),
35089 => conv_std_logic_vector(2329, 16),
35090 => conv_std_logic_vector(2466, 16),
35091 => conv_std_logic_vector(2603, 16),
35092 => conv_std_logic_vector(2740, 16),
35093 => conv_std_logic_vector(2877, 16),
35094 => conv_std_logic_vector(3014, 16),
35095 => conv_std_logic_vector(3151, 16),
35096 => conv_std_logic_vector(3288, 16),
35097 => conv_std_logic_vector(3425, 16),
35098 => conv_std_logic_vector(3562, 16),
35099 => conv_std_logic_vector(3699, 16),
35100 => conv_std_logic_vector(3836, 16),
35101 => conv_std_logic_vector(3973, 16),
35102 => conv_std_logic_vector(4110, 16),
35103 => conv_std_logic_vector(4247, 16),
35104 => conv_std_logic_vector(4384, 16),
35105 => conv_std_logic_vector(4521, 16),
35106 => conv_std_logic_vector(4658, 16),
35107 => conv_std_logic_vector(4795, 16),
35108 => conv_std_logic_vector(4932, 16),
35109 => conv_std_logic_vector(5069, 16),
35110 => conv_std_logic_vector(5206, 16),
35111 => conv_std_logic_vector(5343, 16),
35112 => conv_std_logic_vector(5480, 16),
35113 => conv_std_logic_vector(5617, 16),
35114 => conv_std_logic_vector(5754, 16),
35115 => conv_std_logic_vector(5891, 16),
35116 => conv_std_logic_vector(6028, 16),
35117 => conv_std_logic_vector(6165, 16),
35118 => conv_std_logic_vector(6302, 16),
35119 => conv_std_logic_vector(6439, 16),
35120 => conv_std_logic_vector(6576, 16),
35121 => conv_std_logic_vector(6713, 16),
35122 => conv_std_logic_vector(6850, 16),
35123 => conv_std_logic_vector(6987, 16),
35124 => conv_std_logic_vector(7124, 16),
35125 => conv_std_logic_vector(7261, 16),
35126 => conv_std_logic_vector(7398, 16),
35127 => conv_std_logic_vector(7535, 16),
35128 => conv_std_logic_vector(7672, 16),
35129 => conv_std_logic_vector(7809, 16),
35130 => conv_std_logic_vector(7946, 16),
35131 => conv_std_logic_vector(8083, 16),
35132 => conv_std_logic_vector(8220, 16),
35133 => conv_std_logic_vector(8357, 16),
35134 => conv_std_logic_vector(8494, 16),
35135 => conv_std_logic_vector(8631, 16),
35136 => conv_std_logic_vector(8768, 16),
35137 => conv_std_logic_vector(8905, 16),
35138 => conv_std_logic_vector(9042, 16),
35139 => conv_std_logic_vector(9179, 16),
35140 => conv_std_logic_vector(9316, 16),
35141 => conv_std_logic_vector(9453, 16),
35142 => conv_std_logic_vector(9590, 16),
35143 => conv_std_logic_vector(9727, 16),
35144 => conv_std_logic_vector(9864, 16),
35145 => conv_std_logic_vector(10001, 16),
35146 => conv_std_logic_vector(10138, 16),
35147 => conv_std_logic_vector(10275, 16),
35148 => conv_std_logic_vector(10412, 16),
35149 => conv_std_logic_vector(10549, 16),
35150 => conv_std_logic_vector(10686, 16),
35151 => conv_std_logic_vector(10823, 16),
35152 => conv_std_logic_vector(10960, 16),
35153 => conv_std_logic_vector(11097, 16),
35154 => conv_std_logic_vector(11234, 16),
35155 => conv_std_logic_vector(11371, 16),
35156 => conv_std_logic_vector(11508, 16),
35157 => conv_std_logic_vector(11645, 16),
35158 => conv_std_logic_vector(11782, 16),
35159 => conv_std_logic_vector(11919, 16),
35160 => conv_std_logic_vector(12056, 16),
35161 => conv_std_logic_vector(12193, 16),
35162 => conv_std_logic_vector(12330, 16),
35163 => conv_std_logic_vector(12467, 16),
35164 => conv_std_logic_vector(12604, 16),
35165 => conv_std_logic_vector(12741, 16),
35166 => conv_std_logic_vector(12878, 16),
35167 => conv_std_logic_vector(13015, 16),
35168 => conv_std_logic_vector(13152, 16),
35169 => conv_std_logic_vector(13289, 16),
35170 => conv_std_logic_vector(13426, 16),
35171 => conv_std_logic_vector(13563, 16),
35172 => conv_std_logic_vector(13700, 16),
35173 => conv_std_logic_vector(13837, 16),
35174 => conv_std_logic_vector(13974, 16),
35175 => conv_std_logic_vector(14111, 16),
35176 => conv_std_logic_vector(14248, 16),
35177 => conv_std_logic_vector(14385, 16),
35178 => conv_std_logic_vector(14522, 16),
35179 => conv_std_logic_vector(14659, 16),
35180 => conv_std_logic_vector(14796, 16),
35181 => conv_std_logic_vector(14933, 16),
35182 => conv_std_logic_vector(15070, 16),
35183 => conv_std_logic_vector(15207, 16),
35184 => conv_std_logic_vector(15344, 16),
35185 => conv_std_logic_vector(15481, 16),
35186 => conv_std_logic_vector(15618, 16),
35187 => conv_std_logic_vector(15755, 16),
35188 => conv_std_logic_vector(15892, 16),
35189 => conv_std_logic_vector(16029, 16),
35190 => conv_std_logic_vector(16166, 16),
35191 => conv_std_logic_vector(16303, 16),
35192 => conv_std_logic_vector(16440, 16),
35193 => conv_std_logic_vector(16577, 16),
35194 => conv_std_logic_vector(16714, 16),
35195 => conv_std_logic_vector(16851, 16),
35196 => conv_std_logic_vector(16988, 16),
35197 => conv_std_logic_vector(17125, 16),
35198 => conv_std_logic_vector(17262, 16),
35199 => conv_std_logic_vector(17399, 16),
35200 => conv_std_logic_vector(17536, 16),
35201 => conv_std_logic_vector(17673, 16),
35202 => conv_std_logic_vector(17810, 16),
35203 => conv_std_logic_vector(17947, 16),
35204 => conv_std_logic_vector(18084, 16),
35205 => conv_std_logic_vector(18221, 16),
35206 => conv_std_logic_vector(18358, 16),
35207 => conv_std_logic_vector(18495, 16),
35208 => conv_std_logic_vector(18632, 16),
35209 => conv_std_logic_vector(18769, 16),
35210 => conv_std_logic_vector(18906, 16),
35211 => conv_std_logic_vector(19043, 16),
35212 => conv_std_logic_vector(19180, 16),
35213 => conv_std_logic_vector(19317, 16),
35214 => conv_std_logic_vector(19454, 16),
35215 => conv_std_logic_vector(19591, 16),
35216 => conv_std_logic_vector(19728, 16),
35217 => conv_std_logic_vector(19865, 16),
35218 => conv_std_logic_vector(20002, 16),
35219 => conv_std_logic_vector(20139, 16),
35220 => conv_std_logic_vector(20276, 16),
35221 => conv_std_logic_vector(20413, 16),
35222 => conv_std_logic_vector(20550, 16),
35223 => conv_std_logic_vector(20687, 16),
35224 => conv_std_logic_vector(20824, 16),
35225 => conv_std_logic_vector(20961, 16),
35226 => conv_std_logic_vector(21098, 16),
35227 => conv_std_logic_vector(21235, 16),
35228 => conv_std_logic_vector(21372, 16),
35229 => conv_std_logic_vector(21509, 16),
35230 => conv_std_logic_vector(21646, 16),
35231 => conv_std_logic_vector(21783, 16),
35232 => conv_std_logic_vector(21920, 16),
35233 => conv_std_logic_vector(22057, 16),
35234 => conv_std_logic_vector(22194, 16),
35235 => conv_std_logic_vector(22331, 16),
35236 => conv_std_logic_vector(22468, 16),
35237 => conv_std_logic_vector(22605, 16),
35238 => conv_std_logic_vector(22742, 16),
35239 => conv_std_logic_vector(22879, 16),
35240 => conv_std_logic_vector(23016, 16),
35241 => conv_std_logic_vector(23153, 16),
35242 => conv_std_logic_vector(23290, 16),
35243 => conv_std_logic_vector(23427, 16),
35244 => conv_std_logic_vector(23564, 16),
35245 => conv_std_logic_vector(23701, 16),
35246 => conv_std_logic_vector(23838, 16),
35247 => conv_std_logic_vector(23975, 16),
35248 => conv_std_logic_vector(24112, 16),
35249 => conv_std_logic_vector(24249, 16),
35250 => conv_std_logic_vector(24386, 16),
35251 => conv_std_logic_vector(24523, 16),
35252 => conv_std_logic_vector(24660, 16),
35253 => conv_std_logic_vector(24797, 16),
35254 => conv_std_logic_vector(24934, 16),
35255 => conv_std_logic_vector(25071, 16),
35256 => conv_std_logic_vector(25208, 16),
35257 => conv_std_logic_vector(25345, 16),
35258 => conv_std_logic_vector(25482, 16),
35259 => conv_std_logic_vector(25619, 16),
35260 => conv_std_logic_vector(25756, 16),
35261 => conv_std_logic_vector(25893, 16),
35262 => conv_std_logic_vector(26030, 16),
35263 => conv_std_logic_vector(26167, 16),
35264 => conv_std_logic_vector(26304, 16),
35265 => conv_std_logic_vector(26441, 16),
35266 => conv_std_logic_vector(26578, 16),
35267 => conv_std_logic_vector(26715, 16),
35268 => conv_std_logic_vector(26852, 16),
35269 => conv_std_logic_vector(26989, 16),
35270 => conv_std_logic_vector(27126, 16),
35271 => conv_std_logic_vector(27263, 16),
35272 => conv_std_logic_vector(27400, 16),
35273 => conv_std_logic_vector(27537, 16),
35274 => conv_std_logic_vector(27674, 16),
35275 => conv_std_logic_vector(27811, 16),
35276 => conv_std_logic_vector(27948, 16),
35277 => conv_std_logic_vector(28085, 16),
35278 => conv_std_logic_vector(28222, 16),
35279 => conv_std_logic_vector(28359, 16),
35280 => conv_std_logic_vector(28496, 16),
35281 => conv_std_logic_vector(28633, 16),
35282 => conv_std_logic_vector(28770, 16),
35283 => conv_std_logic_vector(28907, 16),
35284 => conv_std_logic_vector(29044, 16),
35285 => conv_std_logic_vector(29181, 16),
35286 => conv_std_logic_vector(29318, 16),
35287 => conv_std_logic_vector(29455, 16),
35288 => conv_std_logic_vector(29592, 16),
35289 => conv_std_logic_vector(29729, 16),
35290 => conv_std_logic_vector(29866, 16),
35291 => conv_std_logic_vector(30003, 16),
35292 => conv_std_logic_vector(30140, 16),
35293 => conv_std_logic_vector(30277, 16),
35294 => conv_std_logic_vector(30414, 16),
35295 => conv_std_logic_vector(30551, 16),
35296 => conv_std_logic_vector(30688, 16),
35297 => conv_std_logic_vector(30825, 16),
35298 => conv_std_logic_vector(30962, 16),
35299 => conv_std_logic_vector(31099, 16),
35300 => conv_std_logic_vector(31236, 16),
35301 => conv_std_logic_vector(31373, 16),
35302 => conv_std_logic_vector(31510, 16),
35303 => conv_std_logic_vector(31647, 16),
35304 => conv_std_logic_vector(31784, 16),
35305 => conv_std_logic_vector(31921, 16),
35306 => conv_std_logic_vector(32058, 16),
35307 => conv_std_logic_vector(32195, 16),
35308 => conv_std_logic_vector(32332, 16),
35309 => conv_std_logic_vector(32469, 16),
35310 => conv_std_logic_vector(32606, 16),
35311 => conv_std_logic_vector(32743, 16),
35312 => conv_std_logic_vector(32880, 16),
35313 => conv_std_logic_vector(33017, 16),
35314 => conv_std_logic_vector(33154, 16),
35315 => conv_std_logic_vector(33291, 16),
35316 => conv_std_logic_vector(33428, 16),
35317 => conv_std_logic_vector(33565, 16),
35318 => conv_std_logic_vector(33702, 16),
35319 => conv_std_logic_vector(33839, 16),
35320 => conv_std_logic_vector(33976, 16),
35321 => conv_std_logic_vector(34113, 16),
35322 => conv_std_logic_vector(34250, 16),
35323 => conv_std_logic_vector(34387, 16),
35324 => conv_std_logic_vector(34524, 16),
35325 => conv_std_logic_vector(34661, 16),
35326 => conv_std_logic_vector(34798, 16),
35327 => conv_std_logic_vector(34935, 16),
35328 => conv_std_logic_vector(0, 16),
35329 => conv_std_logic_vector(138, 16),
35330 => conv_std_logic_vector(276, 16),
35331 => conv_std_logic_vector(414, 16),
35332 => conv_std_logic_vector(552, 16),
35333 => conv_std_logic_vector(690, 16),
35334 => conv_std_logic_vector(828, 16),
35335 => conv_std_logic_vector(966, 16),
35336 => conv_std_logic_vector(1104, 16),
35337 => conv_std_logic_vector(1242, 16),
35338 => conv_std_logic_vector(1380, 16),
35339 => conv_std_logic_vector(1518, 16),
35340 => conv_std_logic_vector(1656, 16),
35341 => conv_std_logic_vector(1794, 16),
35342 => conv_std_logic_vector(1932, 16),
35343 => conv_std_logic_vector(2070, 16),
35344 => conv_std_logic_vector(2208, 16),
35345 => conv_std_logic_vector(2346, 16),
35346 => conv_std_logic_vector(2484, 16),
35347 => conv_std_logic_vector(2622, 16),
35348 => conv_std_logic_vector(2760, 16),
35349 => conv_std_logic_vector(2898, 16),
35350 => conv_std_logic_vector(3036, 16),
35351 => conv_std_logic_vector(3174, 16),
35352 => conv_std_logic_vector(3312, 16),
35353 => conv_std_logic_vector(3450, 16),
35354 => conv_std_logic_vector(3588, 16),
35355 => conv_std_logic_vector(3726, 16),
35356 => conv_std_logic_vector(3864, 16),
35357 => conv_std_logic_vector(4002, 16),
35358 => conv_std_logic_vector(4140, 16),
35359 => conv_std_logic_vector(4278, 16),
35360 => conv_std_logic_vector(4416, 16),
35361 => conv_std_logic_vector(4554, 16),
35362 => conv_std_logic_vector(4692, 16),
35363 => conv_std_logic_vector(4830, 16),
35364 => conv_std_logic_vector(4968, 16),
35365 => conv_std_logic_vector(5106, 16),
35366 => conv_std_logic_vector(5244, 16),
35367 => conv_std_logic_vector(5382, 16),
35368 => conv_std_logic_vector(5520, 16),
35369 => conv_std_logic_vector(5658, 16),
35370 => conv_std_logic_vector(5796, 16),
35371 => conv_std_logic_vector(5934, 16),
35372 => conv_std_logic_vector(6072, 16),
35373 => conv_std_logic_vector(6210, 16),
35374 => conv_std_logic_vector(6348, 16),
35375 => conv_std_logic_vector(6486, 16),
35376 => conv_std_logic_vector(6624, 16),
35377 => conv_std_logic_vector(6762, 16),
35378 => conv_std_logic_vector(6900, 16),
35379 => conv_std_logic_vector(7038, 16),
35380 => conv_std_logic_vector(7176, 16),
35381 => conv_std_logic_vector(7314, 16),
35382 => conv_std_logic_vector(7452, 16),
35383 => conv_std_logic_vector(7590, 16),
35384 => conv_std_logic_vector(7728, 16),
35385 => conv_std_logic_vector(7866, 16),
35386 => conv_std_logic_vector(8004, 16),
35387 => conv_std_logic_vector(8142, 16),
35388 => conv_std_logic_vector(8280, 16),
35389 => conv_std_logic_vector(8418, 16),
35390 => conv_std_logic_vector(8556, 16),
35391 => conv_std_logic_vector(8694, 16),
35392 => conv_std_logic_vector(8832, 16),
35393 => conv_std_logic_vector(8970, 16),
35394 => conv_std_logic_vector(9108, 16),
35395 => conv_std_logic_vector(9246, 16),
35396 => conv_std_logic_vector(9384, 16),
35397 => conv_std_logic_vector(9522, 16),
35398 => conv_std_logic_vector(9660, 16),
35399 => conv_std_logic_vector(9798, 16),
35400 => conv_std_logic_vector(9936, 16),
35401 => conv_std_logic_vector(10074, 16),
35402 => conv_std_logic_vector(10212, 16),
35403 => conv_std_logic_vector(10350, 16),
35404 => conv_std_logic_vector(10488, 16),
35405 => conv_std_logic_vector(10626, 16),
35406 => conv_std_logic_vector(10764, 16),
35407 => conv_std_logic_vector(10902, 16),
35408 => conv_std_logic_vector(11040, 16),
35409 => conv_std_logic_vector(11178, 16),
35410 => conv_std_logic_vector(11316, 16),
35411 => conv_std_logic_vector(11454, 16),
35412 => conv_std_logic_vector(11592, 16),
35413 => conv_std_logic_vector(11730, 16),
35414 => conv_std_logic_vector(11868, 16),
35415 => conv_std_logic_vector(12006, 16),
35416 => conv_std_logic_vector(12144, 16),
35417 => conv_std_logic_vector(12282, 16),
35418 => conv_std_logic_vector(12420, 16),
35419 => conv_std_logic_vector(12558, 16),
35420 => conv_std_logic_vector(12696, 16),
35421 => conv_std_logic_vector(12834, 16),
35422 => conv_std_logic_vector(12972, 16),
35423 => conv_std_logic_vector(13110, 16),
35424 => conv_std_logic_vector(13248, 16),
35425 => conv_std_logic_vector(13386, 16),
35426 => conv_std_logic_vector(13524, 16),
35427 => conv_std_logic_vector(13662, 16),
35428 => conv_std_logic_vector(13800, 16),
35429 => conv_std_logic_vector(13938, 16),
35430 => conv_std_logic_vector(14076, 16),
35431 => conv_std_logic_vector(14214, 16),
35432 => conv_std_logic_vector(14352, 16),
35433 => conv_std_logic_vector(14490, 16),
35434 => conv_std_logic_vector(14628, 16),
35435 => conv_std_logic_vector(14766, 16),
35436 => conv_std_logic_vector(14904, 16),
35437 => conv_std_logic_vector(15042, 16),
35438 => conv_std_logic_vector(15180, 16),
35439 => conv_std_logic_vector(15318, 16),
35440 => conv_std_logic_vector(15456, 16),
35441 => conv_std_logic_vector(15594, 16),
35442 => conv_std_logic_vector(15732, 16),
35443 => conv_std_logic_vector(15870, 16),
35444 => conv_std_logic_vector(16008, 16),
35445 => conv_std_logic_vector(16146, 16),
35446 => conv_std_logic_vector(16284, 16),
35447 => conv_std_logic_vector(16422, 16),
35448 => conv_std_logic_vector(16560, 16),
35449 => conv_std_logic_vector(16698, 16),
35450 => conv_std_logic_vector(16836, 16),
35451 => conv_std_logic_vector(16974, 16),
35452 => conv_std_logic_vector(17112, 16),
35453 => conv_std_logic_vector(17250, 16),
35454 => conv_std_logic_vector(17388, 16),
35455 => conv_std_logic_vector(17526, 16),
35456 => conv_std_logic_vector(17664, 16),
35457 => conv_std_logic_vector(17802, 16),
35458 => conv_std_logic_vector(17940, 16),
35459 => conv_std_logic_vector(18078, 16),
35460 => conv_std_logic_vector(18216, 16),
35461 => conv_std_logic_vector(18354, 16),
35462 => conv_std_logic_vector(18492, 16),
35463 => conv_std_logic_vector(18630, 16),
35464 => conv_std_logic_vector(18768, 16),
35465 => conv_std_logic_vector(18906, 16),
35466 => conv_std_logic_vector(19044, 16),
35467 => conv_std_logic_vector(19182, 16),
35468 => conv_std_logic_vector(19320, 16),
35469 => conv_std_logic_vector(19458, 16),
35470 => conv_std_logic_vector(19596, 16),
35471 => conv_std_logic_vector(19734, 16),
35472 => conv_std_logic_vector(19872, 16),
35473 => conv_std_logic_vector(20010, 16),
35474 => conv_std_logic_vector(20148, 16),
35475 => conv_std_logic_vector(20286, 16),
35476 => conv_std_logic_vector(20424, 16),
35477 => conv_std_logic_vector(20562, 16),
35478 => conv_std_logic_vector(20700, 16),
35479 => conv_std_logic_vector(20838, 16),
35480 => conv_std_logic_vector(20976, 16),
35481 => conv_std_logic_vector(21114, 16),
35482 => conv_std_logic_vector(21252, 16),
35483 => conv_std_logic_vector(21390, 16),
35484 => conv_std_logic_vector(21528, 16),
35485 => conv_std_logic_vector(21666, 16),
35486 => conv_std_logic_vector(21804, 16),
35487 => conv_std_logic_vector(21942, 16),
35488 => conv_std_logic_vector(22080, 16),
35489 => conv_std_logic_vector(22218, 16),
35490 => conv_std_logic_vector(22356, 16),
35491 => conv_std_logic_vector(22494, 16),
35492 => conv_std_logic_vector(22632, 16),
35493 => conv_std_logic_vector(22770, 16),
35494 => conv_std_logic_vector(22908, 16),
35495 => conv_std_logic_vector(23046, 16),
35496 => conv_std_logic_vector(23184, 16),
35497 => conv_std_logic_vector(23322, 16),
35498 => conv_std_logic_vector(23460, 16),
35499 => conv_std_logic_vector(23598, 16),
35500 => conv_std_logic_vector(23736, 16),
35501 => conv_std_logic_vector(23874, 16),
35502 => conv_std_logic_vector(24012, 16),
35503 => conv_std_logic_vector(24150, 16),
35504 => conv_std_logic_vector(24288, 16),
35505 => conv_std_logic_vector(24426, 16),
35506 => conv_std_logic_vector(24564, 16),
35507 => conv_std_logic_vector(24702, 16),
35508 => conv_std_logic_vector(24840, 16),
35509 => conv_std_logic_vector(24978, 16),
35510 => conv_std_logic_vector(25116, 16),
35511 => conv_std_logic_vector(25254, 16),
35512 => conv_std_logic_vector(25392, 16),
35513 => conv_std_logic_vector(25530, 16),
35514 => conv_std_logic_vector(25668, 16),
35515 => conv_std_logic_vector(25806, 16),
35516 => conv_std_logic_vector(25944, 16),
35517 => conv_std_logic_vector(26082, 16),
35518 => conv_std_logic_vector(26220, 16),
35519 => conv_std_logic_vector(26358, 16),
35520 => conv_std_logic_vector(26496, 16),
35521 => conv_std_logic_vector(26634, 16),
35522 => conv_std_logic_vector(26772, 16),
35523 => conv_std_logic_vector(26910, 16),
35524 => conv_std_logic_vector(27048, 16),
35525 => conv_std_logic_vector(27186, 16),
35526 => conv_std_logic_vector(27324, 16),
35527 => conv_std_logic_vector(27462, 16),
35528 => conv_std_logic_vector(27600, 16),
35529 => conv_std_logic_vector(27738, 16),
35530 => conv_std_logic_vector(27876, 16),
35531 => conv_std_logic_vector(28014, 16),
35532 => conv_std_logic_vector(28152, 16),
35533 => conv_std_logic_vector(28290, 16),
35534 => conv_std_logic_vector(28428, 16),
35535 => conv_std_logic_vector(28566, 16),
35536 => conv_std_logic_vector(28704, 16),
35537 => conv_std_logic_vector(28842, 16),
35538 => conv_std_logic_vector(28980, 16),
35539 => conv_std_logic_vector(29118, 16),
35540 => conv_std_logic_vector(29256, 16),
35541 => conv_std_logic_vector(29394, 16),
35542 => conv_std_logic_vector(29532, 16),
35543 => conv_std_logic_vector(29670, 16),
35544 => conv_std_logic_vector(29808, 16),
35545 => conv_std_logic_vector(29946, 16),
35546 => conv_std_logic_vector(30084, 16),
35547 => conv_std_logic_vector(30222, 16),
35548 => conv_std_logic_vector(30360, 16),
35549 => conv_std_logic_vector(30498, 16),
35550 => conv_std_logic_vector(30636, 16),
35551 => conv_std_logic_vector(30774, 16),
35552 => conv_std_logic_vector(30912, 16),
35553 => conv_std_logic_vector(31050, 16),
35554 => conv_std_logic_vector(31188, 16),
35555 => conv_std_logic_vector(31326, 16),
35556 => conv_std_logic_vector(31464, 16),
35557 => conv_std_logic_vector(31602, 16),
35558 => conv_std_logic_vector(31740, 16),
35559 => conv_std_logic_vector(31878, 16),
35560 => conv_std_logic_vector(32016, 16),
35561 => conv_std_logic_vector(32154, 16),
35562 => conv_std_logic_vector(32292, 16),
35563 => conv_std_logic_vector(32430, 16),
35564 => conv_std_logic_vector(32568, 16),
35565 => conv_std_logic_vector(32706, 16),
35566 => conv_std_logic_vector(32844, 16),
35567 => conv_std_logic_vector(32982, 16),
35568 => conv_std_logic_vector(33120, 16),
35569 => conv_std_logic_vector(33258, 16),
35570 => conv_std_logic_vector(33396, 16),
35571 => conv_std_logic_vector(33534, 16),
35572 => conv_std_logic_vector(33672, 16),
35573 => conv_std_logic_vector(33810, 16),
35574 => conv_std_logic_vector(33948, 16),
35575 => conv_std_logic_vector(34086, 16),
35576 => conv_std_logic_vector(34224, 16),
35577 => conv_std_logic_vector(34362, 16),
35578 => conv_std_logic_vector(34500, 16),
35579 => conv_std_logic_vector(34638, 16),
35580 => conv_std_logic_vector(34776, 16),
35581 => conv_std_logic_vector(34914, 16),
35582 => conv_std_logic_vector(35052, 16),
35583 => conv_std_logic_vector(35190, 16),
35584 => conv_std_logic_vector(0, 16),
35585 => conv_std_logic_vector(139, 16),
35586 => conv_std_logic_vector(278, 16),
35587 => conv_std_logic_vector(417, 16),
35588 => conv_std_logic_vector(556, 16),
35589 => conv_std_logic_vector(695, 16),
35590 => conv_std_logic_vector(834, 16),
35591 => conv_std_logic_vector(973, 16),
35592 => conv_std_logic_vector(1112, 16),
35593 => conv_std_logic_vector(1251, 16),
35594 => conv_std_logic_vector(1390, 16),
35595 => conv_std_logic_vector(1529, 16),
35596 => conv_std_logic_vector(1668, 16),
35597 => conv_std_logic_vector(1807, 16),
35598 => conv_std_logic_vector(1946, 16),
35599 => conv_std_logic_vector(2085, 16),
35600 => conv_std_logic_vector(2224, 16),
35601 => conv_std_logic_vector(2363, 16),
35602 => conv_std_logic_vector(2502, 16),
35603 => conv_std_logic_vector(2641, 16),
35604 => conv_std_logic_vector(2780, 16),
35605 => conv_std_logic_vector(2919, 16),
35606 => conv_std_logic_vector(3058, 16),
35607 => conv_std_logic_vector(3197, 16),
35608 => conv_std_logic_vector(3336, 16),
35609 => conv_std_logic_vector(3475, 16),
35610 => conv_std_logic_vector(3614, 16),
35611 => conv_std_logic_vector(3753, 16),
35612 => conv_std_logic_vector(3892, 16),
35613 => conv_std_logic_vector(4031, 16),
35614 => conv_std_logic_vector(4170, 16),
35615 => conv_std_logic_vector(4309, 16),
35616 => conv_std_logic_vector(4448, 16),
35617 => conv_std_logic_vector(4587, 16),
35618 => conv_std_logic_vector(4726, 16),
35619 => conv_std_logic_vector(4865, 16),
35620 => conv_std_logic_vector(5004, 16),
35621 => conv_std_logic_vector(5143, 16),
35622 => conv_std_logic_vector(5282, 16),
35623 => conv_std_logic_vector(5421, 16),
35624 => conv_std_logic_vector(5560, 16),
35625 => conv_std_logic_vector(5699, 16),
35626 => conv_std_logic_vector(5838, 16),
35627 => conv_std_logic_vector(5977, 16),
35628 => conv_std_logic_vector(6116, 16),
35629 => conv_std_logic_vector(6255, 16),
35630 => conv_std_logic_vector(6394, 16),
35631 => conv_std_logic_vector(6533, 16),
35632 => conv_std_logic_vector(6672, 16),
35633 => conv_std_logic_vector(6811, 16),
35634 => conv_std_logic_vector(6950, 16),
35635 => conv_std_logic_vector(7089, 16),
35636 => conv_std_logic_vector(7228, 16),
35637 => conv_std_logic_vector(7367, 16),
35638 => conv_std_logic_vector(7506, 16),
35639 => conv_std_logic_vector(7645, 16),
35640 => conv_std_logic_vector(7784, 16),
35641 => conv_std_logic_vector(7923, 16),
35642 => conv_std_logic_vector(8062, 16),
35643 => conv_std_logic_vector(8201, 16),
35644 => conv_std_logic_vector(8340, 16),
35645 => conv_std_logic_vector(8479, 16),
35646 => conv_std_logic_vector(8618, 16),
35647 => conv_std_logic_vector(8757, 16),
35648 => conv_std_logic_vector(8896, 16),
35649 => conv_std_logic_vector(9035, 16),
35650 => conv_std_logic_vector(9174, 16),
35651 => conv_std_logic_vector(9313, 16),
35652 => conv_std_logic_vector(9452, 16),
35653 => conv_std_logic_vector(9591, 16),
35654 => conv_std_logic_vector(9730, 16),
35655 => conv_std_logic_vector(9869, 16),
35656 => conv_std_logic_vector(10008, 16),
35657 => conv_std_logic_vector(10147, 16),
35658 => conv_std_logic_vector(10286, 16),
35659 => conv_std_logic_vector(10425, 16),
35660 => conv_std_logic_vector(10564, 16),
35661 => conv_std_logic_vector(10703, 16),
35662 => conv_std_logic_vector(10842, 16),
35663 => conv_std_logic_vector(10981, 16),
35664 => conv_std_logic_vector(11120, 16),
35665 => conv_std_logic_vector(11259, 16),
35666 => conv_std_logic_vector(11398, 16),
35667 => conv_std_logic_vector(11537, 16),
35668 => conv_std_logic_vector(11676, 16),
35669 => conv_std_logic_vector(11815, 16),
35670 => conv_std_logic_vector(11954, 16),
35671 => conv_std_logic_vector(12093, 16),
35672 => conv_std_logic_vector(12232, 16),
35673 => conv_std_logic_vector(12371, 16),
35674 => conv_std_logic_vector(12510, 16),
35675 => conv_std_logic_vector(12649, 16),
35676 => conv_std_logic_vector(12788, 16),
35677 => conv_std_logic_vector(12927, 16),
35678 => conv_std_logic_vector(13066, 16),
35679 => conv_std_logic_vector(13205, 16),
35680 => conv_std_logic_vector(13344, 16),
35681 => conv_std_logic_vector(13483, 16),
35682 => conv_std_logic_vector(13622, 16),
35683 => conv_std_logic_vector(13761, 16),
35684 => conv_std_logic_vector(13900, 16),
35685 => conv_std_logic_vector(14039, 16),
35686 => conv_std_logic_vector(14178, 16),
35687 => conv_std_logic_vector(14317, 16),
35688 => conv_std_logic_vector(14456, 16),
35689 => conv_std_logic_vector(14595, 16),
35690 => conv_std_logic_vector(14734, 16),
35691 => conv_std_logic_vector(14873, 16),
35692 => conv_std_logic_vector(15012, 16),
35693 => conv_std_logic_vector(15151, 16),
35694 => conv_std_logic_vector(15290, 16),
35695 => conv_std_logic_vector(15429, 16),
35696 => conv_std_logic_vector(15568, 16),
35697 => conv_std_logic_vector(15707, 16),
35698 => conv_std_logic_vector(15846, 16),
35699 => conv_std_logic_vector(15985, 16),
35700 => conv_std_logic_vector(16124, 16),
35701 => conv_std_logic_vector(16263, 16),
35702 => conv_std_logic_vector(16402, 16),
35703 => conv_std_logic_vector(16541, 16),
35704 => conv_std_logic_vector(16680, 16),
35705 => conv_std_logic_vector(16819, 16),
35706 => conv_std_logic_vector(16958, 16),
35707 => conv_std_logic_vector(17097, 16),
35708 => conv_std_logic_vector(17236, 16),
35709 => conv_std_logic_vector(17375, 16),
35710 => conv_std_logic_vector(17514, 16),
35711 => conv_std_logic_vector(17653, 16),
35712 => conv_std_logic_vector(17792, 16),
35713 => conv_std_logic_vector(17931, 16),
35714 => conv_std_logic_vector(18070, 16),
35715 => conv_std_logic_vector(18209, 16),
35716 => conv_std_logic_vector(18348, 16),
35717 => conv_std_logic_vector(18487, 16),
35718 => conv_std_logic_vector(18626, 16),
35719 => conv_std_logic_vector(18765, 16),
35720 => conv_std_logic_vector(18904, 16),
35721 => conv_std_logic_vector(19043, 16),
35722 => conv_std_logic_vector(19182, 16),
35723 => conv_std_logic_vector(19321, 16),
35724 => conv_std_logic_vector(19460, 16),
35725 => conv_std_logic_vector(19599, 16),
35726 => conv_std_logic_vector(19738, 16),
35727 => conv_std_logic_vector(19877, 16),
35728 => conv_std_logic_vector(20016, 16),
35729 => conv_std_logic_vector(20155, 16),
35730 => conv_std_logic_vector(20294, 16),
35731 => conv_std_logic_vector(20433, 16),
35732 => conv_std_logic_vector(20572, 16),
35733 => conv_std_logic_vector(20711, 16),
35734 => conv_std_logic_vector(20850, 16),
35735 => conv_std_logic_vector(20989, 16),
35736 => conv_std_logic_vector(21128, 16),
35737 => conv_std_logic_vector(21267, 16),
35738 => conv_std_logic_vector(21406, 16),
35739 => conv_std_logic_vector(21545, 16),
35740 => conv_std_logic_vector(21684, 16),
35741 => conv_std_logic_vector(21823, 16),
35742 => conv_std_logic_vector(21962, 16),
35743 => conv_std_logic_vector(22101, 16),
35744 => conv_std_logic_vector(22240, 16),
35745 => conv_std_logic_vector(22379, 16),
35746 => conv_std_logic_vector(22518, 16),
35747 => conv_std_logic_vector(22657, 16),
35748 => conv_std_logic_vector(22796, 16),
35749 => conv_std_logic_vector(22935, 16),
35750 => conv_std_logic_vector(23074, 16),
35751 => conv_std_logic_vector(23213, 16),
35752 => conv_std_logic_vector(23352, 16),
35753 => conv_std_logic_vector(23491, 16),
35754 => conv_std_logic_vector(23630, 16),
35755 => conv_std_logic_vector(23769, 16),
35756 => conv_std_logic_vector(23908, 16),
35757 => conv_std_logic_vector(24047, 16),
35758 => conv_std_logic_vector(24186, 16),
35759 => conv_std_logic_vector(24325, 16),
35760 => conv_std_logic_vector(24464, 16),
35761 => conv_std_logic_vector(24603, 16),
35762 => conv_std_logic_vector(24742, 16),
35763 => conv_std_logic_vector(24881, 16),
35764 => conv_std_logic_vector(25020, 16),
35765 => conv_std_logic_vector(25159, 16),
35766 => conv_std_logic_vector(25298, 16),
35767 => conv_std_logic_vector(25437, 16),
35768 => conv_std_logic_vector(25576, 16),
35769 => conv_std_logic_vector(25715, 16),
35770 => conv_std_logic_vector(25854, 16),
35771 => conv_std_logic_vector(25993, 16),
35772 => conv_std_logic_vector(26132, 16),
35773 => conv_std_logic_vector(26271, 16),
35774 => conv_std_logic_vector(26410, 16),
35775 => conv_std_logic_vector(26549, 16),
35776 => conv_std_logic_vector(26688, 16),
35777 => conv_std_logic_vector(26827, 16),
35778 => conv_std_logic_vector(26966, 16),
35779 => conv_std_logic_vector(27105, 16),
35780 => conv_std_logic_vector(27244, 16),
35781 => conv_std_logic_vector(27383, 16),
35782 => conv_std_logic_vector(27522, 16),
35783 => conv_std_logic_vector(27661, 16),
35784 => conv_std_logic_vector(27800, 16),
35785 => conv_std_logic_vector(27939, 16),
35786 => conv_std_logic_vector(28078, 16),
35787 => conv_std_logic_vector(28217, 16),
35788 => conv_std_logic_vector(28356, 16),
35789 => conv_std_logic_vector(28495, 16),
35790 => conv_std_logic_vector(28634, 16),
35791 => conv_std_logic_vector(28773, 16),
35792 => conv_std_logic_vector(28912, 16),
35793 => conv_std_logic_vector(29051, 16),
35794 => conv_std_logic_vector(29190, 16),
35795 => conv_std_logic_vector(29329, 16),
35796 => conv_std_logic_vector(29468, 16),
35797 => conv_std_logic_vector(29607, 16),
35798 => conv_std_logic_vector(29746, 16),
35799 => conv_std_logic_vector(29885, 16),
35800 => conv_std_logic_vector(30024, 16),
35801 => conv_std_logic_vector(30163, 16),
35802 => conv_std_logic_vector(30302, 16),
35803 => conv_std_logic_vector(30441, 16),
35804 => conv_std_logic_vector(30580, 16),
35805 => conv_std_logic_vector(30719, 16),
35806 => conv_std_logic_vector(30858, 16),
35807 => conv_std_logic_vector(30997, 16),
35808 => conv_std_logic_vector(31136, 16),
35809 => conv_std_logic_vector(31275, 16),
35810 => conv_std_logic_vector(31414, 16),
35811 => conv_std_logic_vector(31553, 16),
35812 => conv_std_logic_vector(31692, 16),
35813 => conv_std_logic_vector(31831, 16),
35814 => conv_std_logic_vector(31970, 16),
35815 => conv_std_logic_vector(32109, 16),
35816 => conv_std_logic_vector(32248, 16),
35817 => conv_std_logic_vector(32387, 16),
35818 => conv_std_logic_vector(32526, 16),
35819 => conv_std_logic_vector(32665, 16),
35820 => conv_std_logic_vector(32804, 16),
35821 => conv_std_logic_vector(32943, 16),
35822 => conv_std_logic_vector(33082, 16),
35823 => conv_std_logic_vector(33221, 16),
35824 => conv_std_logic_vector(33360, 16),
35825 => conv_std_logic_vector(33499, 16),
35826 => conv_std_logic_vector(33638, 16),
35827 => conv_std_logic_vector(33777, 16),
35828 => conv_std_logic_vector(33916, 16),
35829 => conv_std_logic_vector(34055, 16),
35830 => conv_std_logic_vector(34194, 16),
35831 => conv_std_logic_vector(34333, 16),
35832 => conv_std_logic_vector(34472, 16),
35833 => conv_std_logic_vector(34611, 16),
35834 => conv_std_logic_vector(34750, 16),
35835 => conv_std_logic_vector(34889, 16),
35836 => conv_std_logic_vector(35028, 16),
35837 => conv_std_logic_vector(35167, 16),
35838 => conv_std_logic_vector(35306, 16),
35839 => conv_std_logic_vector(35445, 16),
35840 => conv_std_logic_vector(0, 16),
35841 => conv_std_logic_vector(140, 16),
35842 => conv_std_logic_vector(280, 16),
35843 => conv_std_logic_vector(420, 16),
35844 => conv_std_logic_vector(560, 16),
35845 => conv_std_logic_vector(700, 16),
35846 => conv_std_logic_vector(840, 16),
35847 => conv_std_logic_vector(980, 16),
35848 => conv_std_logic_vector(1120, 16),
35849 => conv_std_logic_vector(1260, 16),
35850 => conv_std_logic_vector(1400, 16),
35851 => conv_std_logic_vector(1540, 16),
35852 => conv_std_logic_vector(1680, 16),
35853 => conv_std_logic_vector(1820, 16),
35854 => conv_std_logic_vector(1960, 16),
35855 => conv_std_logic_vector(2100, 16),
35856 => conv_std_logic_vector(2240, 16),
35857 => conv_std_logic_vector(2380, 16),
35858 => conv_std_logic_vector(2520, 16),
35859 => conv_std_logic_vector(2660, 16),
35860 => conv_std_logic_vector(2800, 16),
35861 => conv_std_logic_vector(2940, 16),
35862 => conv_std_logic_vector(3080, 16),
35863 => conv_std_logic_vector(3220, 16),
35864 => conv_std_logic_vector(3360, 16),
35865 => conv_std_logic_vector(3500, 16),
35866 => conv_std_logic_vector(3640, 16),
35867 => conv_std_logic_vector(3780, 16),
35868 => conv_std_logic_vector(3920, 16),
35869 => conv_std_logic_vector(4060, 16),
35870 => conv_std_logic_vector(4200, 16),
35871 => conv_std_logic_vector(4340, 16),
35872 => conv_std_logic_vector(4480, 16),
35873 => conv_std_logic_vector(4620, 16),
35874 => conv_std_logic_vector(4760, 16),
35875 => conv_std_logic_vector(4900, 16),
35876 => conv_std_logic_vector(5040, 16),
35877 => conv_std_logic_vector(5180, 16),
35878 => conv_std_logic_vector(5320, 16),
35879 => conv_std_logic_vector(5460, 16),
35880 => conv_std_logic_vector(5600, 16),
35881 => conv_std_logic_vector(5740, 16),
35882 => conv_std_logic_vector(5880, 16),
35883 => conv_std_logic_vector(6020, 16),
35884 => conv_std_logic_vector(6160, 16),
35885 => conv_std_logic_vector(6300, 16),
35886 => conv_std_logic_vector(6440, 16),
35887 => conv_std_logic_vector(6580, 16),
35888 => conv_std_logic_vector(6720, 16),
35889 => conv_std_logic_vector(6860, 16),
35890 => conv_std_logic_vector(7000, 16),
35891 => conv_std_logic_vector(7140, 16),
35892 => conv_std_logic_vector(7280, 16),
35893 => conv_std_logic_vector(7420, 16),
35894 => conv_std_logic_vector(7560, 16),
35895 => conv_std_logic_vector(7700, 16),
35896 => conv_std_logic_vector(7840, 16),
35897 => conv_std_logic_vector(7980, 16),
35898 => conv_std_logic_vector(8120, 16),
35899 => conv_std_logic_vector(8260, 16),
35900 => conv_std_logic_vector(8400, 16),
35901 => conv_std_logic_vector(8540, 16),
35902 => conv_std_logic_vector(8680, 16),
35903 => conv_std_logic_vector(8820, 16),
35904 => conv_std_logic_vector(8960, 16),
35905 => conv_std_logic_vector(9100, 16),
35906 => conv_std_logic_vector(9240, 16),
35907 => conv_std_logic_vector(9380, 16),
35908 => conv_std_logic_vector(9520, 16),
35909 => conv_std_logic_vector(9660, 16),
35910 => conv_std_logic_vector(9800, 16),
35911 => conv_std_logic_vector(9940, 16),
35912 => conv_std_logic_vector(10080, 16),
35913 => conv_std_logic_vector(10220, 16),
35914 => conv_std_logic_vector(10360, 16),
35915 => conv_std_logic_vector(10500, 16),
35916 => conv_std_logic_vector(10640, 16),
35917 => conv_std_logic_vector(10780, 16),
35918 => conv_std_logic_vector(10920, 16),
35919 => conv_std_logic_vector(11060, 16),
35920 => conv_std_logic_vector(11200, 16),
35921 => conv_std_logic_vector(11340, 16),
35922 => conv_std_logic_vector(11480, 16),
35923 => conv_std_logic_vector(11620, 16),
35924 => conv_std_logic_vector(11760, 16),
35925 => conv_std_logic_vector(11900, 16),
35926 => conv_std_logic_vector(12040, 16),
35927 => conv_std_logic_vector(12180, 16),
35928 => conv_std_logic_vector(12320, 16),
35929 => conv_std_logic_vector(12460, 16),
35930 => conv_std_logic_vector(12600, 16),
35931 => conv_std_logic_vector(12740, 16),
35932 => conv_std_logic_vector(12880, 16),
35933 => conv_std_logic_vector(13020, 16),
35934 => conv_std_logic_vector(13160, 16),
35935 => conv_std_logic_vector(13300, 16),
35936 => conv_std_logic_vector(13440, 16),
35937 => conv_std_logic_vector(13580, 16),
35938 => conv_std_logic_vector(13720, 16),
35939 => conv_std_logic_vector(13860, 16),
35940 => conv_std_logic_vector(14000, 16),
35941 => conv_std_logic_vector(14140, 16),
35942 => conv_std_logic_vector(14280, 16),
35943 => conv_std_logic_vector(14420, 16),
35944 => conv_std_logic_vector(14560, 16),
35945 => conv_std_logic_vector(14700, 16),
35946 => conv_std_logic_vector(14840, 16),
35947 => conv_std_logic_vector(14980, 16),
35948 => conv_std_logic_vector(15120, 16),
35949 => conv_std_logic_vector(15260, 16),
35950 => conv_std_logic_vector(15400, 16),
35951 => conv_std_logic_vector(15540, 16),
35952 => conv_std_logic_vector(15680, 16),
35953 => conv_std_logic_vector(15820, 16),
35954 => conv_std_logic_vector(15960, 16),
35955 => conv_std_logic_vector(16100, 16),
35956 => conv_std_logic_vector(16240, 16),
35957 => conv_std_logic_vector(16380, 16),
35958 => conv_std_logic_vector(16520, 16),
35959 => conv_std_logic_vector(16660, 16),
35960 => conv_std_logic_vector(16800, 16),
35961 => conv_std_logic_vector(16940, 16),
35962 => conv_std_logic_vector(17080, 16),
35963 => conv_std_logic_vector(17220, 16),
35964 => conv_std_logic_vector(17360, 16),
35965 => conv_std_logic_vector(17500, 16),
35966 => conv_std_logic_vector(17640, 16),
35967 => conv_std_logic_vector(17780, 16),
35968 => conv_std_logic_vector(17920, 16),
35969 => conv_std_logic_vector(18060, 16),
35970 => conv_std_logic_vector(18200, 16),
35971 => conv_std_logic_vector(18340, 16),
35972 => conv_std_logic_vector(18480, 16),
35973 => conv_std_logic_vector(18620, 16),
35974 => conv_std_logic_vector(18760, 16),
35975 => conv_std_logic_vector(18900, 16),
35976 => conv_std_logic_vector(19040, 16),
35977 => conv_std_logic_vector(19180, 16),
35978 => conv_std_logic_vector(19320, 16),
35979 => conv_std_logic_vector(19460, 16),
35980 => conv_std_logic_vector(19600, 16),
35981 => conv_std_logic_vector(19740, 16),
35982 => conv_std_logic_vector(19880, 16),
35983 => conv_std_logic_vector(20020, 16),
35984 => conv_std_logic_vector(20160, 16),
35985 => conv_std_logic_vector(20300, 16),
35986 => conv_std_logic_vector(20440, 16),
35987 => conv_std_logic_vector(20580, 16),
35988 => conv_std_logic_vector(20720, 16),
35989 => conv_std_logic_vector(20860, 16),
35990 => conv_std_logic_vector(21000, 16),
35991 => conv_std_logic_vector(21140, 16),
35992 => conv_std_logic_vector(21280, 16),
35993 => conv_std_logic_vector(21420, 16),
35994 => conv_std_logic_vector(21560, 16),
35995 => conv_std_logic_vector(21700, 16),
35996 => conv_std_logic_vector(21840, 16),
35997 => conv_std_logic_vector(21980, 16),
35998 => conv_std_logic_vector(22120, 16),
35999 => conv_std_logic_vector(22260, 16),
36000 => conv_std_logic_vector(22400, 16),
36001 => conv_std_logic_vector(22540, 16),
36002 => conv_std_logic_vector(22680, 16),
36003 => conv_std_logic_vector(22820, 16),
36004 => conv_std_logic_vector(22960, 16),
36005 => conv_std_logic_vector(23100, 16),
36006 => conv_std_logic_vector(23240, 16),
36007 => conv_std_logic_vector(23380, 16),
36008 => conv_std_logic_vector(23520, 16),
36009 => conv_std_logic_vector(23660, 16),
36010 => conv_std_logic_vector(23800, 16),
36011 => conv_std_logic_vector(23940, 16),
36012 => conv_std_logic_vector(24080, 16),
36013 => conv_std_logic_vector(24220, 16),
36014 => conv_std_logic_vector(24360, 16),
36015 => conv_std_logic_vector(24500, 16),
36016 => conv_std_logic_vector(24640, 16),
36017 => conv_std_logic_vector(24780, 16),
36018 => conv_std_logic_vector(24920, 16),
36019 => conv_std_logic_vector(25060, 16),
36020 => conv_std_logic_vector(25200, 16),
36021 => conv_std_logic_vector(25340, 16),
36022 => conv_std_logic_vector(25480, 16),
36023 => conv_std_logic_vector(25620, 16),
36024 => conv_std_logic_vector(25760, 16),
36025 => conv_std_logic_vector(25900, 16),
36026 => conv_std_logic_vector(26040, 16),
36027 => conv_std_logic_vector(26180, 16),
36028 => conv_std_logic_vector(26320, 16),
36029 => conv_std_logic_vector(26460, 16),
36030 => conv_std_logic_vector(26600, 16),
36031 => conv_std_logic_vector(26740, 16),
36032 => conv_std_logic_vector(26880, 16),
36033 => conv_std_logic_vector(27020, 16),
36034 => conv_std_logic_vector(27160, 16),
36035 => conv_std_logic_vector(27300, 16),
36036 => conv_std_logic_vector(27440, 16),
36037 => conv_std_logic_vector(27580, 16),
36038 => conv_std_logic_vector(27720, 16),
36039 => conv_std_logic_vector(27860, 16),
36040 => conv_std_logic_vector(28000, 16),
36041 => conv_std_logic_vector(28140, 16),
36042 => conv_std_logic_vector(28280, 16),
36043 => conv_std_logic_vector(28420, 16),
36044 => conv_std_logic_vector(28560, 16),
36045 => conv_std_logic_vector(28700, 16),
36046 => conv_std_logic_vector(28840, 16),
36047 => conv_std_logic_vector(28980, 16),
36048 => conv_std_logic_vector(29120, 16),
36049 => conv_std_logic_vector(29260, 16),
36050 => conv_std_logic_vector(29400, 16),
36051 => conv_std_logic_vector(29540, 16),
36052 => conv_std_logic_vector(29680, 16),
36053 => conv_std_logic_vector(29820, 16),
36054 => conv_std_logic_vector(29960, 16),
36055 => conv_std_logic_vector(30100, 16),
36056 => conv_std_logic_vector(30240, 16),
36057 => conv_std_logic_vector(30380, 16),
36058 => conv_std_logic_vector(30520, 16),
36059 => conv_std_logic_vector(30660, 16),
36060 => conv_std_logic_vector(30800, 16),
36061 => conv_std_logic_vector(30940, 16),
36062 => conv_std_logic_vector(31080, 16),
36063 => conv_std_logic_vector(31220, 16),
36064 => conv_std_logic_vector(31360, 16),
36065 => conv_std_logic_vector(31500, 16),
36066 => conv_std_logic_vector(31640, 16),
36067 => conv_std_logic_vector(31780, 16),
36068 => conv_std_logic_vector(31920, 16),
36069 => conv_std_logic_vector(32060, 16),
36070 => conv_std_logic_vector(32200, 16),
36071 => conv_std_logic_vector(32340, 16),
36072 => conv_std_logic_vector(32480, 16),
36073 => conv_std_logic_vector(32620, 16),
36074 => conv_std_logic_vector(32760, 16),
36075 => conv_std_logic_vector(32900, 16),
36076 => conv_std_logic_vector(33040, 16),
36077 => conv_std_logic_vector(33180, 16),
36078 => conv_std_logic_vector(33320, 16),
36079 => conv_std_logic_vector(33460, 16),
36080 => conv_std_logic_vector(33600, 16),
36081 => conv_std_logic_vector(33740, 16),
36082 => conv_std_logic_vector(33880, 16),
36083 => conv_std_logic_vector(34020, 16),
36084 => conv_std_logic_vector(34160, 16),
36085 => conv_std_logic_vector(34300, 16),
36086 => conv_std_logic_vector(34440, 16),
36087 => conv_std_logic_vector(34580, 16),
36088 => conv_std_logic_vector(34720, 16),
36089 => conv_std_logic_vector(34860, 16),
36090 => conv_std_logic_vector(35000, 16),
36091 => conv_std_logic_vector(35140, 16),
36092 => conv_std_logic_vector(35280, 16),
36093 => conv_std_logic_vector(35420, 16),
36094 => conv_std_logic_vector(35560, 16),
36095 => conv_std_logic_vector(35700, 16),
36096 => conv_std_logic_vector(0, 16),
36097 => conv_std_logic_vector(141, 16),
36098 => conv_std_logic_vector(282, 16),
36099 => conv_std_logic_vector(423, 16),
36100 => conv_std_logic_vector(564, 16),
36101 => conv_std_logic_vector(705, 16),
36102 => conv_std_logic_vector(846, 16),
36103 => conv_std_logic_vector(987, 16),
36104 => conv_std_logic_vector(1128, 16),
36105 => conv_std_logic_vector(1269, 16),
36106 => conv_std_logic_vector(1410, 16),
36107 => conv_std_logic_vector(1551, 16),
36108 => conv_std_logic_vector(1692, 16),
36109 => conv_std_logic_vector(1833, 16),
36110 => conv_std_logic_vector(1974, 16),
36111 => conv_std_logic_vector(2115, 16),
36112 => conv_std_logic_vector(2256, 16),
36113 => conv_std_logic_vector(2397, 16),
36114 => conv_std_logic_vector(2538, 16),
36115 => conv_std_logic_vector(2679, 16),
36116 => conv_std_logic_vector(2820, 16),
36117 => conv_std_logic_vector(2961, 16),
36118 => conv_std_logic_vector(3102, 16),
36119 => conv_std_logic_vector(3243, 16),
36120 => conv_std_logic_vector(3384, 16),
36121 => conv_std_logic_vector(3525, 16),
36122 => conv_std_logic_vector(3666, 16),
36123 => conv_std_logic_vector(3807, 16),
36124 => conv_std_logic_vector(3948, 16),
36125 => conv_std_logic_vector(4089, 16),
36126 => conv_std_logic_vector(4230, 16),
36127 => conv_std_logic_vector(4371, 16),
36128 => conv_std_logic_vector(4512, 16),
36129 => conv_std_logic_vector(4653, 16),
36130 => conv_std_logic_vector(4794, 16),
36131 => conv_std_logic_vector(4935, 16),
36132 => conv_std_logic_vector(5076, 16),
36133 => conv_std_logic_vector(5217, 16),
36134 => conv_std_logic_vector(5358, 16),
36135 => conv_std_logic_vector(5499, 16),
36136 => conv_std_logic_vector(5640, 16),
36137 => conv_std_logic_vector(5781, 16),
36138 => conv_std_logic_vector(5922, 16),
36139 => conv_std_logic_vector(6063, 16),
36140 => conv_std_logic_vector(6204, 16),
36141 => conv_std_logic_vector(6345, 16),
36142 => conv_std_logic_vector(6486, 16),
36143 => conv_std_logic_vector(6627, 16),
36144 => conv_std_logic_vector(6768, 16),
36145 => conv_std_logic_vector(6909, 16),
36146 => conv_std_logic_vector(7050, 16),
36147 => conv_std_logic_vector(7191, 16),
36148 => conv_std_logic_vector(7332, 16),
36149 => conv_std_logic_vector(7473, 16),
36150 => conv_std_logic_vector(7614, 16),
36151 => conv_std_logic_vector(7755, 16),
36152 => conv_std_logic_vector(7896, 16),
36153 => conv_std_logic_vector(8037, 16),
36154 => conv_std_logic_vector(8178, 16),
36155 => conv_std_logic_vector(8319, 16),
36156 => conv_std_logic_vector(8460, 16),
36157 => conv_std_logic_vector(8601, 16),
36158 => conv_std_logic_vector(8742, 16),
36159 => conv_std_logic_vector(8883, 16),
36160 => conv_std_logic_vector(9024, 16),
36161 => conv_std_logic_vector(9165, 16),
36162 => conv_std_logic_vector(9306, 16),
36163 => conv_std_logic_vector(9447, 16),
36164 => conv_std_logic_vector(9588, 16),
36165 => conv_std_logic_vector(9729, 16),
36166 => conv_std_logic_vector(9870, 16),
36167 => conv_std_logic_vector(10011, 16),
36168 => conv_std_logic_vector(10152, 16),
36169 => conv_std_logic_vector(10293, 16),
36170 => conv_std_logic_vector(10434, 16),
36171 => conv_std_logic_vector(10575, 16),
36172 => conv_std_logic_vector(10716, 16),
36173 => conv_std_logic_vector(10857, 16),
36174 => conv_std_logic_vector(10998, 16),
36175 => conv_std_logic_vector(11139, 16),
36176 => conv_std_logic_vector(11280, 16),
36177 => conv_std_logic_vector(11421, 16),
36178 => conv_std_logic_vector(11562, 16),
36179 => conv_std_logic_vector(11703, 16),
36180 => conv_std_logic_vector(11844, 16),
36181 => conv_std_logic_vector(11985, 16),
36182 => conv_std_logic_vector(12126, 16),
36183 => conv_std_logic_vector(12267, 16),
36184 => conv_std_logic_vector(12408, 16),
36185 => conv_std_logic_vector(12549, 16),
36186 => conv_std_logic_vector(12690, 16),
36187 => conv_std_logic_vector(12831, 16),
36188 => conv_std_logic_vector(12972, 16),
36189 => conv_std_logic_vector(13113, 16),
36190 => conv_std_logic_vector(13254, 16),
36191 => conv_std_logic_vector(13395, 16),
36192 => conv_std_logic_vector(13536, 16),
36193 => conv_std_logic_vector(13677, 16),
36194 => conv_std_logic_vector(13818, 16),
36195 => conv_std_logic_vector(13959, 16),
36196 => conv_std_logic_vector(14100, 16),
36197 => conv_std_logic_vector(14241, 16),
36198 => conv_std_logic_vector(14382, 16),
36199 => conv_std_logic_vector(14523, 16),
36200 => conv_std_logic_vector(14664, 16),
36201 => conv_std_logic_vector(14805, 16),
36202 => conv_std_logic_vector(14946, 16),
36203 => conv_std_logic_vector(15087, 16),
36204 => conv_std_logic_vector(15228, 16),
36205 => conv_std_logic_vector(15369, 16),
36206 => conv_std_logic_vector(15510, 16),
36207 => conv_std_logic_vector(15651, 16),
36208 => conv_std_logic_vector(15792, 16),
36209 => conv_std_logic_vector(15933, 16),
36210 => conv_std_logic_vector(16074, 16),
36211 => conv_std_logic_vector(16215, 16),
36212 => conv_std_logic_vector(16356, 16),
36213 => conv_std_logic_vector(16497, 16),
36214 => conv_std_logic_vector(16638, 16),
36215 => conv_std_logic_vector(16779, 16),
36216 => conv_std_logic_vector(16920, 16),
36217 => conv_std_logic_vector(17061, 16),
36218 => conv_std_logic_vector(17202, 16),
36219 => conv_std_logic_vector(17343, 16),
36220 => conv_std_logic_vector(17484, 16),
36221 => conv_std_logic_vector(17625, 16),
36222 => conv_std_logic_vector(17766, 16),
36223 => conv_std_logic_vector(17907, 16),
36224 => conv_std_logic_vector(18048, 16),
36225 => conv_std_logic_vector(18189, 16),
36226 => conv_std_logic_vector(18330, 16),
36227 => conv_std_logic_vector(18471, 16),
36228 => conv_std_logic_vector(18612, 16),
36229 => conv_std_logic_vector(18753, 16),
36230 => conv_std_logic_vector(18894, 16),
36231 => conv_std_logic_vector(19035, 16),
36232 => conv_std_logic_vector(19176, 16),
36233 => conv_std_logic_vector(19317, 16),
36234 => conv_std_logic_vector(19458, 16),
36235 => conv_std_logic_vector(19599, 16),
36236 => conv_std_logic_vector(19740, 16),
36237 => conv_std_logic_vector(19881, 16),
36238 => conv_std_logic_vector(20022, 16),
36239 => conv_std_logic_vector(20163, 16),
36240 => conv_std_logic_vector(20304, 16),
36241 => conv_std_logic_vector(20445, 16),
36242 => conv_std_logic_vector(20586, 16),
36243 => conv_std_logic_vector(20727, 16),
36244 => conv_std_logic_vector(20868, 16),
36245 => conv_std_logic_vector(21009, 16),
36246 => conv_std_logic_vector(21150, 16),
36247 => conv_std_logic_vector(21291, 16),
36248 => conv_std_logic_vector(21432, 16),
36249 => conv_std_logic_vector(21573, 16),
36250 => conv_std_logic_vector(21714, 16),
36251 => conv_std_logic_vector(21855, 16),
36252 => conv_std_logic_vector(21996, 16),
36253 => conv_std_logic_vector(22137, 16),
36254 => conv_std_logic_vector(22278, 16),
36255 => conv_std_logic_vector(22419, 16),
36256 => conv_std_logic_vector(22560, 16),
36257 => conv_std_logic_vector(22701, 16),
36258 => conv_std_logic_vector(22842, 16),
36259 => conv_std_logic_vector(22983, 16),
36260 => conv_std_logic_vector(23124, 16),
36261 => conv_std_logic_vector(23265, 16),
36262 => conv_std_logic_vector(23406, 16),
36263 => conv_std_logic_vector(23547, 16),
36264 => conv_std_logic_vector(23688, 16),
36265 => conv_std_logic_vector(23829, 16),
36266 => conv_std_logic_vector(23970, 16),
36267 => conv_std_logic_vector(24111, 16),
36268 => conv_std_logic_vector(24252, 16),
36269 => conv_std_logic_vector(24393, 16),
36270 => conv_std_logic_vector(24534, 16),
36271 => conv_std_logic_vector(24675, 16),
36272 => conv_std_logic_vector(24816, 16),
36273 => conv_std_logic_vector(24957, 16),
36274 => conv_std_logic_vector(25098, 16),
36275 => conv_std_logic_vector(25239, 16),
36276 => conv_std_logic_vector(25380, 16),
36277 => conv_std_logic_vector(25521, 16),
36278 => conv_std_logic_vector(25662, 16),
36279 => conv_std_logic_vector(25803, 16),
36280 => conv_std_logic_vector(25944, 16),
36281 => conv_std_logic_vector(26085, 16),
36282 => conv_std_logic_vector(26226, 16),
36283 => conv_std_logic_vector(26367, 16),
36284 => conv_std_logic_vector(26508, 16),
36285 => conv_std_logic_vector(26649, 16),
36286 => conv_std_logic_vector(26790, 16),
36287 => conv_std_logic_vector(26931, 16),
36288 => conv_std_logic_vector(27072, 16),
36289 => conv_std_logic_vector(27213, 16),
36290 => conv_std_logic_vector(27354, 16),
36291 => conv_std_logic_vector(27495, 16),
36292 => conv_std_logic_vector(27636, 16),
36293 => conv_std_logic_vector(27777, 16),
36294 => conv_std_logic_vector(27918, 16),
36295 => conv_std_logic_vector(28059, 16),
36296 => conv_std_logic_vector(28200, 16),
36297 => conv_std_logic_vector(28341, 16),
36298 => conv_std_logic_vector(28482, 16),
36299 => conv_std_logic_vector(28623, 16),
36300 => conv_std_logic_vector(28764, 16),
36301 => conv_std_logic_vector(28905, 16),
36302 => conv_std_logic_vector(29046, 16),
36303 => conv_std_logic_vector(29187, 16),
36304 => conv_std_logic_vector(29328, 16),
36305 => conv_std_logic_vector(29469, 16),
36306 => conv_std_logic_vector(29610, 16),
36307 => conv_std_logic_vector(29751, 16),
36308 => conv_std_logic_vector(29892, 16),
36309 => conv_std_logic_vector(30033, 16),
36310 => conv_std_logic_vector(30174, 16),
36311 => conv_std_logic_vector(30315, 16),
36312 => conv_std_logic_vector(30456, 16),
36313 => conv_std_logic_vector(30597, 16),
36314 => conv_std_logic_vector(30738, 16),
36315 => conv_std_logic_vector(30879, 16),
36316 => conv_std_logic_vector(31020, 16),
36317 => conv_std_logic_vector(31161, 16),
36318 => conv_std_logic_vector(31302, 16),
36319 => conv_std_logic_vector(31443, 16),
36320 => conv_std_logic_vector(31584, 16),
36321 => conv_std_logic_vector(31725, 16),
36322 => conv_std_logic_vector(31866, 16),
36323 => conv_std_logic_vector(32007, 16),
36324 => conv_std_logic_vector(32148, 16),
36325 => conv_std_logic_vector(32289, 16),
36326 => conv_std_logic_vector(32430, 16),
36327 => conv_std_logic_vector(32571, 16),
36328 => conv_std_logic_vector(32712, 16),
36329 => conv_std_logic_vector(32853, 16),
36330 => conv_std_logic_vector(32994, 16),
36331 => conv_std_logic_vector(33135, 16),
36332 => conv_std_logic_vector(33276, 16),
36333 => conv_std_logic_vector(33417, 16),
36334 => conv_std_logic_vector(33558, 16),
36335 => conv_std_logic_vector(33699, 16),
36336 => conv_std_logic_vector(33840, 16),
36337 => conv_std_logic_vector(33981, 16),
36338 => conv_std_logic_vector(34122, 16),
36339 => conv_std_logic_vector(34263, 16),
36340 => conv_std_logic_vector(34404, 16),
36341 => conv_std_logic_vector(34545, 16),
36342 => conv_std_logic_vector(34686, 16),
36343 => conv_std_logic_vector(34827, 16),
36344 => conv_std_logic_vector(34968, 16),
36345 => conv_std_logic_vector(35109, 16),
36346 => conv_std_logic_vector(35250, 16),
36347 => conv_std_logic_vector(35391, 16),
36348 => conv_std_logic_vector(35532, 16),
36349 => conv_std_logic_vector(35673, 16),
36350 => conv_std_logic_vector(35814, 16),
36351 => conv_std_logic_vector(35955, 16),
36352 => conv_std_logic_vector(0, 16),
36353 => conv_std_logic_vector(142, 16),
36354 => conv_std_logic_vector(284, 16),
36355 => conv_std_logic_vector(426, 16),
36356 => conv_std_logic_vector(568, 16),
36357 => conv_std_logic_vector(710, 16),
36358 => conv_std_logic_vector(852, 16),
36359 => conv_std_logic_vector(994, 16),
36360 => conv_std_logic_vector(1136, 16),
36361 => conv_std_logic_vector(1278, 16),
36362 => conv_std_logic_vector(1420, 16),
36363 => conv_std_logic_vector(1562, 16),
36364 => conv_std_logic_vector(1704, 16),
36365 => conv_std_logic_vector(1846, 16),
36366 => conv_std_logic_vector(1988, 16),
36367 => conv_std_logic_vector(2130, 16),
36368 => conv_std_logic_vector(2272, 16),
36369 => conv_std_logic_vector(2414, 16),
36370 => conv_std_logic_vector(2556, 16),
36371 => conv_std_logic_vector(2698, 16),
36372 => conv_std_logic_vector(2840, 16),
36373 => conv_std_logic_vector(2982, 16),
36374 => conv_std_logic_vector(3124, 16),
36375 => conv_std_logic_vector(3266, 16),
36376 => conv_std_logic_vector(3408, 16),
36377 => conv_std_logic_vector(3550, 16),
36378 => conv_std_logic_vector(3692, 16),
36379 => conv_std_logic_vector(3834, 16),
36380 => conv_std_logic_vector(3976, 16),
36381 => conv_std_logic_vector(4118, 16),
36382 => conv_std_logic_vector(4260, 16),
36383 => conv_std_logic_vector(4402, 16),
36384 => conv_std_logic_vector(4544, 16),
36385 => conv_std_logic_vector(4686, 16),
36386 => conv_std_logic_vector(4828, 16),
36387 => conv_std_logic_vector(4970, 16),
36388 => conv_std_logic_vector(5112, 16),
36389 => conv_std_logic_vector(5254, 16),
36390 => conv_std_logic_vector(5396, 16),
36391 => conv_std_logic_vector(5538, 16),
36392 => conv_std_logic_vector(5680, 16),
36393 => conv_std_logic_vector(5822, 16),
36394 => conv_std_logic_vector(5964, 16),
36395 => conv_std_logic_vector(6106, 16),
36396 => conv_std_logic_vector(6248, 16),
36397 => conv_std_logic_vector(6390, 16),
36398 => conv_std_logic_vector(6532, 16),
36399 => conv_std_logic_vector(6674, 16),
36400 => conv_std_logic_vector(6816, 16),
36401 => conv_std_logic_vector(6958, 16),
36402 => conv_std_logic_vector(7100, 16),
36403 => conv_std_logic_vector(7242, 16),
36404 => conv_std_logic_vector(7384, 16),
36405 => conv_std_logic_vector(7526, 16),
36406 => conv_std_logic_vector(7668, 16),
36407 => conv_std_logic_vector(7810, 16),
36408 => conv_std_logic_vector(7952, 16),
36409 => conv_std_logic_vector(8094, 16),
36410 => conv_std_logic_vector(8236, 16),
36411 => conv_std_logic_vector(8378, 16),
36412 => conv_std_logic_vector(8520, 16),
36413 => conv_std_logic_vector(8662, 16),
36414 => conv_std_logic_vector(8804, 16),
36415 => conv_std_logic_vector(8946, 16),
36416 => conv_std_logic_vector(9088, 16),
36417 => conv_std_logic_vector(9230, 16),
36418 => conv_std_logic_vector(9372, 16),
36419 => conv_std_logic_vector(9514, 16),
36420 => conv_std_logic_vector(9656, 16),
36421 => conv_std_logic_vector(9798, 16),
36422 => conv_std_logic_vector(9940, 16),
36423 => conv_std_logic_vector(10082, 16),
36424 => conv_std_logic_vector(10224, 16),
36425 => conv_std_logic_vector(10366, 16),
36426 => conv_std_logic_vector(10508, 16),
36427 => conv_std_logic_vector(10650, 16),
36428 => conv_std_logic_vector(10792, 16),
36429 => conv_std_logic_vector(10934, 16),
36430 => conv_std_logic_vector(11076, 16),
36431 => conv_std_logic_vector(11218, 16),
36432 => conv_std_logic_vector(11360, 16),
36433 => conv_std_logic_vector(11502, 16),
36434 => conv_std_logic_vector(11644, 16),
36435 => conv_std_logic_vector(11786, 16),
36436 => conv_std_logic_vector(11928, 16),
36437 => conv_std_logic_vector(12070, 16),
36438 => conv_std_logic_vector(12212, 16),
36439 => conv_std_logic_vector(12354, 16),
36440 => conv_std_logic_vector(12496, 16),
36441 => conv_std_logic_vector(12638, 16),
36442 => conv_std_logic_vector(12780, 16),
36443 => conv_std_logic_vector(12922, 16),
36444 => conv_std_logic_vector(13064, 16),
36445 => conv_std_logic_vector(13206, 16),
36446 => conv_std_logic_vector(13348, 16),
36447 => conv_std_logic_vector(13490, 16),
36448 => conv_std_logic_vector(13632, 16),
36449 => conv_std_logic_vector(13774, 16),
36450 => conv_std_logic_vector(13916, 16),
36451 => conv_std_logic_vector(14058, 16),
36452 => conv_std_logic_vector(14200, 16),
36453 => conv_std_logic_vector(14342, 16),
36454 => conv_std_logic_vector(14484, 16),
36455 => conv_std_logic_vector(14626, 16),
36456 => conv_std_logic_vector(14768, 16),
36457 => conv_std_logic_vector(14910, 16),
36458 => conv_std_logic_vector(15052, 16),
36459 => conv_std_logic_vector(15194, 16),
36460 => conv_std_logic_vector(15336, 16),
36461 => conv_std_logic_vector(15478, 16),
36462 => conv_std_logic_vector(15620, 16),
36463 => conv_std_logic_vector(15762, 16),
36464 => conv_std_logic_vector(15904, 16),
36465 => conv_std_logic_vector(16046, 16),
36466 => conv_std_logic_vector(16188, 16),
36467 => conv_std_logic_vector(16330, 16),
36468 => conv_std_logic_vector(16472, 16),
36469 => conv_std_logic_vector(16614, 16),
36470 => conv_std_logic_vector(16756, 16),
36471 => conv_std_logic_vector(16898, 16),
36472 => conv_std_logic_vector(17040, 16),
36473 => conv_std_logic_vector(17182, 16),
36474 => conv_std_logic_vector(17324, 16),
36475 => conv_std_logic_vector(17466, 16),
36476 => conv_std_logic_vector(17608, 16),
36477 => conv_std_logic_vector(17750, 16),
36478 => conv_std_logic_vector(17892, 16),
36479 => conv_std_logic_vector(18034, 16),
36480 => conv_std_logic_vector(18176, 16),
36481 => conv_std_logic_vector(18318, 16),
36482 => conv_std_logic_vector(18460, 16),
36483 => conv_std_logic_vector(18602, 16),
36484 => conv_std_logic_vector(18744, 16),
36485 => conv_std_logic_vector(18886, 16),
36486 => conv_std_logic_vector(19028, 16),
36487 => conv_std_logic_vector(19170, 16),
36488 => conv_std_logic_vector(19312, 16),
36489 => conv_std_logic_vector(19454, 16),
36490 => conv_std_logic_vector(19596, 16),
36491 => conv_std_logic_vector(19738, 16),
36492 => conv_std_logic_vector(19880, 16),
36493 => conv_std_logic_vector(20022, 16),
36494 => conv_std_logic_vector(20164, 16),
36495 => conv_std_logic_vector(20306, 16),
36496 => conv_std_logic_vector(20448, 16),
36497 => conv_std_logic_vector(20590, 16),
36498 => conv_std_logic_vector(20732, 16),
36499 => conv_std_logic_vector(20874, 16),
36500 => conv_std_logic_vector(21016, 16),
36501 => conv_std_logic_vector(21158, 16),
36502 => conv_std_logic_vector(21300, 16),
36503 => conv_std_logic_vector(21442, 16),
36504 => conv_std_logic_vector(21584, 16),
36505 => conv_std_logic_vector(21726, 16),
36506 => conv_std_logic_vector(21868, 16),
36507 => conv_std_logic_vector(22010, 16),
36508 => conv_std_logic_vector(22152, 16),
36509 => conv_std_logic_vector(22294, 16),
36510 => conv_std_logic_vector(22436, 16),
36511 => conv_std_logic_vector(22578, 16),
36512 => conv_std_logic_vector(22720, 16),
36513 => conv_std_logic_vector(22862, 16),
36514 => conv_std_logic_vector(23004, 16),
36515 => conv_std_logic_vector(23146, 16),
36516 => conv_std_logic_vector(23288, 16),
36517 => conv_std_logic_vector(23430, 16),
36518 => conv_std_logic_vector(23572, 16),
36519 => conv_std_logic_vector(23714, 16),
36520 => conv_std_logic_vector(23856, 16),
36521 => conv_std_logic_vector(23998, 16),
36522 => conv_std_logic_vector(24140, 16),
36523 => conv_std_logic_vector(24282, 16),
36524 => conv_std_logic_vector(24424, 16),
36525 => conv_std_logic_vector(24566, 16),
36526 => conv_std_logic_vector(24708, 16),
36527 => conv_std_logic_vector(24850, 16),
36528 => conv_std_logic_vector(24992, 16),
36529 => conv_std_logic_vector(25134, 16),
36530 => conv_std_logic_vector(25276, 16),
36531 => conv_std_logic_vector(25418, 16),
36532 => conv_std_logic_vector(25560, 16),
36533 => conv_std_logic_vector(25702, 16),
36534 => conv_std_logic_vector(25844, 16),
36535 => conv_std_logic_vector(25986, 16),
36536 => conv_std_logic_vector(26128, 16),
36537 => conv_std_logic_vector(26270, 16),
36538 => conv_std_logic_vector(26412, 16),
36539 => conv_std_logic_vector(26554, 16),
36540 => conv_std_logic_vector(26696, 16),
36541 => conv_std_logic_vector(26838, 16),
36542 => conv_std_logic_vector(26980, 16),
36543 => conv_std_logic_vector(27122, 16),
36544 => conv_std_logic_vector(27264, 16),
36545 => conv_std_logic_vector(27406, 16),
36546 => conv_std_logic_vector(27548, 16),
36547 => conv_std_logic_vector(27690, 16),
36548 => conv_std_logic_vector(27832, 16),
36549 => conv_std_logic_vector(27974, 16),
36550 => conv_std_logic_vector(28116, 16),
36551 => conv_std_logic_vector(28258, 16),
36552 => conv_std_logic_vector(28400, 16),
36553 => conv_std_logic_vector(28542, 16),
36554 => conv_std_logic_vector(28684, 16),
36555 => conv_std_logic_vector(28826, 16),
36556 => conv_std_logic_vector(28968, 16),
36557 => conv_std_logic_vector(29110, 16),
36558 => conv_std_logic_vector(29252, 16),
36559 => conv_std_logic_vector(29394, 16),
36560 => conv_std_logic_vector(29536, 16),
36561 => conv_std_logic_vector(29678, 16),
36562 => conv_std_logic_vector(29820, 16),
36563 => conv_std_logic_vector(29962, 16),
36564 => conv_std_logic_vector(30104, 16),
36565 => conv_std_logic_vector(30246, 16),
36566 => conv_std_logic_vector(30388, 16),
36567 => conv_std_logic_vector(30530, 16),
36568 => conv_std_logic_vector(30672, 16),
36569 => conv_std_logic_vector(30814, 16),
36570 => conv_std_logic_vector(30956, 16),
36571 => conv_std_logic_vector(31098, 16),
36572 => conv_std_logic_vector(31240, 16),
36573 => conv_std_logic_vector(31382, 16),
36574 => conv_std_logic_vector(31524, 16),
36575 => conv_std_logic_vector(31666, 16),
36576 => conv_std_logic_vector(31808, 16),
36577 => conv_std_logic_vector(31950, 16),
36578 => conv_std_logic_vector(32092, 16),
36579 => conv_std_logic_vector(32234, 16),
36580 => conv_std_logic_vector(32376, 16),
36581 => conv_std_logic_vector(32518, 16),
36582 => conv_std_logic_vector(32660, 16),
36583 => conv_std_logic_vector(32802, 16),
36584 => conv_std_logic_vector(32944, 16),
36585 => conv_std_logic_vector(33086, 16),
36586 => conv_std_logic_vector(33228, 16),
36587 => conv_std_logic_vector(33370, 16),
36588 => conv_std_logic_vector(33512, 16),
36589 => conv_std_logic_vector(33654, 16),
36590 => conv_std_logic_vector(33796, 16),
36591 => conv_std_logic_vector(33938, 16),
36592 => conv_std_logic_vector(34080, 16),
36593 => conv_std_logic_vector(34222, 16),
36594 => conv_std_logic_vector(34364, 16),
36595 => conv_std_logic_vector(34506, 16),
36596 => conv_std_logic_vector(34648, 16),
36597 => conv_std_logic_vector(34790, 16),
36598 => conv_std_logic_vector(34932, 16),
36599 => conv_std_logic_vector(35074, 16),
36600 => conv_std_logic_vector(35216, 16),
36601 => conv_std_logic_vector(35358, 16),
36602 => conv_std_logic_vector(35500, 16),
36603 => conv_std_logic_vector(35642, 16),
36604 => conv_std_logic_vector(35784, 16),
36605 => conv_std_logic_vector(35926, 16),
36606 => conv_std_logic_vector(36068, 16),
36607 => conv_std_logic_vector(36210, 16),
36608 => conv_std_logic_vector(0, 16),
36609 => conv_std_logic_vector(143, 16),
36610 => conv_std_logic_vector(286, 16),
36611 => conv_std_logic_vector(429, 16),
36612 => conv_std_logic_vector(572, 16),
36613 => conv_std_logic_vector(715, 16),
36614 => conv_std_logic_vector(858, 16),
36615 => conv_std_logic_vector(1001, 16),
36616 => conv_std_logic_vector(1144, 16),
36617 => conv_std_logic_vector(1287, 16),
36618 => conv_std_logic_vector(1430, 16),
36619 => conv_std_logic_vector(1573, 16),
36620 => conv_std_logic_vector(1716, 16),
36621 => conv_std_logic_vector(1859, 16),
36622 => conv_std_logic_vector(2002, 16),
36623 => conv_std_logic_vector(2145, 16),
36624 => conv_std_logic_vector(2288, 16),
36625 => conv_std_logic_vector(2431, 16),
36626 => conv_std_logic_vector(2574, 16),
36627 => conv_std_logic_vector(2717, 16),
36628 => conv_std_logic_vector(2860, 16),
36629 => conv_std_logic_vector(3003, 16),
36630 => conv_std_logic_vector(3146, 16),
36631 => conv_std_logic_vector(3289, 16),
36632 => conv_std_logic_vector(3432, 16),
36633 => conv_std_logic_vector(3575, 16),
36634 => conv_std_logic_vector(3718, 16),
36635 => conv_std_logic_vector(3861, 16),
36636 => conv_std_logic_vector(4004, 16),
36637 => conv_std_logic_vector(4147, 16),
36638 => conv_std_logic_vector(4290, 16),
36639 => conv_std_logic_vector(4433, 16),
36640 => conv_std_logic_vector(4576, 16),
36641 => conv_std_logic_vector(4719, 16),
36642 => conv_std_logic_vector(4862, 16),
36643 => conv_std_logic_vector(5005, 16),
36644 => conv_std_logic_vector(5148, 16),
36645 => conv_std_logic_vector(5291, 16),
36646 => conv_std_logic_vector(5434, 16),
36647 => conv_std_logic_vector(5577, 16),
36648 => conv_std_logic_vector(5720, 16),
36649 => conv_std_logic_vector(5863, 16),
36650 => conv_std_logic_vector(6006, 16),
36651 => conv_std_logic_vector(6149, 16),
36652 => conv_std_logic_vector(6292, 16),
36653 => conv_std_logic_vector(6435, 16),
36654 => conv_std_logic_vector(6578, 16),
36655 => conv_std_logic_vector(6721, 16),
36656 => conv_std_logic_vector(6864, 16),
36657 => conv_std_logic_vector(7007, 16),
36658 => conv_std_logic_vector(7150, 16),
36659 => conv_std_logic_vector(7293, 16),
36660 => conv_std_logic_vector(7436, 16),
36661 => conv_std_logic_vector(7579, 16),
36662 => conv_std_logic_vector(7722, 16),
36663 => conv_std_logic_vector(7865, 16),
36664 => conv_std_logic_vector(8008, 16),
36665 => conv_std_logic_vector(8151, 16),
36666 => conv_std_logic_vector(8294, 16),
36667 => conv_std_logic_vector(8437, 16),
36668 => conv_std_logic_vector(8580, 16),
36669 => conv_std_logic_vector(8723, 16),
36670 => conv_std_logic_vector(8866, 16),
36671 => conv_std_logic_vector(9009, 16),
36672 => conv_std_logic_vector(9152, 16),
36673 => conv_std_logic_vector(9295, 16),
36674 => conv_std_logic_vector(9438, 16),
36675 => conv_std_logic_vector(9581, 16),
36676 => conv_std_logic_vector(9724, 16),
36677 => conv_std_logic_vector(9867, 16),
36678 => conv_std_logic_vector(10010, 16),
36679 => conv_std_logic_vector(10153, 16),
36680 => conv_std_logic_vector(10296, 16),
36681 => conv_std_logic_vector(10439, 16),
36682 => conv_std_logic_vector(10582, 16),
36683 => conv_std_logic_vector(10725, 16),
36684 => conv_std_logic_vector(10868, 16),
36685 => conv_std_logic_vector(11011, 16),
36686 => conv_std_logic_vector(11154, 16),
36687 => conv_std_logic_vector(11297, 16),
36688 => conv_std_logic_vector(11440, 16),
36689 => conv_std_logic_vector(11583, 16),
36690 => conv_std_logic_vector(11726, 16),
36691 => conv_std_logic_vector(11869, 16),
36692 => conv_std_logic_vector(12012, 16),
36693 => conv_std_logic_vector(12155, 16),
36694 => conv_std_logic_vector(12298, 16),
36695 => conv_std_logic_vector(12441, 16),
36696 => conv_std_logic_vector(12584, 16),
36697 => conv_std_logic_vector(12727, 16),
36698 => conv_std_logic_vector(12870, 16),
36699 => conv_std_logic_vector(13013, 16),
36700 => conv_std_logic_vector(13156, 16),
36701 => conv_std_logic_vector(13299, 16),
36702 => conv_std_logic_vector(13442, 16),
36703 => conv_std_logic_vector(13585, 16),
36704 => conv_std_logic_vector(13728, 16),
36705 => conv_std_logic_vector(13871, 16),
36706 => conv_std_logic_vector(14014, 16),
36707 => conv_std_logic_vector(14157, 16),
36708 => conv_std_logic_vector(14300, 16),
36709 => conv_std_logic_vector(14443, 16),
36710 => conv_std_logic_vector(14586, 16),
36711 => conv_std_logic_vector(14729, 16),
36712 => conv_std_logic_vector(14872, 16),
36713 => conv_std_logic_vector(15015, 16),
36714 => conv_std_logic_vector(15158, 16),
36715 => conv_std_logic_vector(15301, 16),
36716 => conv_std_logic_vector(15444, 16),
36717 => conv_std_logic_vector(15587, 16),
36718 => conv_std_logic_vector(15730, 16),
36719 => conv_std_logic_vector(15873, 16),
36720 => conv_std_logic_vector(16016, 16),
36721 => conv_std_logic_vector(16159, 16),
36722 => conv_std_logic_vector(16302, 16),
36723 => conv_std_logic_vector(16445, 16),
36724 => conv_std_logic_vector(16588, 16),
36725 => conv_std_logic_vector(16731, 16),
36726 => conv_std_logic_vector(16874, 16),
36727 => conv_std_logic_vector(17017, 16),
36728 => conv_std_logic_vector(17160, 16),
36729 => conv_std_logic_vector(17303, 16),
36730 => conv_std_logic_vector(17446, 16),
36731 => conv_std_logic_vector(17589, 16),
36732 => conv_std_logic_vector(17732, 16),
36733 => conv_std_logic_vector(17875, 16),
36734 => conv_std_logic_vector(18018, 16),
36735 => conv_std_logic_vector(18161, 16),
36736 => conv_std_logic_vector(18304, 16),
36737 => conv_std_logic_vector(18447, 16),
36738 => conv_std_logic_vector(18590, 16),
36739 => conv_std_logic_vector(18733, 16),
36740 => conv_std_logic_vector(18876, 16),
36741 => conv_std_logic_vector(19019, 16),
36742 => conv_std_logic_vector(19162, 16),
36743 => conv_std_logic_vector(19305, 16),
36744 => conv_std_logic_vector(19448, 16),
36745 => conv_std_logic_vector(19591, 16),
36746 => conv_std_logic_vector(19734, 16),
36747 => conv_std_logic_vector(19877, 16),
36748 => conv_std_logic_vector(20020, 16),
36749 => conv_std_logic_vector(20163, 16),
36750 => conv_std_logic_vector(20306, 16),
36751 => conv_std_logic_vector(20449, 16),
36752 => conv_std_logic_vector(20592, 16),
36753 => conv_std_logic_vector(20735, 16),
36754 => conv_std_logic_vector(20878, 16),
36755 => conv_std_logic_vector(21021, 16),
36756 => conv_std_logic_vector(21164, 16),
36757 => conv_std_logic_vector(21307, 16),
36758 => conv_std_logic_vector(21450, 16),
36759 => conv_std_logic_vector(21593, 16),
36760 => conv_std_logic_vector(21736, 16),
36761 => conv_std_logic_vector(21879, 16),
36762 => conv_std_logic_vector(22022, 16),
36763 => conv_std_logic_vector(22165, 16),
36764 => conv_std_logic_vector(22308, 16),
36765 => conv_std_logic_vector(22451, 16),
36766 => conv_std_logic_vector(22594, 16),
36767 => conv_std_logic_vector(22737, 16),
36768 => conv_std_logic_vector(22880, 16),
36769 => conv_std_logic_vector(23023, 16),
36770 => conv_std_logic_vector(23166, 16),
36771 => conv_std_logic_vector(23309, 16),
36772 => conv_std_logic_vector(23452, 16),
36773 => conv_std_logic_vector(23595, 16),
36774 => conv_std_logic_vector(23738, 16),
36775 => conv_std_logic_vector(23881, 16),
36776 => conv_std_logic_vector(24024, 16),
36777 => conv_std_logic_vector(24167, 16),
36778 => conv_std_logic_vector(24310, 16),
36779 => conv_std_logic_vector(24453, 16),
36780 => conv_std_logic_vector(24596, 16),
36781 => conv_std_logic_vector(24739, 16),
36782 => conv_std_logic_vector(24882, 16),
36783 => conv_std_logic_vector(25025, 16),
36784 => conv_std_logic_vector(25168, 16),
36785 => conv_std_logic_vector(25311, 16),
36786 => conv_std_logic_vector(25454, 16),
36787 => conv_std_logic_vector(25597, 16),
36788 => conv_std_logic_vector(25740, 16),
36789 => conv_std_logic_vector(25883, 16),
36790 => conv_std_logic_vector(26026, 16),
36791 => conv_std_logic_vector(26169, 16),
36792 => conv_std_logic_vector(26312, 16),
36793 => conv_std_logic_vector(26455, 16),
36794 => conv_std_logic_vector(26598, 16),
36795 => conv_std_logic_vector(26741, 16),
36796 => conv_std_logic_vector(26884, 16),
36797 => conv_std_logic_vector(27027, 16),
36798 => conv_std_logic_vector(27170, 16),
36799 => conv_std_logic_vector(27313, 16),
36800 => conv_std_logic_vector(27456, 16),
36801 => conv_std_logic_vector(27599, 16),
36802 => conv_std_logic_vector(27742, 16),
36803 => conv_std_logic_vector(27885, 16),
36804 => conv_std_logic_vector(28028, 16),
36805 => conv_std_logic_vector(28171, 16),
36806 => conv_std_logic_vector(28314, 16),
36807 => conv_std_logic_vector(28457, 16),
36808 => conv_std_logic_vector(28600, 16),
36809 => conv_std_logic_vector(28743, 16),
36810 => conv_std_logic_vector(28886, 16),
36811 => conv_std_logic_vector(29029, 16),
36812 => conv_std_logic_vector(29172, 16),
36813 => conv_std_logic_vector(29315, 16),
36814 => conv_std_logic_vector(29458, 16),
36815 => conv_std_logic_vector(29601, 16),
36816 => conv_std_logic_vector(29744, 16),
36817 => conv_std_logic_vector(29887, 16),
36818 => conv_std_logic_vector(30030, 16),
36819 => conv_std_logic_vector(30173, 16),
36820 => conv_std_logic_vector(30316, 16),
36821 => conv_std_logic_vector(30459, 16),
36822 => conv_std_logic_vector(30602, 16),
36823 => conv_std_logic_vector(30745, 16),
36824 => conv_std_logic_vector(30888, 16),
36825 => conv_std_logic_vector(31031, 16),
36826 => conv_std_logic_vector(31174, 16),
36827 => conv_std_logic_vector(31317, 16),
36828 => conv_std_logic_vector(31460, 16),
36829 => conv_std_logic_vector(31603, 16),
36830 => conv_std_logic_vector(31746, 16),
36831 => conv_std_logic_vector(31889, 16),
36832 => conv_std_logic_vector(32032, 16),
36833 => conv_std_logic_vector(32175, 16),
36834 => conv_std_logic_vector(32318, 16),
36835 => conv_std_logic_vector(32461, 16),
36836 => conv_std_logic_vector(32604, 16),
36837 => conv_std_logic_vector(32747, 16),
36838 => conv_std_logic_vector(32890, 16),
36839 => conv_std_logic_vector(33033, 16),
36840 => conv_std_logic_vector(33176, 16),
36841 => conv_std_logic_vector(33319, 16),
36842 => conv_std_logic_vector(33462, 16),
36843 => conv_std_logic_vector(33605, 16),
36844 => conv_std_logic_vector(33748, 16),
36845 => conv_std_logic_vector(33891, 16),
36846 => conv_std_logic_vector(34034, 16),
36847 => conv_std_logic_vector(34177, 16),
36848 => conv_std_logic_vector(34320, 16),
36849 => conv_std_logic_vector(34463, 16),
36850 => conv_std_logic_vector(34606, 16),
36851 => conv_std_logic_vector(34749, 16),
36852 => conv_std_logic_vector(34892, 16),
36853 => conv_std_logic_vector(35035, 16),
36854 => conv_std_logic_vector(35178, 16),
36855 => conv_std_logic_vector(35321, 16),
36856 => conv_std_logic_vector(35464, 16),
36857 => conv_std_logic_vector(35607, 16),
36858 => conv_std_logic_vector(35750, 16),
36859 => conv_std_logic_vector(35893, 16),
36860 => conv_std_logic_vector(36036, 16),
36861 => conv_std_logic_vector(36179, 16),
36862 => conv_std_logic_vector(36322, 16),
36863 => conv_std_logic_vector(36465, 16),
36864 => conv_std_logic_vector(0, 16),
36865 => conv_std_logic_vector(144, 16),
36866 => conv_std_logic_vector(288, 16),
36867 => conv_std_logic_vector(432, 16),
36868 => conv_std_logic_vector(576, 16),
36869 => conv_std_logic_vector(720, 16),
36870 => conv_std_logic_vector(864, 16),
36871 => conv_std_logic_vector(1008, 16),
36872 => conv_std_logic_vector(1152, 16),
36873 => conv_std_logic_vector(1296, 16),
36874 => conv_std_logic_vector(1440, 16),
36875 => conv_std_logic_vector(1584, 16),
36876 => conv_std_logic_vector(1728, 16),
36877 => conv_std_logic_vector(1872, 16),
36878 => conv_std_logic_vector(2016, 16),
36879 => conv_std_logic_vector(2160, 16),
36880 => conv_std_logic_vector(2304, 16),
36881 => conv_std_logic_vector(2448, 16),
36882 => conv_std_logic_vector(2592, 16),
36883 => conv_std_logic_vector(2736, 16),
36884 => conv_std_logic_vector(2880, 16),
36885 => conv_std_logic_vector(3024, 16),
36886 => conv_std_logic_vector(3168, 16),
36887 => conv_std_logic_vector(3312, 16),
36888 => conv_std_logic_vector(3456, 16),
36889 => conv_std_logic_vector(3600, 16),
36890 => conv_std_logic_vector(3744, 16),
36891 => conv_std_logic_vector(3888, 16),
36892 => conv_std_logic_vector(4032, 16),
36893 => conv_std_logic_vector(4176, 16),
36894 => conv_std_logic_vector(4320, 16),
36895 => conv_std_logic_vector(4464, 16),
36896 => conv_std_logic_vector(4608, 16),
36897 => conv_std_logic_vector(4752, 16),
36898 => conv_std_logic_vector(4896, 16),
36899 => conv_std_logic_vector(5040, 16),
36900 => conv_std_logic_vector(5184, 16),
36901 => conv_std_logic_vector(5328, 16),
36902 => conv_std_logic_vector(5472, 16),
36903 => conv_std_logic_vector(5616, 16),
36904 => conv_std_logic_vector(5760, 16),
36905 => conv_std_logic_vector(5904, 16),
36906 => conv_std_logic_vector(6048, 16),
36907 => conv_std_logic_vector(6192, 16),
36908 => conv_std_logic_vector(6336, 16),
36909 => conv_std_logic_vector(6480, 16),
36910 => conv_std_logic_vector(6624, 16),
36911 => conv_std_logic_vector(6768, 16),
36912 => conv_std_logic_vector(6912, 16),
36913 => conv_std_logic_vector(7056, 16),
36914 => conv_std_logic_vector(7200, 16),
36915 => conv_std_logic_vector(7344, 16),
36916 => conv_std_logic_vector(7488, 16),
36917 => conv_std_logic_vector(7632, 16),
36918 => conv_std_logic_vector(7776, 16),
36919 => conv_std_logic_vector(7920, 16),
36920 => conv_std_logic_vector(8064, 16),
36921 => conv_std_logic_vector(8208, 16),
36922 => conv_std_logic_vector(8352, 16),
36923 => conv_std_logic_vector(8496, 16),
36924 => conv_std_logic_vector(8640, 16),
36925 => conv_std_logic_vector(8784, 16),
36926 => conv_std_logic_vector(8928, 16),
36927 => conv_std_logic_vector(9072, 16),
36928 => conv_std_logic_vector(9216, 16),
36929 => conv_std_logic_vector(9360, 16),
36930 => conv_std_logic_vector(9504, 16),
36931 => conv_std_logic_vector(9648, 16),
36932 => conv_std_logic_vector(9792, 16),
36933 => conv_std_logic_vector(9936, 16),
36934 => conv_std_logic_vector(10080, 16),
36935 => conv_std_logic_vector(10224, 16),
36936 => conv_std_logic_vector(10368, 16),
36937 => conv_std_logic_vector(10512, 16),
36938 => conv_std_logic_vector(10656, 16),
36939 => conv_std_logic_vector(10800, 16),
36940 => conv_std_logic_vector(10944, 16),
36941 => conv_std_logic_vector(11088, 16),
36942 => conv_std_logic_vector(11232, 16),
36943 => conv_std_logic_vector(11376, 16),
36944 => conv_std_logic_vector(11520, 16),
36945 => conv_std_logic_vector(11664, 16),
36946 => conv_std_logic_vector(11808, 16),
36947 => conv_std_logic_vector(11952, 16),
36948 => conv_std_logic_vector(12096, 16),
36949 => conv_std_logic_vector(12240, 16),
36950 => conv_std_logic_vector(12384, 16),
36951 => conv_std_logic_vector(12528, 16),
36952 => conv_std_logic_vector(12672, 16),
36953 => conv_std_logic_vector(12816, 16),
36954 => conv_std_logic_vector(12960, 16),
36955 => conv_std_logic_vector(13104, 16),
36956 => conv_std_logic_vector(13248, 16),
36957 => conv_std_logic_vector(13392, 16),
36958 => conv_std_logic_vector(13536, 16),
36959 => conv_std_logic_vector(13680, 16),
36960 => conv_std_logic_vector(13824, 16),
36961 => conv_std_logic_vector(13968, 16),
36962 => conv_std_logic_vector(14112, 16),
36963 => conv_std_logic_vector(14256, 16),
36964 => conv_std_logic_vector(14400, 16),
36965 => conv_std_logic_vector(14544, 16),
36966 => conv_std_logic_vector(14688, 16),
36967 => conv_std_logic_vector(14832, 16),
36968 => conv_std_logic_vector(14976, 16),
36969 => conv_std_logic_vector(15120, 16),
36970 => conv_std_logic_vector(15264, 16),
36971 => conv_std_logic_vector(15408, 16),
36972 => conv_std_logic_vector(15552, 16),
36973 => conv_std_logic_vector(15696, 16),
36974 => conv_std_logic_vector(15840, 16),
36975 => conv_std_logic_vector(15984, 16),
36976 => conv_std_logic_vector(16128, 16),
36977 => conv_std_logic_vector(16272, 16),
36978 => conv_std_logic_vector(16416, 16),
36979 => conv_std_logic_vector(16560, 16),
36980 => conv_std_logic_vector(16704, 16),
36981 => conv_std_logic_vector(16848, 16),
36982 => conv_std_logic_vector(16992, 16),
36983 => conv_std_logic_vector(17136, 16),
36984 => conv_std_logic_vector(17280, 16),
36985 => conv_std_logic_vector(17424, 16),
36986 => conv_std_logic_vector(17568, 16),
36987 => conv_std_logic_vector(17712, 16),
36988 => conv_std_logic_vector(17856, 16),
36989 => conv_std_logic_vector(18000, 16),
36990 => conv_std_logic_vector(18144, 16),
36991 => conv_std_logic_vector(18288, 16),
36992 => conv_std_logic_vector(18432, 16),
36993 => conv_std_logic_vector(18576, 16),
36994 => conv_std_logic_vector(18720, 16),
36995 => conv_std_logic_vector(18864, 16),
36996 => conv_std_logic_vector(19008, 16),
36997 => conv_std_logic_vector(19152, 16),
36998 => conv_std_logic_vector(19296, 16),
36999 => conv_std_logic_vector(19440, 16),
37000 => conv_std_logic_vector(19584, 16),
37001 => conv_std_logic_vector(19728, 16),
37002 => conv_std_logic_vector(19872, 16),
37003 => conv_std_logic_vector(20016, 16),
37004 => conv_std_logic_vector(20160, 16),
37005 => conv_std_logic_vector(20304, 16),
37006 => conv_std_logic_vector(20448, 16),
37007 => conv_std_logic_vector(20592, 16),
37008 => conv_std_logic_vector(20736, 16),
37009 => conv_std_logic_vector(20880, 16),
37010 => conv_std_logic_vector(21024, 16),
37011 => conv_std_logic_vector(21168, 16),
37012 => conv_std_logic_vector(21312, 16),
37013 => conv_std_logic_vector(21456, 16),
37014 => conv_std_logic_vector(21600, 16),
37015 => conv_std_logic_vector(21744, 16),
37016 => conv_std_logic_vector(21888, 16),
37017 => conv_std_logic_vector(22032, 16),
37018 => conv_std_logic_vector(22176, 16),
37019 => conv_std_logic_vector(22320, 16),
37020 => conv_std_logic_vector(22464, 16),
37021 => conv_std_logic_vector(22608, 16),
37022 => conv_std_logic_vector(22752, 16),
37023 => conv_std_logic_vector(22896, 16),
37024 => conv_std_logic_vector(23040, 16),
37025 => conv_std_logic_vector(23184, 16),
37026 => conv_std_logic_vector(23328, 16),
37027 => conv_std_logic_vector(23472, 16),
37028 => conv_std_logic_vector(23616, 16),
37029 => conv_std_logic_vector(23760, 16),
37030 => conv_std_logic_vector(23904, 16),
37031 => conv_std_logic_vector(24048, 16),
37032 => conv_std_logic_vector(24192, 16),
37033 => conv_std_logic_vector(24336, 16),
37034 => conv_std_logic_vector(24480, 16),
37035 => conv_std_logic_vector(24624, 16),
37036 => conv_std_logic_vector(24768, 16),
37037 => conv_std_logic_vector(24912, 16),
37038 => conv_std_logic_vector(25056, 16),
37039 => conv_std_logic_vector(25200, 16),
37040 => conv_std_logic_vector(25344, 16),
37041 => conv_std_logic_vector(25488, 16),
37042 => conv_std_logic_vector(25632, 16),
37043 => conv_std_logic_vector(25776, 16),
37044 => conv_std_logic_vector(25920, 16),
37045 => conv_std_logic_vector(26064, 16),
37046 => conv_std_logic_vector(26208, 16),
37047 => conv_std_logic_vector(26352, 16),
37048 => conv_std_logic_vector(26496, 16),
37049 => conv_std_logic_vector(26640, 16),
37050 => conv_std_logic_vector(26784, 16),
37051 => conv_std_logic_vector(26928, 16),
37052 => conv_std_logic_vector(27072, 16),
37053 => conv_std_logic_vector(27216, 16),
37054 => conv_std_logic_vector(27360, 16),
37055 => conv_std_logic_vector(27504, 16),
37056 => conv_std_logic_vector(27648, 16),
37057 => conv_std_logic_vector(27792, 16),
37058 => conv_std_logic_vector(27936, 16),
37059 => conv_std_logic_vector(28080, 16),
37060 => conv_std_logic_vector(28224, 16),
37061 => conv_std_logic_vector(28368, 16),
37062 => conv_std_logic_vector(28512, 16),
37063 => conv_std_logic_vector(28656, 16),
37064 => conv_std_logic_vector(28800, 16),
37065 => conv_std_logic_vector(28944, 16),
37066 => conv_std_logic_vector(29088, 16),
37067 => conv_std_logic_vector(29232, 16),
37068 => conv_std_logic_vector(29376, 16),
37069 => conv_std_logic_vector(29520, 16),
37070 => conv_std_logic_vector(29664, 16),
37071 => conv_std_logic_vector(29808, 16),
37072 => conv_std_logic_vector(29952, 16),
37073 => conv_std_logic_vector(30096, 16),
37074 => conv_std_logic_vector(30240, 16),
37075 => conv_std_logic_vector(30384, 16),
37076 => conv_std_logic_vector(30528, 16),
37077 => conv_std_logic_vector(30672, 16),
37078 => conv_std_logic_vector(30816, 16),
37079 => conv_std_logic_vector(30960, 16),
37080 => conv_std_logic_vector(31104, 16),
37081 => conv_std_logic_vector(31248, 16),
37082 => conv_std_logic_vector(31392, 16),
37083 => conv_std_logic_vector(31536, 16),
37084 => conv_std_logic_vector(31680, 16),
37085 => conv_std_logic_vector(31824, 16),
37086 => conv_std_logic_vector(31968, 16),
37087 => conv_std_logic_vector(32112, 16),
37088 => conv_std_logic_vector(32256, 16),
37089 => conv_std_logic_vector(32400, 16),
37090 => conv_std_logic_vector(32544, 16),
37091 => conv_std_logic_vector(32688, 16),
37092 => conv_std_logic_vector(32832, 16),
37093 => conv_std_logic_vector(32976, 16),
37094 => conv_std_logic_vector(33120, 16),
37095 => conv_std_logic_vector(33264, 16),
37096 => conv_std_logic_vector(33408, 16),
37097 => conv_std_logic_vector(33552, 16),
37098 => conv_std_logic_vector(33696, 16),
37099 => conv_std_logic_vector(33840, 16),
37100 => conv_std_logic_vector(33984, 16),
37101 => conv_std_logic_vector(34128, 16),
37102 => conv_std_logic_vector(34272, 16),
37103 => conv_std_logic_vector(34416, 16),
37104 => conv_std_logic_vector(34560, 16),
37105 => conv_std_logic_vector(34704, 16),
37106 => conv_std_logic_vector(34848, 16),
37107 => conv_std_logic_vector(34992, 16),
37108 => conv_std_logic_vector(35136, 16),
37109 => conv_std_logic_vector(35280, 16),
37110 => conv_std_logic_vector(35424, 16),
37111 => conv_std_logic_vector(35568, 16),
37112 => conv_std_logic_vector(35712, 16),
37113 => conv_std_logic_vector(35856, 16),
37114 => conv_std_logic_vector(36000, 16),
37115 => conv_std_logic_vector(36144, 16),
37116 => conv_std_logic_vector(36288, 16),
37117 => conv_std_logic_vector(36432, 16),
37118 => conv_std_logic_vector(36576, 16),
37119 => conv_std_logic_vector(36720, 16),
37120 => conv_std_logic_vector(0, 16),
37121 => conv_std_logic_vector(145, 16),
37122 => conv_std_logic_vector(290, 16),
37123 => conv_std_logic_vector(435, 16),
37124 => conv_std_logic_vector(580, 16),
37125 => conv_std_logic_vector(725, 16),
37126 => conv_std_logic_vector(870, 16),
37127 => conv_std_logic_vector(1015, 16),
37128 => conv_std_logic_vector(1160, 16),
37129 => conv_std_logic_vector(1305, 16),
37130 => conv_std_logic_vector(1450, 16),
37131 => conv_std_logic_vector(1595, 16),
37132 => conv_std_logic_vector(1740, 16),
37133 => conv_std_logic_vector(1885, 16),
37134 => conv_std_logic_vector(2030, 16),
37135 => conv_std_logic_vector(2175, 16),
37136 => conv_std_logic_vector(2320, 16),
37137 => conv_std_logic_vector(2465, 16),
37138 => conv_std_logic_vector(2610, 16),
37139 => conv_std_logic_vector(2755, 16),
37140 => conv_std_logic_vector(2900, 16),
37141 => conv_std_logic_vector(3045, 16),
37142 => conv_std_logic_vector(3190, 16),
37143 => conv_std_logic_vector(3335, 16),
37144 => conv_std_logic_vector(3480, 16),
37145 => conv_std_logic_vector(3625, 16),
37146 => conv_std_logic_vector(3770, 16),
37147 => conv_std_logic_vector(3915, 16),
37148 => conv_std_logic_vector(4060, 16),
37149 => conv_std_logic_vector(4205, 16),
37150 => conv_std_logic_vector(4350, 16),
37151 => conv_std_logic_vector(4495, 16),
37152 => conv_std_logic_vector(4640, 16),
37153 => conv_std_logic_vector(4785, 16),
37154 => conv_std_logic_vector(4930, 16),
37155 => conv_std_logic_vector(5075, 16),
37156 => conv_std_logic_vector(5220, 16),
37157 => conv_std_logic_vector(5365, 16),
37158 => conv_std_logic_vector(5510, 16),
37159 => conv_std_logic_vector(5655, 16),
37160 => conv_std_logic_vector(5800, 16),
37161 => conv_std_logic_vector(5945, 16),
37162 => conv_std_logic_vector(6090, 16),
37163 => conv_std_logic_vector(6235, 16),
37164 => conv_std_logic_vector(6380, 16),
37165 => conv_std_logic_vector(6525, 16),
37166 => conv_std_logic_vector(6670, 16),
37167 => conv_std_logic_vector(6815, 16),
37168 => conv_std_logic_vector(6960, 16),
37169 => conv_std_logic_vector(7105, 16),
37170 => conv_std_logic_vector(7250, 16),
37171 => conv_std_logic_vector(7395, 16),
37172 => conv_std_logic_vector(7540, 16),
37173 => conv_std_logic_vector(7685, 16),
37174 => conv_std_logic_vector(7830, 16),
37175 => conv_std_logic_vector(7975, 16),
37176 => conv_std_logic_vector(8120, 16),
37177 => conv_std_logic_vector(8265, 16),
37178 => conv_std_logic_vector(8410, 16),
37179 => conv_std_logic_vector(8555, 16),
37180 => conv_std_logic_vector(8700, 16),
37181 => conv_std_logic_vector(8845, 16),
37182 => conv_std_logic_vector(8990, 16),
37183 => conv_std_logic_vector(9135, 16),
37184 => conv_std_logic_vector(9280, 16),
37185 => conv_std_logic_vector(9425, 16),
37186 => conv_std_logic_vector(9570, 16),
37187 => conv_std_logic_vector(9715, 16),
37188 => conv_std_logic_vector(9860, 16),
37189 => conv_std_logic_vector(10005, 16),
37190 => conv_std_logic_vector(10150, 16),
37191 => conv_std_logic_vector(10295, 16),
37192 => conv_std_logic_vector(10440, 16),
37193 => conv_std_logic_vector(10585, 16),
37194 => conv_std_logic_vector(10730, 16),
37195 => conv_std_logic_vector(10875, 16),
37196 => conv_std_logic_vector(11020, 16),
37197 => conv_std_logic_vector(11165, 16),
37198 => conv_std_logic_vector(11310, 16),
37199 => conv_std_logic_vector(11455, 16),
37200 => conv_std_logic_vector(11600, 16),
37201 => conv_std_logic_vector(11745, 16),
37202 => conv_std_logic_vector(11890, 16),
37203 => conv_std_logic_vector(12035, 16),
37204 => conv_std_logic_vector(12180, 16),
37205 => conv_std_logic_vector(12325, 16),
37206 => conv_std_logic_vector(12470, 16),
37207 => conv_std_logic_vector(12615, 16),
37208 => conv_std_logic_vector(12760, 16),
37209 => conv_std_logic_vector(12905, 16),
37210 => conv_std_logic_vector(13050, 16),
37211 => conv_std_logic_vector(13195, 16),
37212 => conv_std_logic_vector(13340, 16),
37213 => conv_std_logic_vector(13485, 16),
37214 => conv_std_logic_vector(13630, 16),
37215 => conv_std_logic_vector(13775, 16),
37216 => conv_std_logic_vector(13920, 16),
37217 => conv_std_logic_vector(14065, 16),
37218 => conv_std_logic_vector(14210, 16),
37219 => conv_std_logic_vector(14355, 16),
37220 => conv_std_logic_vector(14500, 16),
37221 => conv_std_logic_vector(14645, 16),
37222 => conv_std_logic_vector(14790, 16),
37223 => conv_std_logic_vector(14935, 16),
37224 => conv_std_logic_vector(15080, 16),
37225 => conv_std_logic_vector(15225, 16),
37226 => conv_std_logic_vector(15370, 16),
37227 => conv_std_logic_vector(15515, 16),
37228 => conv_std_logic_vector(15660, 16),
37229 => conv_std_logic_vector(15805, 16),
37230 => conv_std_logic_vector(15950, 16),
37231 => conv_std_logic_vector(16095, 16),
37232 => conv_std_logic_vector(16240, 16),
37233 => conv_std_logic_vector(16385, 16),
37234 => conv_std_logic_vector(16530, 16),
37235 => conv_std_logic_vector(16675, 16),
37236 => conv_std_logic_vector(16820, 16),
37237 => conv_std_logic_vector(16965, 16),
37238 => conv_std_logic_vector(17110, 16),
37239 => conv_std_logic_vector(17255, 16),
37240 => conv_std_logic_vector(17400, 16),
37241 => conv_std_logic_vector(17545, 16),
37242 => conv_std_logic_vector(17690, 16),
37243 => conv_std_logic_vector(17835, 16),
37244 => conv_std_logic_vector(17980, 16),
37245 => conv_std_logic_vector(18125, 16),
37246 => conv_std_logic_vector(18270, 16),
37247 => conv_std_logic_vector(18415, 16),
37248 => conv_std_logic_vector(18560, 16),
37249 => conv_std_logic_vector(18705, 16),
37250 => conv_std_logic_vector(18850, 16),
37251 => conv_std_logic_vector(18995, 16),
37252 => conv_std_logic_vector(19140, 16),
37253 => conv_std_logic_vector(19285, 16),
37254 => conv_std_logic_vector(19430, 16),
37255 => conv_std_logic_vector(19575, 16),
37256 => conv_std_logic_vector(19720, 16),
37257 => conv_std_logic_vector(19865, 16),
37258 => conv_std_logic_vector(20010, 16),
37259 => conv_std_logic_vector(20155, 16),
37260 => conv_std_logic_vector(20300, 16),
37261 => conv_std_logic_vector(20445, 16),
37262 => conv_std_logic_vector(20590, 16),
37263 => conv_std_logic_vector(20735, 16),
37264 => conv_std_logic_vector(20880, 16),
37265 => conv_std_logic_vector(21025, 16),
37266 => conv_std_logic_vector(21170, 16),
37267 => conv_std_logic_vector(21315, 16),
37268 => conv_std_logic_vector(21460, 16),
37269 => conv_std_logic_vector(21605, 16),
37270 => conv_std_logic_vector(21750, 16),
37271 => conv_std_logic_vector(21895, 16),
37272 => conv_std_logic_vector(22040, 16),
37273 => conv_std_logic_vector(22185, 16),
37274 => conv_std_logic_vector(22330, 16),
37275 => conv_std_logic_vector(22475, 16),
37276 => conv_std_logic_vector(22620, 16),
37277 => conv_std_logic_vector(22765, 16),
37278 => conv_std_logic_vector(22910, 16),
37279 => conv_std_logic_vector(23055, 16),
37280 => conv_std_logic_vector(23200, 16),
37281 => conv_std_logic_vector(23345, 16),
37282 => conv_std_logic_vector(23490, 16),
37283 => conv_std_logic_vector(23635, 16),
37284 => conv_std_logic_vector(23780, 16),
37285 => conv_std_logic_vector(23925, 16),
37286 => conv_std_logic_vector(24070, 16),
37287 => conv_std_logic_vector(24215, 16),
37288 => conv_std_logic_vector(24360, 16),
37289 => conv_std_logic_vector(24505, 16),
37290 => conv_std_logic_vector(24650, 16),
37291 => conv_std_logic_vector(24795, 16),
37292 => conv_std_logic_vector(24940, 16),
37293 => conv_std_logic_vector(25085, 16),
37294 => conv_std_logic_vector(25230, 16),
37295 => conv_std_logic_vector(25375, 16),
37296 => conv_std_logic_vector(25520, 16),
37297 => conv_std_logic_vector(25665, 16),
37298 => conv_std_logic_vector(25810, 16),
37299 => conv_std_logic_vector(25955, 16),
37300 => conv_std_logic_vector(26100, 16),
37301 => conv_std_logic_vector(26245, 16),
37302 => conv_std_logic_vector(26390, 16),
37303 => conv_std_logic_vector(26535, 16),
37304 => conv_std_logic_vector(26680, 16),
37305 => conv_std_logic_vector(26825, 16),
37306 => conv_std_logic_vector(26970, 16),
37307 => conv_std_logic_vector(27115, 16),
37308 => conv_std_logic_vector(27260, 16),
37309 => conv_std_logic_vector(27405, 16),
37310 => conv_std_logic_vector(27550, 16),
37311 => conv_std_logic_vector(27695, 16),
37312 => conv_std_logic_vector(27840, 16),
37313 => conv_std_logic_vector(27985, 16),
37314 => conv_std_logic_vector(28130, 16),
37315 => conv_std_logic_vector(28275, 16),
37316 => conv_std_logic_vector(28420, 16),
37317 => conv_std_logic_vector(28565, 16),
37318 => conv_std_logic_vector(28710, 16),
37319 => conv_std_logic_vector(28855, 16),
37320 => conv_std_logic_vector(29000, 16),
37321 => conv_std_logic_vector(29145, 16),
37322 => conv_std_logic_vector(29290, 16),
37323 => conv_std_logic_vector(29435, 16),
37324 => conv_std_logic_vector(29580, 16),
37325 => conv_std_logic_vector(29725, 16),
37326 => conv_std_logic_vector(29870, 16),
37327 => conv_std_logic_vector(30015, 16),
37328 => conv_std_logic_vector(30160, 16),
37329 => conv_std_logic_vector(30305, 16),
37330 => conv_std_logic_vector(30450, 16),
37331 => conv_std_logic_vector(30595, 16),
37332 => conv_std_logic_vector(30740, 16),
37333 => conv_std_logic_vector(30885, 16),
37334 => conv_std_logic_vector(31030, 16),
37335 => conv_std_logic_vector(31175, 16),
37336 => conv_std_logic_vector(31320, 16),
37337 => conv_std_logic_vector(31465, 16),
37338 => conv_std_logic_vector(31610, 16),
37339 => conv_std_logic_vector(31755, 16),
37340 => conv_std_logic_vector(31900, 16),
37341 => conv_std_logic_vector(32045, 16),
37342 => conv_std_logic_vector(32190, 16),
37343 => conv_std_logic_vector(32335, 16),
37344 => conv_std_logic_vector(32480, 16),
37345 => conv_std_logic_vector(32625, 16),
37346 => conv_std_logic_vector(32770, 16),
37347 => conv_std_logic_vector(32915, 16),
37348 => conv_std_logic_vector(33060, 16),
37349 => conv_std_logic_vector(33205, 16),
37350 => conv_std_logic_vector(33350, 16),
37351 => conv_std_logic_vector(33495, 16),
37352 => conv_std_logic_vector(33640, 16),
37353 => conv_std_logic_vector(33785, 16),
37354 => conv_std_logic_vector(33930, 16),
37355 => conv_std_logic_vector(34075, 16),
37356 => conv_std_logic_vector(34220, 16),
37357 => conv_std_logic_vector(34365, 16),
37358 => conv_std_logic_vector(34510, 16),
37359 => conv_std_logic_vector(34655, 16),
37360 => conv_std_logic_vector(34800, 16),
37361 => conv_std_logic_vector(34945, 16),
37362 => conv_std_logic_vector(35090, 16),
37363 => conv_std_logic_vector(35235, 16),
37364 => conv_std_logic_vector(35380, 16),
37365 => conv_std_logic_vector(35525, 16),
37366 => conv_std_logic_vector(35670, 16),
37367 => conv_std_logic_vector(35815, 16),
37368 => conv_std_logic_vector(35960, 16),
37369 => conv_std_logic_vector(36105, 16),
37370 => conv_std_logic_vector(36250, 16),
37371 => conv_std_logic_vector(36395, 16),
37372 => conv_std_logic_vector(36540, 16),
37373 => conv_std_logic_vector(36685, 16),
37374 => conv_std_logic_vector(36830, 16),
37375 => conv_std_logic_vector(36975, 16),
37376 => conv_std_logic_vector(0, 16),
37377 => conv_std_logic_vector(146, 16),
37378 => conv_std_logic_vector(292, 16),
37379 => conv_std_logic_vector(438, 16),
37380 => conv_std_logic_vector(584, 16),
37381 => conv_std_logic_vector(730, 16),
37382 => conv_std_logic_vector(876, 16),
37383 => conv_std_logic_vector(1022, 16),
37384 => conv_std_logic_vector(1168, 16),
37385 => conv_std_logic_vector(1314, 16),
37386 => conv_std_logic_vector(1460, 16),
37387 => conv_std_logic_vector(1606, 16),
37388 => conv_std_logic_vector(1752, 16),
37389 => conv_std_logic_vector(1898, 16),
37390 => conv_std_logic_vector(2044, 16),
37391 => conv_std_logic_vector(2190, 16),
37392 => conv_std_logic_vector(2336, 16),
37393 => conv_std_logic_vector(2482, 16),
37394 => conv_std_logic_vector(2628, 16),
37395 => conv_std_logic_vector(2774, 16),
37396 => conv_std_logic_vector(2920, 16),
37397 => conv_std_logic_vector(3066, 16),
37398 => conv_std_logic_vector(3212, 16),
37399 => conv_std_logic_vector(3358, 16),
37400 => conv_std_logic_vector(3504, 16),
37401 => conv_std_logic_vector(3650, 16),
37402 => conv_std_logic_vector(3796, 16),
37403 => conv_std_logic_vector(3942, 16),
37404 => conv_std_logic_vector(4088, 16),
37405 => conv_std_logic_vector(4234, 16),
37406 => conv_std_logic_vector(4380, 16),
37407 => conv_std_logic_vector(4526, 16),
37408 => conv_std_logic_vector(4672, 16),
37409 => conv_std_logic_vector(4818, 16),
37410 => conv_std_logic_vector(4964, 16),
37411 => conv_std_logic_vector(5110, 16),
37412 => conv_std_logic_vector(5256, 16),
37413 => conv_std_logic_vector(5402, 16),
37414 => conv_std_logic_vector(5548, 16),
37415 => conv_std_logic_vector(5694, 16),
37416 => conv_std_logic_vector(5840, 16),
37417 => conv_std_logic_vector(5986, 16),
37418 => conv_std_logic_vector(6132, 16),
37419 => conv_std_logic_vector(6278, 16),
37420 => conv_std_logic_vector(6424, 16),
37421 => conv_std_logic_vector(6570, 16),
37422 => conv_std_logic_vector(6716, 16),
37423 => conv_std_logic_vector(6862, 16),
37424 => conv_std_logic_vector(7008, 16),
37425 => conv_std_logic_vector(7154, 16),
37426 => conv_std_logic_vector(7300, 16),
37427 => conv_std_logic_vector(7446, 16),
37428 => conv_std_logic_vector(7592, 16),
37429 => conv_std_logic_vector(7738, 16),
37430 => conv_std_logic_vector(7884, 16),
37431 => conv_std_logic_vector(8030, 16),
37432 => conv_std_logic_vector(8176, 16),
37433 => conv_std_logic_vector(8322, 16),
37434 => conv_std_logic_vector(8468, 16),
37435 => conv_std_logic_vector(8614, 16),
37436 => conv_std_logic_vector(8760, 16),
37437 => conv_std_logic_vector(8906, 16),
37438 => conv_std_logic_vector(9052, 16),
37439 => conv_std_logic_vector(9198, 16),
37440 => conv_std_logic_vector(9344, 16),
37441 => conv_std_logic_vector(9490, 16),
37442 => conv_std_logic_vector(9636, 16),
37443 => conv_std_logic_vector(9782, 16),
37444 => conv_std_logic_vector(9928, 16),
37445 => conv_std_logic_vector(10074, 16),
37446 => conv_std_logic_vector(10220, 16),
37447 => conv_std_logic_vector(10366, 16),
37448 => conv_std_logic_vector(10512, 16),
37449 => conv_std_logic_vector(10658, 16),
37450 => conv_std_logic_vector(10804, 16),
37451 => conv_std_logic_vector(10950, 16),
37452 => conv_std_logic_vector(11096, 16),
37453 => conv_std_logic_vector(11242, 16),
37454 => conv_std_logic_vector(11388, 16),
37455 => conv_std_logic_vector(11534, 16),
37456 => conv_std_logic_vector(11680, 16),
37457 => conv_std_logic_vector(11826, 16),
37458 => conv_std_logic_vector(11972, 16),
37459 => conv_std_logic_vector(12118, 16),
37460 => conv_std_logic_vector(12264, 16),
37461 => conv_std_logic_vector(12410, 16),
37462 => conv_std_logic_vector(12556, 16),
37463 => conv_std_logic_vector(12702, 16),
37464 => conv_std_logic_vector(12848, 16),
37465 => conv_std_logic_vector(12994, 16),
37466 => conv_std_logic_vector(13140, 16),
37467 => conv_std_logic_vector(13286, 16),
37468 => conv_std_logic_vector(13432, 16),
37469 => conv_std_logic_vector(13578, 16),
37470 => conv_std_logic_vector(13724, 16),
37471 => conv_std_logic_vector(13870, 16),
37472 => conv_std_logic_vector(14016, 16),
37473 => conv_std_logic_vector(14162, 16),
37474 => conv_std_logic_vector(14308, 16),
37475 => conv_std_logic_vector(14454, 16),
37476 => conv_std_logic_vector(14600, 16),
37477 => conv_std_logic_vector(14746, 16),
37478 => conv_std_logic_vector(14892, 16),
37479 => conv_std_logic_vector(15038, 16),
37480 => conv_std_logic_vector(15184, 16),
37481 => conv_std_logic_vector(15330, 16),
37482 => conv_std_logic_vector(15476, 16),
37483 => conv_std_logic_vector(15622, 16),
37484 => conv_std_logic_vector(15768, 16),
37485 => conv_std_logic_vector(15914, 16),
37486 => conv_std_logic_vector(16060, 16),
37487 => conv_std_logic_vector(16206, 16),
37488 => conv_std_logic_vector(16352, 16),
37489 => conv_std_logic_vector(16498, 16),
37490 => conv_std_logic_vector(16644, 16),
37491 => conv_std_logic_vector(16790, 16),
37492 => conv_std_logic_vector(16936, 16),
37493 => conv_std_logic_vector(17082, 16),
37494 => conv_std_logic_vector(17228, 16),
37495 => conv_std_logic_vector(17374, 16),
37496 => conv_std_logic_vector(17520, 16),
37497 => conv_std_logic_vector(17666, 16),
37498 => conv_std_logic_vector(17812, 16),
37499 => conv_std_logic_vector(17958, 16),
37500 => conv_std_logic_vector(18104, 16),
37501 => conv_std_logic_vector(18250, 16),
37502 => conv_std_logic_vector(18396, 16),
37503 => conv_std_logic_vector(18542, 16),
37504 => conv_std_logic_vector(18688, 16),
37505 => conv_std_logic_vector(18834, 16),
37506 => conv_std_logic_vector(18980, 16),
37507 => conv_std_logic_vector(19126, 16),
37508 => conv_std_logic_vector(19272, 16),
37509 => conv_std_logic_vector(19418, 16),
37510 => conv_std_logic_vector(19564, 16),
37511 => conv_std_logic_vector(19710, 16),
37512 => conv_std_logic_vector(19856, 16),
37513 => conv_std_logic_vector(20002, 16),
37514 => conv_std_logic_vector(20148, 16),
37515 => conv_std_logic_vector(20294, 16),
37516 => conv_std_logic_vector(20440, 16),
37517 => conv_std_logic_vector(20586, 16),
37518 => conv_std_logic_vector(20732, 16),
37519 => conv_std_logic_vector(20878, 16),
37520 => conv_std_logic_vector(21024, 16),
37521 => conv_std_logic_vector(21170, 16),
37522 => conv_std_logic_vector(21316, 16),
37523 => conv_std_logic_vector(21462, 16),
37524 => conv_std_logic_vector(21608, 16),
37525 => conv_std_logic_vector(21754, 16),
37526 => conv_std_logic_vector(21900, 16),
37527 => conv_std_logic_vector(22046, 16),
37528 => conv_std_logic_vector(22192, 16),
37529 => conv_std_logic_vector(22338, 16),
37530 => conv_std_logic_vector(22484, 16),
37531 => conv_std_logic_vector(22630, 16),
37532 => conv_std_logic_vector(22776, 16),
37533 => conv_std_logic_vector(22922, 16),
37534 => conv_std_logic_vector(23068, 16),
37535 => conv_std_logic_vector(23214, 16),
37536 => conv_std_logic_vector(23360, 16),
37537 => conv_std_logic_vector(23506, 16),
37538 => conv_std_logic_vector(23652, 16),
37539 => conv_std_logic_vector(23798, 16),
37540 => conv_std_logic_vector(23944, 16),
37541 => conv_std_logic_vector(24090, 16),
37542 => conv_std_logic_vector(24236, 16),
37543 => conv_std_logic_vector(24382, 16),
37544 => conv_std_logic_vector(24528, 16),
37545 => conv_std_logic_vector(24674, 16),
37546 => conv_std_logic_vector(24820, 16),
37547 => conv_std_logic_vector(24966, 16),
37548 => conv_std_logic_vector(25112, 16),
37549 => conv_std_logic_vector(25258, 16),
37550 => conv_std_logic_vector(25404, 16),
37551 => conv_std_logic_vector(25550, 16),
37552 => conv_std_logic_vector(25696, 16),
37553 => conv_std_logic_vector(25842, 16),
37554 => conv_std_logic_vector(25988, 16),
37555 => conv_std_logic_vector(26134, 16),
37556 => conv_std_logic_vector(26280, 16),
37557 => conv_std_logic_vector(26426, 16),
37558 => conv_std_logic_vector(26572, 16),
37559 => conv_std_logic_vector(26718, 16),
37560 => conv_std_logic_vector(26864, 16),
37561 => conv_std_logic_vector(27010, 16),
37562 => conv_std_logic_vector(27156, 16),
37563 => conv_std_logic_vector(27302, 16),
37564 => conv_std_logic_vector(27448, 16),
37565 => conv_std_logic_vector(27594, 16),
37566 => conv_std_logic_vector(27740, 16),
37567 => conv_std_logic_vector(27886, 16),
37568 => conv_std_logic_vector(28032, 16),
37569 => conv_std_logic_vector(28178, 16),
37570 => conv_std_logic_vector(28324, 16),
37571 => conv_std_logic_vector(28470, 16),
37572 => conv_std_logic_vector(28616, 16),
37573 => conv_std_logic_vector(28762, 16),
37574 => conv_std_logic_vector(28908, 16),
37575 => conv_std_logic_vector(29054, 16),
37576 => conv_std_logic_vector(29200, 16),
37577 => conv_std_logic_vector(29346, 16),
37578 => conv_std_logic_vector(29492, 16),
37579 => conv_std_logic_vector(29638, 16),
37580 => conv_std_logic_vector(29784, 16),
37581 => conv_std_logic_vector(29930, 16),
37582 => conv_std_logic_vector(30076, 16),
37583 => conv_std_logic_vector(30222, 16),
37584 => conv_std_logic_vector(30368, 16),
37585 => conv_std_logic_vector(30514, 16),
37586 => conv_std_logic_vector(30660, 16),
37587 => conv_std_logic_vector(30806, 16),
37588 => conv_std_logic_vector(30952, 16),
37589 => conv_std_logic_vector(31098, 16),
37590 => conv_std_logic_vector(31244, 16),
37591 => conv_std_logic_vector(31390, 16),
37592 => conv_std_logic_vector(31536, 16),
37593 => conv_std_logic_vector(31682, 16),
37594 => conv_std_logic_vector(31828, 16),
37595 => conv_std_logic_vector(31974, 16),
37596 => conv_std_logic_vector(32120, 16),
37597 => conv_std_logic_vector(32266, 16),
37598 => conv_std_logic_vector(32412, 16),
37599 => conv_std_logic_vector(32558, 16),
37600 => conv_std_logic_vector(32704, 16),
37601 => conv_std_logic_vector(32850, 16),
37602 => conv_std_logic_vector(32996, 16),
37603 => conv_std_logic_vector(33142, 16),
37604 => conv_std_logic_vector(33288, 16),
37605 => conv_std_logic_vector(33434, 16),
37606 => conv_std_logic_vector(33580, 16),
37607 => conv_std_logic_vector(33726, 16),
37608 => conv_std_logic_vector(33872, 16),
37609 => conv_std_logic_vector(34018, 16),
37610 => conv_std_logic_vector(34164, 16),
37611 => conv_std_logic_vector(34310, 16),
37612 => conv_std_logic_vector(34456, 16),
37613 => conv_std_logic_vector(34602, 16),
37614 => conv_std_logic_vector(34748, 16),
37615 => conv_std_logic_vector(34894, 16),
37616 => conv_std_logic_vector(35040, 16),
37617 => conv_std_logic_vector(35186, 16),
37618 => conv_std_logic_vector(35332, 16),
37619 => conv_std_logic_vector(35478, 16),
37620 => conv_std_logic_vector(35624, 16),
37621 => conv_std_logic_vector(35770, 16),
37622 => conv_std_logic_vector(35916, 16),
37623 => conv_std_logic_vector(36062, 16),
37624 => conv_std_logic_vector(36208, 16),
37625 => conv_std_logic_vector(36354, 16),
37626 => conv_std_logic_vector(36500, 16),
37627 => conv_std_logic_vector(36646, 16),
37628 => conv_std_logic_vector(36792, 16),
37629 => conv_std_logic_vector(36938, 16),
37630 => conv_std_logic_vector(37084, 16),
37631 => conv_std_logic_vector(37230, 16),
37632 => conv_std_logic_vector(0, 16),
37633 => conv_std_logic_vector(147, 16),
37634 => conv_std_logic_vector(294, 16),
37635 => conv_std_logic_vector(441, 16),
37636 => conv_std_logic_vector(588, 16),
37637 => conv_std_logic_vector(735, 16),
37638 => conv_std_logic_vector(882, 16),
37639 => conv_std_logic_vector(1029, 16),
37640 => conv_std_logic_vector(1176, 16),
37641 => conv_std_logic_vector(1323, 16),
37642 => conv_std_logic_vector(1470, 16),
37643 => conv_std_logic_vector(1617, 16),
37644 => conv_std_logic_vector(1764, 16),
37645 => conv_std_logic_vector(1911, 16),
37646 => conv_std_logic_vector(2058, 16),
37647 => conv_std_logic_vector(2205, 16),
37648 => conv_std_logic_vector(2352, 16),
37649 => conv_std_logic_vector(2499, 16),
37650 => conv_std_logic_vector(2646, 16),
37651 => conv_std_logic_vector(2793, 16),
37652 => conv_std_logic_vector(2940, 16),
37653 => conv_std_logic_vector(3087, 16),
37654 => conv_std_logic_vector(3234, 16),
37655 => conv_std_logic_vector(3381, 16),
37656 => conv_std_logic_vector(3528, 16),
37657 => conv_std_logic_vector(3675, 16),
37658 => conv_std_logic_vector(3822, 16),
37659 => conv_std_logic_vector(3969, 16),
37660 => conv_std_logic_vector(4116, 16),
37661 => conv_std_logic_vector(4263, 16),
37662 => conv_std_logic_vector(4410, 16),
37663 => conv_std_logic_vector(4557, 16),
37664 => conv_std_logic_vector(4704, 16),
37665 => conv_std_logic_vector(4851, 16),
37666 => conv_std_logic_vector(4998, 16),
37667 => conv_std_logic_vector(5145, 16),
37668 => conv_std_logic_vector(5292, 16),
37669 => conv_std_logic_vector(5439, 16),
37670 => conv_std_logic_vector(5586, 16),
37671 => conv_std_logic_vector(5733, 16),
37672 => conv_std_logic_vector(5880, 16),
37673 => conv_std_logic_vector(6027, 16),
37674 => conv_std_logic_vector(6174, 16),
37675 => conv_std_logic_vector(6321, 16),
37676 => conv_std_logic_vector(6468, 16),
37677 => conv_std_logic_vector(6615, 16),
37678 => conv_std_logic_vector(6762, 16),
37679 => conv_std_logic_vector(6909, 16),
37680 => conv_std_logic_vector(7056, 16),
37681 => conv_std_logic_vector(7203, 16),
37682 => conv_std_logic_vector(7350, 16),
37683 => conv_std_logic_vector(7497, 16),
37684 => conv_std_logic_vector(7644, 16),
37685 => conv_std_logic_vector(7791, 16),
37686 => conv_std_logic_vector(7938, 16),
37687 => conv_std_logic_vector(8085, 16),
37688 => conv_std_logic_vector(8232, 16),
37689 => conv_std_logic_vector(8379, 16),
37690 => conv_std_logic_vector(8526, 16),
37691 => conv_std_logic_vector(8673, 16),
37692 => conv_std_logic_vector(8820, 16),
37693 => conv_std_logic_vector(8967, 16),
37694 => conv_std_logic_vector(9114, 16),
37695 => conv_std_logic_vector(9261, 16),
37696 => conv_std_logic_vector(9408, 16),
37697 => conv_std_logic_vector(9555, 16),
37698 => conv_std_logic_vector(9702, 16),
37699 => conv_std_logic_vector(9849, 16),
37700 => conv_std_logic_vector(9996, 16),
37701 => conv_std_logic_vector(10143, 16),
37702 => conv_std_logic_vector(10290, 16),
37703 => conv_std_logic_vector(10437, 16),
37704 => conv_std_logic_vector(10584, 16),
37705 => conv_std_logic_vector(10731, 16),
37706 => conv_std_logic_vector(10878, 16),
37707 => conv_std_logic_vector(11025, 16),
37708 => conv_std_logic_vector(11172, 16),
37709 => conv_std_logic_vector(11319, 16),
37710 => conv_std_logic_vector(11466, 16),
37711 => conv_std_logic_vector(11613, 16),
37712 => conv_std_logic_vector(11760, 16),
37713 => conv_std_logic_vector(11907, 16),
37714 => conv_std_logic_vector(12054, 16),
37715 => conv_std_logic_vector(12201, 16),
37716 => conv_std_logic_vector(12348, 16),
37717 => conv_std_logic_vector(12495, 16),
37718 => conv_std_logic_vector(12642, 16),
37719 => conv_std_logic_vector(12789, 16),
37720 => conv_std_logic_vector(12936, 16),
37721 => conv_std_logic_vector(13083, 16),
37722 => conv_std_logic_vector(13230, 16),
37723 => conv_std_logic_vector(13377, 16),
37724 => conv_std_logic_vector(13524, 16),
37725 => conv_std_logic_vector(13671, 16),
37726 => conv_std_logic_vector(13818, 16),
37727 => conv_std_logic_vector(13965, 16),
37728 => conv_std_logic_vector(14112, 16),
37729 => conv_std_logic_vector(14259, 16),
37730 => conv_std_logic_vector(14406, 16),
37731 => conv_std_logic_vector(14553, 16),
37732 => conv_std_logic_vector(14700, 16),
37733 => conv_std_logic_vector(14847, 16),
37734 => conv_std_logic_vector(14994, 16),
37735 => conv_std_logic_vector(15141, 16),
37736 => conv_std_logic_vector(15288, 16),
37737 => conv_std_logic_vector(15435, 16),
37738 => conv_std_logic_vector(15582, 16),
37739 => conv_std_logic_vector(15729, 16),
37740 => conv_std_logic_vector(15876, 16),
37741 => conv_std_logic_vector(16023, 16),
37742 => conv_std_logic_vector(16170, 16),
37743 => conv_std_logic_vector(16317, 16),
37744 => conv_std_logic_vector(16464, 16),
37745 => conv_std_logic_vector(16611, 16),
37746 => conv_std_logic_vector(16758, 16),
37747 => conv_std_logic_vector(16905, 16),
37748 => conv_std_logic_vector(17052, 16),
37749 => conv_std_logic_vector(17199, 16),
37750 => conv_std_logic_vector(17346, 16),
37751 => conv_std_logic_vector(17493, 16),
37752 => conv_std_logic_vector(17640, 16),
37753 => conv_std_logic_vector(17787, 16),
37754 => conv_std_logic_vector(17934, 16),
37755 => conv_std_logic_vector(18081, 16),
37756 => conv_std_logic_vector(18228, 16),
37757 => conv_std_logic_vector(18375, 16),
37758 => conv_std_logic_vector(18522, 16),
37759 => conv_std_logic_vector(18669, 16),
37760 => conv_std_logic_vector(18816, 16),
37761 => conv_std_logic_vector(18963, 16),
37762 => conv_std_logic_vector(19110, 16),
37763 => conv_std_logic_vector(19257, 16),
37764 => conv_std_logic_vector(19404, 16),
37765 => conv_std_logic_vector(19551, 16),
37766 => conv_std_logic_vector(19698, 16),
37767 => conv_std_logic_vector(19845, 16),
37768 => conv_std_logic_vector(19992, 16),
37769 => conv_std_logic_vector(20139, 16),
37770 => conv_std_logic_vector(20286, 16),
37771 => conv_std_logic_vector(20433, 16),
37772 => conv_std_logic_vector(20580, 16),
37773 => conv_std_logic_vector(20727, 16),
37774 => conv_std_logic_vector(20874, 16),
37775 => conv_std_logic_vector(21021, 16),
37776 => conv_std_logic_vector(21168, 16),
37777 => conv_std_logic_vector(21315, 16),
37778 => conv_std_logic_vector(21462, 16),
37779 => conv_std_logic_vector(21609, 16),
37780 => conv_std_logic_vector(21756, 16),
37781 => conv_std_logic_vector(21903, 16),
37782 => conv_std_logic_vector(22050, 16),
37783 => conv_std_logic_vector(22197, 16),
37784 => conv_std_logic_vector(22344, 16),
37785 => conv_std_logic_vector(22491, 16),
37786 => conv_std_logic_vector(22638, 16),
37787 => conv_std_logic_vector(22785, 16),
37788 => conv_std_logic_vector(22932, 16),
37789 => conv_std_logic_vector(23079, 16),
37790 => conv_std_logic_vector(23226, 16),
37791 => conv_std_logic_vector(23373, 16),
37792 => conv_std_logic_vector(23520, 16),
37793 => conv_std_logic_vector(23667, 16),
37794 => conv_std_logic_vector(23814, 16),
37795 => conv_std_logic_vector(23961, 16),
37796 => conv_std_logic_vector(24108, 16),
37797 => conv_std_logic_vector(24255, 16),
37798 => conv_std_logic_vector(24402, 16),
37799 => conv_std_logic_vector(24549, 16),
37800 => conv_std_logic_vector(24696, 16),
37801 => conv_std_logic_vector(24843, 16),
37802 => conv_std_logic_vector(24990, 16),
37803 => conv_std_logic_vector(25137, 16),
37804 => conv_std_logic_vector(25284, 16),
37805 => conv_std_logic_vector(25431, 16),
37806 => conv_std_logic_vector(25578, 16),
37807 => conv_std_logic_vector(25725, 16),
37808 => conv_std_logic_vector(25872, 16),
37809 => conv_std_logic_vector(26019, 16),
37810 => conv_std_logic_vector(26166, 16),
37811 => conv_std_logic_vector(26313, 16),
37812 => conv_std_logic_vector(26460, 16),
37813 => conv_std_logic_vector(26607, 16),
37814 => conv_std_logic_vector(26754, 16),
37815 => conv_std_logic_vector(26901, 16),
37816 => conv_std_logic_vector(27048, 16),
37817 => conv_std_logic_vector(27195, 16),
37818 => conv_std_logic_vector(27342, 16),
37819 => conv_std_logic_vector(27489, 16),
37820 => conv_std_logic_vector(27636, 16),
37821 => conv_std_logic_vector(27783, 16),
37822 => conv_std_logic_vector(27930, 16),
37823 => conv_std_logic_vector(28077, 16),
37824 => conv_std_logic_vector(28224, 16),
37825 => conv_std_logic_vector(28371, 16),
37826 => conv_std_logic_vector(28518, 16),
37827 => conv_std_logic_vector(28665, 16),
37828 => conv_std_logic_vector(28812, 16),
37829 => conv_std_logic_vector(28959, 16),
37830 => conv_std_logic_vector(29106, 16),
37831 => conv_std_logic_vector(29253, 16),
37832 => conv_std_logic_vector(29400, 16),
37833 => conv_std_logic_vector(29547, 16),
37834 => conv_std_logic_vector(29694, 16),
37835 => conv_std_logic_vector(29841, 16),
37836 => conv_std_logic_vector(29988, 16),
37837 => conv_std_logic_vector(30135, 16),
37838 => conv_std_logic_vector(30282, 16),
37839 => conv_std_logic_vector(30429, 16),
37840 => conv_std_logic_vector(30576, 16),
37841 => conv_std_logic_vector(30723, 16),
37842 => conv_std_logic_vector(30870, 16),
37843 => conv_std_logic_vector(31017, 16),
37844 => conv_std_logic_vector(31164, 16),
37845 => conv_std_logic_vector(31311, 16),
37846 => conv_std_logic_vector(31458, 16),
37847 => conv_std_logic_vector(31605, 16),
37848 => conv_std_logic_vector(31752, 16),
37849 => conv_std_logic_vector(31899, 16),
37850 => conv_std_logic_vector(32046, 16),
37851 => conv_std_logic_vector(32193, 16),
37852 => conv_std_logic_vector(32340, 16),
37853 => conv_std_logic_vector(32487, 16),
37854 => conv_std_logic_vector(32634, 16),
37855 => conv_std_logic_vector(32781, 16),
37856 => conv_std_logic_vector(32928, 16),
37857 => conv_std_logic_vector(33075, 16),
37858 => conv_std_logic_vector(33222, 16),
37859 => conv_std_logic_vector(33369, 16),
37860 => conv_std_logic_vector(33516, 16),
37861 => conv_std_logic_vector(33663, 16),
37862 => conv_std_logic_vector(33810, 16),
37863 => conv_std_logic_vector(33957, 16),
37864 => conv_std_logic_vector(34104, 16),
37865 => conv_std_logic_vector(34251, 16),
37866 => conv_std_logic_vector(34398, 16),
37867 => conv_std_logic_vector(34545, 16),
37868 => conv_std_logic_vector(34692, 16),
37869 => conv_std_logic_vector(34839, 16),
37870 => conv_std_logic_vector(34986, 16),
37871 => conv_std_logic_vector(35133, 16),
37872 => conv_std_logic_vector(35280, 16),
37873 => conv_std_logic_vector(35427, 16),
37874 => conv_std_logic_vector(35574, 16),
37875 => conv_std_logic_vector(35721, 16),
37876 => conv_std_logic_vector(35868, 16),
37877 => conv_std_logic_vector(36015, 16),
37878 => conv_std_logic_vector(36162, 16),
37879 => conv_std_logic_vector(36309, 16),
37880 => conv_std_logic_vector(36456, 16),
37881 => conv_std_logic_vector(36603, 16),
37882 => conv_std_logic_vector(36750, 16),
37883 => conv_std_logic_vector(36897, 16),
37884 => conv_std_logic_vector(37044, 16),
37885 => conv_std_logic_vector(37191, 16),
37886 => conv_std_logic_vector(37338, 16),
37887 => conv_std_logic_vector(37485, 16),
37888 => conv_std_logic_vector(0, 16),
37889 => conv_std_logic_vector(148, 16),
37890 => conv_std_logic_vector(296, 16),
37891 => conv_std_logic_vector(444, 16),
37892 => conv_std_logic_vector(592, 16),
37893 => conv_std_logic_vector(740, 16),
37894 => conv_std_logic_vector(888, 16),
37895 => conv_std_logic_vector(1036, 16),
37896 => conv_std_logic_vector(1184, 16),
37897 => conv_std_logic_vector(1332, 16),
37898 => conv_std_logic_vector(1480, 16),
37899 => conv_std_logic_vector(1628, 16),
37900 => conv_std_logic_vector(1776, 16),
37901 => conv_std_logic_vector(1924, 16),
37902 => conv_std_logic_vector(2072, 16),
37903 => conv_std_logic_vector(2220, 16),
37904 => conv_std_logic_vector(2368, 16),
37905 => conv_std_logic_vector(2516, 16),
37906 => conv_std_logic_vector(2664, 16),
37907 => conv_std_logic_vector(2812, 16),
37908 => conv_std_logic_vector(2960, 16),
37909 => conv_std_logic_vector(3108, 16),
37910 => conv_std_logic_vector(3256, 16),
37911 => conv_std_logic_vector(3404, 16),
37912 => conv_std_logic_vector(3552, 16),
37913 => conv_std_logic_vector(3700, 16),
37914 => conv_std_logic_vector(3848, 16),
37915 => conv_std_logic_vector(3996, 16),
37916 => conv_std_logic_vector(4144, 16),
37917 => conv_std_logic_vector(4292, 16),
37918 => conv_std_logic_vector(4440, 16),
37919 => conv_std_logic_vector(4588, 16),
37920 => conv_std_logic_vector(4736, 16),
37921 => conv_std_logic_vector(4884, 16),
37922 => conv_std_logic_vector(5032, 16),
37923 => conv_std_logic_vector(5180, 16),
37924 => conv_std_logic_vector(5328, 16),
37925 => conv_std_logic_vector(5476, 16),
37926 => conv_std_logic_vector(5624, 16),
37927 => conv_std_logic_vector(5772, 16),
37928 => conv_std_logic_vector(5920, 16),
37929 => conv_std_logic_vector(6068, 16),
37930 => conv_std_logic_vector(6216, 16),
37931 => conv_std_logic_vector(6364, 16),
37932 => conv_std_logic_vector(6512, 16),
37933 => conv_std_logic_vector(6660, 16),
37934 => conv_std_logic_vector(6808, 16),
37935 => conv_std_logic_vector(6956, 16),
37936 => conv_std_logic_vector(7104, 16),
37937 => conv_std_logic_vector(7252, 16),
37938 => conv_std_logic_vector(7400, 16),
37939 => conv_std_logic_vector(7548, 16),
37940 => conv_std_logic_vector(7696, 16),
37941 => conv_std_logic_vector(7844, 16),
37942 => conv_std_logic_vector(7992, 16),
37943 => conv_std_logic_vector(8140, 16),
37944 => conv_std_logic_vector(8288, 16),
37945 => conv_std_logic_vector(8436, 16),
37946 => conv_std_logic_vector(8584, 16),
37947 => conv_std_logic_vector(8732, 16),
37948 => conv_std_logic_vector(8880, 16),
37949 => conv_std_logic_vector(9028, 16),
37950 => conv_std_logic_vector(9176, 16),
37951 => conv_std_logic_vector(9324, 16),
37952 => conv_std_logic_vector(9472, 16),
37953 => conv_std_logic_vector(9620, 16),
37954 => conv_std_logic_vector(9768, 16),
37955 => conv_std_logic_vector(9916, 16),
37956 => conv_std_logic_vector(10064, 16),
37957 => conv_std_logic_vector(10212, 16),
37958 => conv_std_logic_vector(10360, 16),
37959 => conv_std_logic_vector(10508, 16),
37960 => conv_std_logic_vector(10656, 16),
37961 => conv_std_logic_vector(10804, 16),
37962 => conv_std_logic_vector(10952, 16),
37963 => conv_std_logic_vector(11100, 16),
37964 => conv_std_logic_vector(11248, 16),
37965 => conv_std_logic_vector(11396, 16),
37966 => conv_std_logic_vector(11544, 16),
37967 => conv_std_logic_vector(11692, 16),
37968 => conv_std_logic_vector(11840, 16),
37969 => conv_std_logic_vector(11988, 16),
37970 => conv_std_logic_vector(12136, 16),
37971 => conv_std_logic_vector(12284, 16),
37972 => conv_std_logic_vector(12432, 16),
37973 => conv_std_logic_vector(12580, 16),
37974 => conv_std_logic_vector(12728, 16),
37975 => conv_std_logic_vector(12876, 16),
37976 => conv_std_logic_vector(13024, 16),
37977 => conv_std_logic_vector(13172, 16),
37978 => conv_std_logic_vector(13320, 16),
37979 => conv_std_logic_vector(13468, 16),
37980 => conv_std_logic_vector(13616, 16),
37981 => conv_std_logic_vector(13764, 16),
37982 => conv_std_logic_vector(13912, 16),
37983 => conv_std_logic_vector(14060, 16),
37984 => conv_std_logic_vector(14208, 16),
37985 => conv_std_logic_vector(14356, 16),
37986 => conv_std_logic_vector(14504, 16),
37987 => conv_std_logic_vector(14652, 16),
37988 => conv_std_logic_vector(14800, 16),
37989 => conv_std_logic_vector(14948, 16),
37990 => conv_std_logic_vector(15096, 16),
37991 => conv_std_logic_vector(15244, 16),
37992 => conv_std_logic_vector(15392, 16),
37993 => conv_std_logic_vector(15540, 16),
37994 => conv_std_logic_vector(15688, 16),
37995 => conv_std_logic_vector(15836, 16),
37996 => conv_std_logic_vector(15984, 16),
37997 => conv_std_logic_vector(16132, 16),
37998 => conv_std_logic_vector(16280, 16),
37999 => conv_std_logic_vector(16428, 16),
38000 => conv_std_logic_vector(16576, 16),
38001 => conv_std_logic_vector(16724, 16),
38002 => conv_std_logic_vector(16872, 16),
38003 => conv_std_logic_vector(17020, 16),
38004 => conv_std_logic_vector(17168, 16),
38005 => conv_std_logic_vector(17316, 16),
38006 => conv_std_logic_vector(17464, 16),
38007 => conv_std_logic_vector(17612, 16),
38008 => conv_std_logic_vector(17760, 16),
38009 => conv_std_logic_vector(17908, 16),
38010 => conv_std_logic_vector(18056, 16),
38011 => conv_std_logic_vector(18204, 16),
38012 => conv_std_logic_vector(18352, 16),
38013 => conv_std_logic_vector(18500, 16),
38014 => conv_std_logic_vector(18648, 16),
38015 => conv_std_logic_vector(18796, 16),
38016 => conv_std_logic_vector(18944, 16),
38017 => conv_std_logic_vector(19092, 16),
38018 => conv_std_logic_vector(19240, 16),
38019 => conv_std_logic_vector(19388, 16),
38020 => conv_std_logic_vector(19536, 16),
38021 => conv_std_logic_vector(19684, 16),
38022 => conv_std_logic_vector(19832, 16),
38023 => conv_std_logic_vector(19980, 16),
38024 => conv_std_logic_vector(20128, 16),
38025 => conv_std_logic_vector(20276, 16),
38026 => conv_std_logic_vector(20424, 16),
38027 => conv_std_logic_vector(20572, 16),
38028 => conv_std_logic_vector(20720, 16),
38029 => conv_std_logic_vector(20868, 16),
38030 => conv_std_logic_vector(21016, 16),
38031 => conv_std_logic_vector(21164, 16),
38032 => conv_std_logic_vector(21312, 16),
38033 => conv_std_logic_vector(21460, 16),
38034 => conv_std_logic_vector(21608, 16),
38035 => conv_std_logic_vector(21756, 16),
38036 => conv_std_logic_vector(21904, 16),
38037 => conv_std_logic_vector(22052, 16),
38038 => conv_std_logic_vector(22200, 16),
38039 => conv_std_logic_vector(22348, 16),
38040 => conv_std_logic_vector(22496, 16),
38041 => conv_std_logic_vector(22644, 16),
38042 => conv_std_logic_vector(22792, 16),
38043 => conv_std_logic_vector(22940, 16),
38044 => conv_std_logic_vector(23088, 16),
38045 => conv_std_logic_vector(23236, 16),
38046 => conv_std_logic_vector(23384, 16),
38047 => conv_std_logic_vector(23532, 16),
38048 => conv_std_logic_vector(23680, 16),
38049 => conv_std_logic_vector(23828, 16),
38050 => conv_std_logic_vector(23976, 16),
38051 => conv_std_logic_vector(24124, 16),
38052 => conv_std_logic_vector(24272, 16),
38053 => conv_std_logic_vector(24420, 16),
38054 => conv_std_logic_vector(24568, 16),
38055 => conv_std_logic_vector(24716, 16),
38056 => conv_std_logic_vector(24864, 16),
38057 => conv_std_logic_vector(25012, 16),
38058 => conv_std_logic_vector(25160, 16),
38059 => conv_std_logic_vector(25308, 16),
38060 => conv_std_logic_vector(25456, 16),
38061 => conv_std_logic_vector(25604, 16),
38062 => conv_std_logic_vector(25752, 16),
38063 => conv_std_logic_vector(25900, 16),
38064 => conv_std_logic_vector(26048, 16),
38065 => conv_std_logic_vector(26196, 16),
38066 => conv_std_logic_vector(26344, 16),
38067 => conv_std_logic_vector(26492, 16),
38068 => conv_std_logic_vector(26640, 16),
38069 => conv_std_logic_vector(26788, 16),
38070 => conv_std_logic_vector(26936, 16),
38071 => conv_std_logic_vector(27084, 16),
38072 => conv_std_logic_vector(27232, 16),
38073 => conv_std_logic_vector(27380, 16),
38074 => conv_std_logic_vector(27528, 16),
38075 => conv_std_logic_vector(27676, 16),
38076 => conv_std_logic_vector(27824, 16),
38077 => conv_std_logic_vector(27972, 16),
38078 => conv_std_logic_vector(28120, 16),
38079 => conv_std_logic_vector(28268, 16),
38080 => conv_std_logic_vector(28416, 16),
38081 => conv_std_logic_vector(28564, 16),
38082 => conv_std_logic_vector(28712, 16),
38083 => conv_std_logic_vector(28860, 16),
38084 => conv_std_logic_vector(29008, 16),
38085 => conv_std_logic_vector(29156, 16),
38086 => conv_std_logic_vector(29304, 16),
38087 => conv_std_logic_vector(29452, 16),
38088 => conv_std_logic_vector(29600, 16),
38089 => conv_std_logic_vector(29748, 16),
38090 => conv_std_logic_vector(29896, 16),
38091 => conv_std_logic_vector(30044, 16),
38092 => conv_std_logic_vector(30192, 16),
38093 => conv_std_logic_vector(30340, 16),
38094 => conv_std_logic_vector(30488, 16),
38095 => conv_std_logic_vector(30636, 16),
38096 => conv_std_logic_vector(30784, 16),
38097 => conv_std_logic_vector(30932, 16),
38098 => conv_std_logic_vector(31080, 16),
38099 => conv_std_logic_vector(31228, 16),
38100 => conv_std_logic_vector(31376, 16),
38101 => conv_std_logic_vector(31524, 16),
38102 => conv_std_logic_vector(31672, 16),
38103 => conv_std_logic_vector(31820, 16),
38104 => conv_std_logic_vector(31968, 16),
38105 => conv_std_logic_vector(32116, 16),
38106 => conv_std_logic_vector(32264, 16),
38107 => conv_std_logic_vector(32412, 16),
38108 => conv_std_logic_vector(32560, 16),
38109 => conv_std_logic_vector(32708, 16),
38110 => conv_std_logic_vector(32856, 16),
38111 => conv_std_logic_vector(33004, 16),
38112 => conv_std_logic_vector(33152, 16),
38113 => conv_std_logic_vector(33300, 16),
38114 => conv_std_logic_vector(33448, 16),
38115 => conv_std_logic_vector(33596, 16),
38116 => conv_std_logic_vector(33744, 16),
38117 => conv_std_logic_vector(33892, 16),
38118 => conv_std_logic_vector(34040, 16),
38119 => conv_std_logic_vector(34188, 16),
38120 => conv_std_logic_vector(34336, 16),
38121 => conv_std_logic_vector(34484, 16),
38122 => conv_std_logic_vector(34632, 16),
38123 => conv_std_logic_vector(34780, 16),
38124 => conv_std_logic_vector(34928, 16),
38125 => conv_std_logic_vector(35076, 16),
38126 => conv_std_logic_vector(35224, 16),
38127 => conv_std_logic_vector(35372, 16),
38128 => conv_std_logic_vector(35520, 16),
38129 => conv_std_logic_vector(35668, 16),
38130 => conv_std_logic_vector(35816, 16),
38131 => conv_std_logic_vector(35964, 16),
38132 => conv_std_logic_vector(36112, 16),
38133 => conv_std_logic_vector(36260, 16),
38134 => conv_std_logic_vector(36408, 16),
38135 => conv_std_logic_vector(36556, 16),
38136 => conv_std_logic_vector(36704, 16),
38137 => conv_std_logic_vector(36852, 16),
38138 => conv_std_logic_vector(37000, 16),
38139 => conv_std_logic_vector(37148, 16),
38140 => conv_std_logic_vector(37296, 16),
38141 => conv_std_logic_vector(37444, 16),
38142 => conv_std_logic_vector(37592, 16),
38143 => conv_std_logic_vector(37740, 16),
38144 => conv_std_logic_vector(0, 16),
38145 => conv_std_logic_vector(149, 16),
38146 => conv_std_logic_vector(298, 16),
38147 => conv_std_logic_vector(447, 16),
38148 => conv_std_logic_vector(596, 16),
38149 => conv_std_logic_vector(745, 16),
38150 => conv_std_logic_vector(894, 16),
38151 => conv_std_logic_vector(1043, 16),
38152 => conv_std_logic_vector(1192, 16),
38153 => conv_std_logic_vector(1341, 16),
38154 => conv_std_logic_vector(1490, 16),
38155 => conv_std_logic_vector(1639, 16),
38156 => conv_std_logic_vector(1788, 16),
38157 => conv_std_logic_vector(1937, 16),
38158 => conv_std_logic_vector(2086, 16),
38159 => conv_std_logic_vector(2235, 16),
38160 => conv_std_logic_vector(2384, 16),
38161 => conv_std_logic_vector(2533, 16),
38162 => conv_std_logic_vector(2682, 16),
38163 => conv_std_logic_vector(2831, 16),
38164 => conv_std_logic_vector(2980, 16),
38165 => conv_std_logic_vector(3129, 16),
38166 => conv_std_logic_vector(3278, 16),
38167 => conv_std_logic_vector(3427, 16),
38168 => conv_std_logic_vector(3576, 16),
38169 => conv_std_logic_vector(3725, 16),
38170 => conv_std_logic_vector(3874, 16),
38171 => conv_std_logic_vector(4023, 16),
38172 => conv_std_logic_vector(4172, 16),
38173 => conv_std_logic_vector(4321, 16),
38174 => conv_std_logic_vector(4470, 16),
38175 => conv_std_logic_vector(4619, 16),
38176 => conv_std_logic_vector(4768, 16),
38177 => conv_std_logic_vector(4917, 16),
38178 => conv_std_logic_vector(5066, 16),
38179 => conv_std_logic_vector(5215, 16),
38180 => conv_std_logic_vector(5364, 16),
38181 => conv_std_logic_vector(5513, 16),
38182 => conv_std_logic_vector(5662, 16),
38183 => conv_std_logic_vector(5811, 16),
38184 => conv_std_logic_vector(5960, 16),
38185 => conv_std_logic_vector(6109, 16),
38186 => conv_std_logic_vector(6258, 16),
38187 => conv_std_logic_vector(6407, 16),
38188 => conv_std_logic_vector(6556, 16),
38189 => conv_std_logic_vector(6705, 16),
38190 => conv_std_logic_vector(6854, 16),
38191 => conv_std_logic_vector(7003, 16),
38192 => conv_std_logic_vector(7152, 16),
38193 => conv_std_logic_vector(7301, 16),
38194 => conv_std_logic_vector(7450, 16),
38195 => conv_std_logic_vector(7599, 16),
38196 => conv_std_logic_vector(7748, 16),
38197 => conv_std_logic_vector(7897, 16),
38198 => conv_std_logic_vector(8046, 16),
38199 => conv_std_logic_vector(8195, 16),
38200 => conv_std_logic_vector(8344, 16),
38201 => conv_std_logic_vector(8493, 16),
38202 => conv_std_logic_vector(8642, 16),
38203 => conv_std_logic_vector(8791, 16),
38204 => conv_std_logic_vector(8940, 16),
38205 => conv_std_logic_vector(9089, 16),
38206 => conv_std_logic_vector(9238, 16),
38207 => conv_std_logic_vector(9387, 16),
38208 => conv_std_logic_vector(9536, 16),
38209 => conv_std_logic_vector(9685, 16),
38210 => conv_std_logic_vector(9834, 16),
38211 => conv_std_logic_vector(9983, 16),
38212 => conv_std_logic_vector(10132, 16),
38213 => conv_std_logic_vector(10281, 16),
38214 => conv_std_logic_vector(10430, 16),
38215 => conv_std_logic_vector(10579, 16),
38216 => conv_std_logic_vector(10728, 16),
38217 => conv_std_logic_vector(10877, 16),
38218 => conv_std_logic_vector(11026, 16),
38219 => conv_std_logic_vector(11175, 16),
38220 => conv_std_logic_vector(11324, 16),
38221 => conv_std_logic_vector(11473, 16),
38222 => conv_std_logic_vector(11622, 16),
38223 => conv_std_logic_vector(11771, 16),
38224 => conv_std_logic_vector(11920, 16),
38225 => conv_std_logic_vector(12069, 16),
38226 => conv_std_logic_vector(12218, 16),
38227 => conv_std_logic_vector(12367, 16),
38228 => conv_std_logic_vector(12516, 16),
38229 => conv_std_logic_vector(12665, 16),
38230 => conv_std_logic_vector(12814, 16),
38231 => conv_std_logic_vector(12963, 16),
38232 => conv_std_logic_vector(13112, 16),
38233 => conv_std_logic_vector(13261, 16),
38234 => conv_std_logic_vector(13410, 16),
38235 => conv_std_logic_vector(13559, 16),
38236 => conv_std_logic_vector(13708, 16),
38237 => conv_std_logic_vector(13857, 16),
38238 => conv_std_logic_vector(14006, 16),
38239 => conv_std_logic_vector(14155, 16),
38240 => conv_std_logic_vector(14304, 16),
38241 => conv_std_logic_vector(14453, 16),
38242 => conv_std_logic_vector(14602, 16),
38243 => conv_std_logic_vector(14751, 16),
38244 => conv_std_logic_vector(14900, 16),
38245 => conv_std_logic_vector(15049, 16),
38246 => conv_std_logic_vector(15198, 16),
38247 => conv_std_logic_vector(15347, 16),
38248 => conv_std_logic_vector(15496, 16),
38249 => conv_std_logic_vector(15645, 16),
38250 => conv_std_logic_vector(15794, 16),
38251 => conv_std_logic_vector(15943, 16),
38252 => conv_std_logic_vector(16092, 16),
38253 => conv_std_logic_vector(16241, 16),
38254 => conv_std_logic_vector(16390, 16),
38255 => conv_std_logic_vector(16539, 16),
38256 => conv_std_logic_vector(16688, 16),
38257 => conv_std_logic_vector(16837, 16),
38258 => conv_std_logic_vector(16986, 16),
38259 => conv_std_logic_vector(17135, 16),
38260 => conv_std_logic_vector(17284, 16),
38261 => conv_std_logic_vector(17433, 16),
38262 => conv_std_logic_vector(17582, 16),
38263 => conv_std_logic_vector(17731, 16),
38264 => conv_std_logic_vector(17880, 16),
38265 => conv_std_logic_vector(18029, 16),
38266 => conv_std_logic_vector(18178, 16),
38267 => conv_std_logic_vector(18327, 16),
38268 => conv_std_logic_vector(18476, 16),
38269 => conv_std_logic_vector(18625, 16),
38270 => conv_std_logic_vector(18774, 16),
38271 => conv_std_logic_vector(18923, 16),
38272 => conv_std_logic_vector(19072, 16),
38273 => conv_std_logic_vector(19221, 16),
38274 => conv_std_logic_vector(19370, 16),
38275 => conv_std_logic_vector(19519, 16),
38276 => conv_std_logic_vector(19668, 16),
38277 => conv_std_logic_vector(19817, 16),
38278 => conv_std_logic_vector(19966, 16),
38279 => conv_std_logic_vector(20115, 16),
38280 => conv_std_logic_vector(20264, 16),
38281 => conv_std_logic_vector(20413, 16),
38282 => conv_std_logic_vector(20562, 16),
38283 => conv_std_logic_vector(20711, 16),
38284 => conv_std_logic_vector(20860, 16),
38285 => conv_std_logic_vector(21009, 16),
38286 => conv_std_logic_vector(21158, 16),
38287 => conv_std_logic_vector(21307, 16),
38288 => conv_std_logic_vector(21456, 16),
38289 => conv_std_logic_vector(21605, 16),
38290 => conv_std_logic_vector(21754, 16),
38291 => conv_std_logic_vector(21903, 16),
38292 => conv_std_logic_vector(22052, 16),
38293 => conv_std_logic_vector(22201, 16),
38294 => conv_std_logic_vector(22350, 16),
38295 => conv_std_logic_vector(22499, 16),
38296 => conv_std_logic_vector(22648, 16),
38297 => conv_std_logic_vector(22797, 16),
38298 => conv_std_logic_vector(22946, 16),
38299 => conv_std_logic_vector(23095, 16),
38300 => conv_std_logic_vector(23244, 16),
38301 => conv_std_logic_vector(23393, 16),
38302 => conv_std_logic_vector(23542, 16),
38303 => conv_std_logic_vector(23691, 16),
38304 => conv_std_logic_vector(23840, 16),
38305 => conv_std_logic_vector(23989, 16),
38306 => conv_std_logic_vector(24138, 16),
38307 => conv_std_logic_vector(24287, 16),
38308 => conv_std_logic_vector(24436, 16),
38309 => conv_std_logic_vector(24585, 16),
38310 => conv_std_logic_vector(24734, 16),
38311 => conv_std_logic_vector(24883, 16),
38312 => conv_std_logic_vector(25032, 16),
38313 => conv_std_logic_vector(25181, 16),
38314 => conv_std_logic_vector(25330, 16),
38315 => conv_std_logic_vector(25479, 16),
38316 => conv_std_logic_vector(25628, 16),
38317 => conv_std_logic_vector(25777, 16),
38318 => conv_std_logic_vector(25926, 16),
38319 => conv_std_logic_vector(26075, 16),
38320 => conv_std_logic_vector(26224, 16),
38321 => conv_std_logic_vector(26373, 16),
38322 => conv_std_logic_vector(26522, 16),
38323 => conv_std_logic_vector(26671, 16),
38324 => conv_std_logic_vector(26820, 16),
38325 => conv_std_logic_vector(26969, 16),
38326 => conv_std_logic_vector(27118, 16),
38327 => conv_std_logic_vector(27267, 16),
38328 => conv_std_logic_vector(27416, 16),
38329 => conv_std_logic_vector(27565, 16),
38330 => conv_std_logic_vector(27714, 16),
38331 => conv_std_logic_vector(27863, 16),
38332 => conv_std_logic_vector(28012, 16),
38333 => conv_std_logic_vector(28161, 16),
38334 => conv_std_logic_vector(28310, 16),
38335 => conv_std_logic_vector(28459, 16),
38336 => conv_std_logic_vector(28608, 16),
38337 => conv_std_logic_vector(28757, 16),
38338 => conv_std_logic_vector(28906, 16),
38339 => conv_std_logic_vector(29055, 16),
38340 => conv_std_logic_vector(29204, 16),
38341 => conv_std_logic_vector(29353, 16),
38342 => conv_std_logic_vector(29502, 16),
38343 => conv_std_logic_vector(29651, 16),
38344 => conv_std_logic_vector(29800, 16),
38345 => conv_std_logic_vector(29949, 16),
38346 => conv_std_logic_vector(30098, 16),
38347 => conv_std_logic_vector(30247, 16),
38348 => conv_std_logic_vector(30396, 16),
38349 => conv_std_logic_vector(30545, 16),
38350 => conv_std_logic_vector(30694, 16),
38351 => conv_std_logic_vector(30843, 16),
38352 => conv_std_logic_vector(30992, 16),
38353 => conv_std_logic_vector(31141, 16),
38354 => conv_std_logic_vector(31290, 16),
38355 => conv_std_logic_vector(31439, 16),
38356 => conv_std_logic_vector(31588, 16),
38357 => conv_std_logic_vector(31737, 16),
38358 => conv_std_logic_vector(31886, 16),
38359 => conv_std_logic_vector(32035, 16),
38360 => conv_std_logic_vector(32184, 16),
38361 => conv_std_logic_vector(32333, 16),
38362 => conv_std_logic_vector(32482, 16),
38363 => conv_std_logic_vector(32631, 16),
38364 => conv_std_logic_vector(32780, 16),
38365 => conv_std_logic_vector(32929, 16),
38366 => conv_std_logic_vector(33078, 16),
38367 => conv_std_logic_vector(33227, 16),
38368 => conv_std_logic_vector(33376, 16),
38369 => conv_std_logic_vector(33525, 16),
38370 => conv_std_logic_vector(33674, 16),
38371 => conv_std_logic_vector(33823, 16),
38372 => conv_std_logic_vector(33972, 16),
38373 => conv_std_logic_vector(34121, 16),
38374 => conv_std_logic_vector(34270, 16),
38375 => conv_std_logic_vector(34419, 16),
38376 => conv_std_logic_vector(34568, 16),
38377 => conv_std_logic_vector(34717, 16),
38378 => conv_std_logic_vector(34866, 16),
38379 => conv_std_logic_vector(35015, 16),
38380 => conv_std_logic_vector(35164, 16),
38381 => conv_std_logic_vector(35313, 16),
38382 => conv_std_logic_vector(35462, 16),
38383 => conv_std_logic_vector(35611, 16),
38384 => conv_std_logic_vector(35760, 16),
38385 => conv_std_logic_vector(35909, 16),
38386 => conv_std_logic_vector(36058, 16),
38387 => conv_std_logic_vector(36207, 16),
38388 => conv_std_logic_vector(36356, 16),
38389 => conv_std_logic_vector(36505, 16),
38390 => conv_std_logic_vector(36654, 16),
38391 => conv_std_logic_vector(36803, 16),
38392 => conv_std_logic_vector(36952, 16),
38393 => conv_std_logic_vector(37101, 16),
38394 => conv_std_logic_vector(37250, 16),
38395 => conv_std_logic_vector(37399, 16),
38396 => conv_std_logic_vector(37548, 16),
38397 => conv_std_logic_vector(37697, 16),
38398 => conv_std_logic_vector(37846, 16),
38399 => conv_std_logic_vector(37995, 16),
38400 => conv_std_logic_vector(0, 16),
38401 => conv_std_logic_vector(150, 16),
38402 => conv_std_logic_vector(300, 16),
38403 => conv_std_logic_vector(450, 16),
38404 => conv_std_logic_vector(600, 16),
38405 => conv_std_logic_vector(750, 16),
38406 => conv_std_logic_vector(900, 16),
38407 => conv_std_logic_vector(1050, 16),
38408 => conv_std_logic_vector(1200, 16),
38409 => conv_std_logic_vector(1350, 16),
38410 => conv_std_logic_vector(1500, 16),
38411 => conv_std_logic_vector(1650, 16),
38412 => conv_std_logic_vector(1800, 16),
38413 => conv_std_logic_vector(1950, 16),
38414 => conv_std_logic_vector(2100, 16),
38415 => conv_std_logic_vector(2250, 16),
38416 => conv_std_logic_vector(2400, 16),
38417 => conv_std_logic_vector(2550, 16),
38418 => conv_std_logic_vector(2700, 16),
38419 => conv_std_logic_vector(2850, 16),
38420 => conv_std_logic_vector(3000, 16),
38421 => conv_std_logic_vector(3150, 16),
38422 => conv_std_logic_vector(3300, 16),
38423 => conv_std_logic_vector(3450, 16),
38424 => conv_std_logic_vector(3600, 16),
38425 => conv_std_logic_vector(3750, 16),
38426 => conv_std_logic_vector(3900, 16),
38427 => conv_std_logic_vector(4050, 16),
38428 => conv_std_logic_vector(4200, 16),
38429 => conv_std_logic_vector(4350, 16),
38430 => conv_std_logic_vector(4500, 16),
38431 => conv_std_logic_vector(4650, 16),
38432 => conv_std_logic_vector(4800, 16),
38433 => conv_std_logic_vector(4950, 16),
38434 => conv_std_logic_vector(5100, 16),
38435 => conv_std_logic_vector(5250, 16),
38436 => conv_std_logic_vector(5400, 16),
38437 => conv_std_logic_vector(5550, 16),
38438 => conv_std_logic_vector(5700, 16),
38439 => conv_std_logic_vector(5850, 16),
38440 => conv_std_logic_vector(6000, 16),
38441 => conv_std_logic_vector(6150, 16),
38442 => conv_std_logic_vector(6300, 16),
38443 => conv_std_logic_vector(6450, 16),
38444 => conv_std_logic_vector(6600, 16),
38445 => conv_std_logic_vector(6750, 16),
38446 => conv_std_logic_vector(6900, 16),
38447 => conv_std_logic_vector(7050, 16),
38448 => conv_std_logic_vector(7200, 16),
38449 => conv_std_logic_vector(7350, 16),
38450 => conv_std_logic_vector(7500, 16),
38451 => conv_std_logic_vector(7650, 16),
38452 => conv_std_logic_vector(7800, 16),
38453 => conv_std_logic_vector(7950, 16),
38454 => conv_std_logic_vector(8100, 16),
38455 => conv_std_logic_vector(8250, 16),
38456 => conv_std_logic_vector(8400, 16),
38457 => conv_std_logic_vector(8550, 16),
38458 => conv_std_logic_vector(8700, 16),
38459 => conv_std_logic_vector(8850, 16),
38460 => conv_std_logic_vector(9000, 16),
38461 => conv_std_logic_vector(9150, 16),
38462 => conv_std_logic_vector(9300, 16),
38463 => conv_std_logic_vector(9450, 16),
38464 => conv_std_logic_vector(9600, 16),
38465 => conv_std_logic_vector(9750, 16),
38466 => conv_std_logic_vector(9900, 16),
38467 => conv_std_logic_vector(10050, 16),
38468 => conv_std_logic_vector(10200, 16),
38469 => conv_std_logic_vector(10350, 16),
38470 => conv_std_logic_vector(10500, 16),
38471 => conv_std_logic_vector(10650, 16),
38472 => conv_std_logic_vector(10800, 16),
38473 => conv_std_logic_vector(10950, 16),
38474 => conv_std_logic_vector(11100, 16),
38475 => conv_std_logic_vector(11250, 16),
38476 => conv_std_logic_vector(11400, 16),
38477 => conv_std_logic_vector(11550, 16),
38478 => conv_std_logic_vector(11700, 16),
38479 => conv_std_logic_vector(11850, 16),
38480 => conv_std_logic_vector(12000, 16),
38481 => conv_std_logic_vector(12150, 16),
38482 => conv_std_logic_vector(12300, 16),
38483 => conv_std_logic_vector(12450, 16),
38484 => conv_std_logic_vector(12600, 16),
38485 => conv_std_logic_vector(12750, 16),
38486 => conv_std_logic_vector(12900, 16),
38487 => conv_std_logic_vector(13050, 16),
38488 => conv_std_logic_vector(13200, 16),
38489 => conv_std_logic_vector(13350, 16),
38490 => conv_std_logic_vector(13500, 16),
38491 => conv_std_logic_vector(13650, 16),
38492 => conv_std_logic_vector(13800, 16),
38493 => conv_std_logic_vector(13950, 16),
38494 => conv_std_logic_vector(14100, 16),
38495 => conv_std_logic_vector(14250, 16),
38496 => conv_std_logic_vector(14400, 16),
38497 => conv_std_logic_vector(14550, 16),
38498 => conv_std_logic_vector(14700, 16),
38499 => conv_std_logic_vector(14850, 16),
38500 => conv_std_logic_vector(15000, 16),
38501 => conv_std_logic_vector(15150, 16),
38502 => conv_std_logic_vector(15300, 16),
38503 => conv_std_logic_vector(15450, 16),
38504 => conv_std_logic_vector(15600, 16),
38505 => conv_std_logic_vector(15750, 16),
38506 => conv_std_logic_vector(15900, 16),
38507 => conv_std_logic_vector(16050, 16),
38508 => conv_std_logic_vector(16200, 16),
38509 => conv_std_logic_vector(16350, 16),
38510 => conv_std_logic_vector(16500, 16),
38511 => conv_std_logic_vector(16650, 16),
38512 => conv_std_logic_vector(16800, 16),
38513 => conv_std_logic_vector(16950, 16),
38514 => conv_std_logic_vector(17100, 16),
38515 => conv_std_logic_vector(17250, 16),
38516 => conv_std_logic_vector(17400, 16),
38517 => conv_std_logic_vector(17550, 16),
38518 => conv_std_logic_vector(17700, 16),
38519 => conv_std_logic_vector(17850, 16),
38520 => conv_std_logic_vector(18000, 16),
38521 => conv_std_logic_vector(18150, 16),
38522 => conv_std_logic_vector(18300, 16),
38523 => conv_std_logic_vector(18450, 16),
38524 => conv_std_logic_vector(18600, 16),
38525 => conv_std_logic_vector(18750, 16),
38526 => conv_std_logic_vector(18900, 16),
38527 => conv_std_logic_vector(19050, 16),
38528 => conv_std_logic_vector(19200, 16),
38529 => conv_std_logic_vector(19350, 16),
38530 => conv_std_logic_vector(19500, 16),
38531 => conv_std_logic_vector(19650, 16),
38532 => conv_std_logic_vector(19800, 16),
38533 => conv_std_logic_vector(19950, 16),
38534 => conv_std_logic_vector(20100, 16),
38535 => conv_std_logic_vector(20250, 16),
38536 => conv_std_logic_vector(20400, 16),
38537 => conv_std_logic_vector(20550, 16),
38538 => conv_std_logic_vector(20700, 16),
38539 => conv_std_logic_vector(20850, 16),
38540 => conv_std_logic_vector(21000, 16),
38541 => conv_std_logic_vector(21150, 16),
38542 => conv_std_logic_vector(21300, 16),
38543 => conv_std_logic_vector(21450, 16),
38544 => conv_std_logic_vector(21600, 16),
38545 => conv_std_logic_vector(21750, 16),
38546 => conv_std_logic_vector(21900, 16),
38547 => conv_std_logic_vector(22050, 16),
38548 => conv_std_logic_vector(22200, 16),
38549 => conv_std_logic_vector(22350, 16),
38550 => conv_std_logic_vector(22500, 16),
38551 => conv_std_logic_vector(22650, 16),
38552 => conv_std_logic_vector(22800, 16),
38553 => conv_std_logic_vector(22950, 16),
38554 => conv_std_logic_vector(23100, 16),
38555 => conv_std_logic_vector(23250, 16),
38556 => conv_std_logic_vector(23400, 16),
38557 => conv_std_logic_vector(23550, 16),
38558 => conv_std_logic_vector(23700, 16),
38559 => conv_std_logic_vector(23850, 16),
38560 => conv_std_logic_vector(24000, 16),
38561 => conv_std_logic_vector(24150, 16),
38562 => conv_std_logic_vector(24300, 16),
38563 => conv_std_logic_vector(24450, 16),
38564 => conv_std_logic_vector(24600, 16),
38565 => conv_std_logic_vector(24750, 16),
38566 => conv_std_logic_vector(24900, 16),
38567 => conv_std_logic_vector(25050, 16),
38568 => conv_std_logic_vector(25200, 16),
38569 => conv_std_logic_vector(25350, 16),
38570 => conv_std_logic_vector(25500, 16),
38571 => conv_std_logic_vector(25650, 16),
38572 => conv_std_logic_vector(25800, 16),
38573 => conv_std_logic_vector(25950, 16),
38574 => conv_std_logic_vector(26100, 16),
38575 => conv_std_logic_vector(26250, 16),
38576 => conv_std_logic_vector(26400, 16),
38577 => conv_std_logic_vector(26550, 16),
38578 => conv_std_logic_vector(26700, 16),
38579 => conv_std_logic_vector(26850, 16),
38580 => conv_std_logic_vector(27000, 16),
38581 => conv_std_logic_vector(27150, 16),
38582 => conv_std_logic_vector(27300, 16),
38583 => conv_std_logic_vector(27450, 16),
38584 => conv_std_logic_vector(27600, 16),
38585 => conv_std_logic_vector(27750, 16),
38586 => conv_std_logic_vector(27900, 16),
38587 => conv_std_logic_vector(28050, 16),
38588 => conv_std_logic_vector(28200, 16),
38589 => conv_std_logic_vector(28350, 16),
38590 => conv_std_logic_vector(28500, 16),
38591 => conv_std_logic_vector(28650, 16),
38592 => conv_std_logic_vector(28800, 16),
38593 => conv_std_logic_vector(28950, 16),
38594 => conv_std_logic_vector(29100, 16),
38595 => conv_std_logic_vector(29250, 16),
38596 => conv_std_logic_vector(29400, 16),
38597 => conv_std_logic_vector(29550, 16),
38598 => conv_std_logic_vector(29700, 16),
38599 => conv_std_logic_vector(29850, 16),
38600 => conv_std_logic_vector(30000, 16),
38601 => conv_std_logic_vector(30150, 16),
38602 => conv_std_logic_vector(30300, 16),
38603 => conv_std_logic_vector(30450, 16),
38604 => conv_std_logic_vector(30600, 16),
38605 => conv_std_logic_vector(30750, 16),
38606 => conv_std_logic_vector(30900, 16),
38607 => conv_std_logic_vector(31050, 16),
38608 => conv_std_logic_vector(31200, 16),
38609 => conv_std_logic_vector(31350, 16),
38610 => conv_std_logic_vector(31500, 16),
38611 => conv_std_logic_vector(31650, 16),
38612 => conv_std_logic_vector(31800, 16),
38613 => conv_std_logic_vector(31950, 16),
38614 => conv_std_logic_vector(32100, 16),
38615 => conv_std_logic_vector(32250, 16),
38616 => conv_std_logic_vector(32400, 16),
38617 => conv_std_logic_vector(32550, 16),
38618 => conv_std_logic_vector(32700, 16),
38619 => conv_std_logic_vector(32850, 16),
38620 => conv_std_logic_vector(33000, 16),
38621 => conv_std_logic_vector(33150, 16),
38622 => conv_std_logic_vector(33300, 16),
38623 => conv_std_logic_vector(33450, 16),
38624 => conv_std_logic_vector(33600, 16),
38625 => conv_std_logic_vector(33750, 16),
38626 => conv_std_logic_vector(33900, 16),
38627 => conv_std_logic_vector(34050, 16),
38628 => conv_std_logic_vector(34200, 16),
38629 => conv_std_logic_vector(34350, 16),
38630 => conv_std_logic_vector(34500, 16),
38631 => conv_std_logic_vector(34650, 16),
38632 => conv_std_logic_vector(34800, 16),
38633 => conv_std_logic_vector(34950, 16),
38634 => conv_std_logic_vector(35100, 16),
38635 => conv_std_logic_vector(35250, 16),
38636 => conv_std_logic_vector(35400, 16),
38637 => conv_std_logic_vector(35550, 16),
38638 => conv_std_logic_vector(35700, 16),
38639 => conv_std_logic_vector(35850, 16),
38640 => conv_std_logic_vector(36000, 16),
38641 => conv_std_logic_vector(36150, 16),
38642 => conv_std_logic_vector(36300, 16),
38643 => conv_std_logic_vector(36450, 16),
38644 => conv_std_logic_vector(36600, 16),
38645 => conv_std_logic_vector(36750, 16),
38646 => conv_std_logic_vector(36900, 16),
38647 => conv_std_logic_vector(37050, 16),
38648 => conv_std_logic_vector(37200, 16),
38649 => conv_std_logic_vector(37350, 16),
38650 => conv_std_logic_vector(37500, 16),
38651 => conv_std_logic_vector(37650, 16),
38652 => conv_std_logic_vector(37800, 16),
38653 => conv_std_logic_vector(37950, 16),
38654 => conv_std_logic_vector(38100, 16),
38655 => conv_std_logic_vector(38250, 16),
38656 => conv_std_logic_vector(0, 16),
38657 => conv_std_logic_vector(151, 16),
38658 => conv_std_logic_vector(302, 16),
38659 => conv_std_logic_vector(453, 16),
38660 => conv_std_logic_vector(604, 16),
38661 => conv_std_logic_vector(755, 16),
38662 => conv_std_logic_vector(906, 16),
38663 => conv_std_logic_vector(1057, 16),
38664 => conv_std_logic_vector(1208, 16),
38665 => conv_std_logic_vector(1359, 16),
38666 => conv_std_logic_vector(1510, 16),
38667 => conv_std_logic_vector(1661, 16),
38668 => conv_std_logic_vector(1812, 16),
38669 => conv_std_logic_vector(1963, 16),
38670 => conv_std_logic_vector(2114, 16),
38671 => conv_std_logic_vector(2265, 16),
38672 => conv_std_logic_vector(2416, 16),
38673 => conv_std_logic_vector(2567, 16),
38674 => conv_std_logic_vector(2718, 16),
38675 => conv_std_logic_vector(2869, 16),
38676 => conv_std_logic_vector(3020, 16),
38677 => conv_std_logic_vector(3171, 16),
38678 => conv_std_logic_vector(3322, 16),
38679 => conv_std_logic_vector(3473, 16),
38680 => conv_std_logic_vector(3624, 16),
38681 => conv_std_logic_vector(3775, 16),
38682 => conv_std_logic_vector(3926, 16),
38683 => conv_std_logic_vector(4077, 16),
38684 => conv_std_logic_vector(4228, 16),
38685 => conv_std_logic_vector(4379, 16),
38686 => conv_std_logic_vector(4530, 16),
38687 => conv_std_logic_vector(4681, 16),
38688 => conv_std_logic_vector(4832, 16),
38689 => conv_std_logic_vector(4983, 16),
38690 => conv_std_logic_vector(5134, 16),
38691 => conv_std_logic_vector(5285, 16),
38692 => conv_std_logic_vector(5436, 16),
38693 => conv_std_logic_vector(5587, 16),
38694 => conv_std_logic_vector(5738, 16),
38695 => conv_std_logic_vector(5889, 16),
38696 => conv_std_logic_vector(6040, 16),
38697 => conv_std_logic_vector(6191, 16),
38698 => conv_std_logic_vector(6342, 16),
38699 => conv_std_logic_vector(6493, 16),
38700 => conv_std_logic_vector(6644, 16),
38701 => conv_std_logic_vector(6795, 16),
38702 => conv_std_logic_vector(6946, 16),
38703 => conv_std_logic_vector(7097, 16),
38704 => conv_std_logic_vector(7248, 16),
38705 => conv_std_logic_vector(7399, 16),
38706 => conv_std_logic_vector(7550, 16),
38707 => conv_std_logic_vector(7701, 16),
38708 => conv_std_logic_vector(7852, 16),
38709 => conv_std_logic_vector(8003, 16),
38710 => conv_std_logic_vector(8154, 16),
38711 => conv_std_logic_vector(8305, 16),
38712 => conv_std_logic_vector(8456, 16),
38713 => conv_std_logic_vector(8607, 16),
38714 => conv_std_logic_vector(8758, 16),
38715 => conv_std_logic_vector(8909, 16),
38716 => conv_std_logic_vector(9060, 16),
38717 => conv_std_logic_vector(9211, 16),
38718 => conv_std_logic_vector(9362, 16),
38719 => conv_std_logic_vector(9513, 16),
38720 => conv_std_logic_vector(9664, 16),
38721 => conv_std_logic_vector(9815, 16),
38722 => conv_std_logic_vector(9966, 16),
38723 => conv_std_logic_vector(10117, 16),
38724 => conv_std_logic_vector(10268, 16),
38725 => conv_std_logic_vector(10419, 16),
38726 => conv_std_logic_vector(10570, 16),
38727 => conv_std_logic_vector(10721, 16),
38728 => conv_std_logic_vector(10872, 16),
38729 => conv_std_logic_vector(11023, 16),
38730 => conv_std_logic_vector(11174, 16),
38731 => conv_std_logic_vector(11325, 16),
38732 => conv_std_logic_vector(11476, 16),
38733 => conv_std_logic_vector(11627, 16),
38734 => conv_std_logic_vector(11778, 16),
38735 => conv_std_logic_vector(11929, 16),
38736 => conv_std_logic_vector(12080, 16),
38737 => conv_std_logic_vector(12231, 16),
38738 => conv_std_logic_vector(12382, 16),
38739 => conv_std_logic_vector(12533, 16),
38740 => conv_std_logic_vector(12684, 16),
38741 => conv_std_logic_vector(12835, 16),
38742 => conv_std_logic_vector(12986, 16),
38743 => conv_std_logic_vector(13137, 16),
38744 => conv_std_logic_vector(13288, 16),
38745 => conv_std_logic_vector(13439, 16),
38746 => conv_std_logic_vector(13590, 16),
38747 => conv_std_logic_vector(13741, 16),
38748 => conv_std_logic_vector(13892, 16),
38749 => conv_std_logic_vector(14043, 16),
38750 => conv_std_logic_vector(14194, 16),
38751 => conv_std_logic_vector(14345, 16),
38752 => conv_std_logic_vector(14496, 16),
38753 => conv_std_logic_vector(14647, 16),
38754 => conv_std_logic_vector(14798, 16),
38755 => conv_std_logic_vector(14949, 16),
38756 => conv_std_logic_vector(15100, 16),
38757 => conv_std_logic_vector(15251, 16),
38758 => conv_std_logic_vector(15402, 16),
38759 => conv_std_logic_vector(15553, 16),
38760 => conv_std_logic_vector(15704, 16),
38761 => conv_std_logic_vector(15855, 16),
38762 => conv_std_logic_vector(16006, 16),
38763 => conv_std_logic_vector(16157, 16),
38764 => conv_std_logic_vector(16308, 16),
38765 => conv_std_logic_vector(16459, 16),
38766 => conv_std_logic_vector(16610, 16),
38767 => conv_std_logic_vector(16761, 16),
38768 => conv_std_logic_vector(16912, 16),
38769 => conv_std_logic_vector(17063, 16),
38770 => conv_std_logic_vector(17214, 16),
38771 => conv_std_logic_vector(17365, 16),
38772 => conv_std_logic_vector(17516, 16),
38773 => conv_std_logic_vector(17667, 16),
38774 => conv_std_logic_vector(17818, 16),
38775 => conv_std_logic_vector(17969, 16),
38776 => conv_std_logic_vector(18120, 16),
38777 => conv_std_logic_vector(18271, 16),
38778 => conv_std_logic_vector(18422, 16),
38779 => conv_std_logic_vector(18573, 16),
38780 => conv_std_logic_vector(18724, 16),
38781 => conv_std_logic_vector(18875, 16),
38782 => conv_std_logic_vector(19026, 16),
38783 => conv_std_logic_vector(19177, 16),
38784 => conv_std_logic_vector(19328, 16),
38785 => conv_std_logic_vector(19479, 16),
38786 => conv_std_logic_vector(19630, 16),
38787 => conv_std_logic_vector(19781, 16),
38788 => conv_std_logic_vector(19932, 16),
38789 => conv_std_logic_vector(20083, 16),
38790 => conv_std_logic_vector(20234, 16),
38791 => conv_std_logic_vector(20385, 16),
38792 => conv_std_logic_vector(20536, 16),
38793 => conv_std_logic_vector(20687, 16),
38794 => conv_std_logic_vector(20838, 16),
38795 => conv_std_logic_vector(20989, 16),
38796 => conv_std_logic_vector(21140, 16),
38797 => conv_std_logic_vector(21291, 16),
38798 => conv_std_logic_vector(21442, 16),
38799 => conv_std_logic_vector(21593, 16),
38800 => conv_std_logic_vector(21744, 16),
38801 => conv_std_logic_vector(21895, 16),
38802 => conv_std_logic_vector(22046, 16),
38803 => conv_std_logic_vector(22197, 16),
38804 => conv_std_logic_vector(22348, 16),
38805 => conv_std_logic_vector(22499, 16),
38806 => conv_std_logic_vector(22650, 16),
38807 => conv_std_logic_vector(22801, 16),
38808 => conv_std_logic_vector(22952, 16),
38809 => conv_std_logic_vector(23103, 16),
38810 => conv_std_logic_vector(23254, 16),
38811 => conv_std_logic_vector(23405, 16),
38812 => conv_std_logic_vector(23556, 16),
38813 => conv_std_logic_vector(23707, 16),
38814 => conv_std_logic_vector(23858, 16),
38815 => conv_std_logic_vector(24009, 16),
38816 => conv_std_logic_vector(24160, 16),
38817 => conv_std_logic_vector(24311, 16),
38818 => conv_std_logic_vector(24462, 16),
38819 => conv_std_logic_vector(24613, 16),
38820 => conv_std_logic_vector(24764, 16),
38821 => conv_std_logic_vector(24915, 16),
38822 => conv_std_logic_vector(25066, 16),
38823 => conv_std_logic_vector(25217, 16),
38824 => conv_std_logic_vector(25368, 16),
38825 => conv_std_logic_vector(25519, 16),
38826 => conv_std_logic_vector(25670, 16),
38827 => conv_std_logic_vector(25821, 16),
38828 => conv_std_logic_vector(25972, 16),
38829 => conv_std_logic_vector(26123, 16),
38830 => conv_std_logic_vector(26274, 16),
38831 => conv_std_logic_vector(26425, 16),
38832 => conv_std_logic_vector(26576, 16),
38833 => conv_std_logic_vector(26727, 16),
38834 => conv_std_logic_vector(26878, 16),
38835 => conv_std_logic_vector(27029, 16),
38836 => conv_std_logic_vector(27180, 16),
38837 => conv_std_logic_vector(27331, 16),
38838 => conv_std_logic_vector(27482, 16),
38839 => conv_std_logic_vector(27633, 16),
38840 => conv_std_logic_vector(27784, 16),
38841 => conv_std_logic_vector(27935, 16),
38842 => conv_std_logic_vector(28086, 16),
38843 => conv_std_logic_vector(28237, 16),
38844 => conv_std_logic_vector(28388, 16),
38845 => conv_std_logic_vector(28539, 16),
38846 => conv_std_logic_vector(28690, 16),
38847 => conv_std_logic_vector(28841, 16),
38848 => conv_std_logic_vector(28992, 16),
38849 => conv_std_logic_vector(29143, 16),
38850 => conv_std_logic_vector(29294, 16),
38851 => conv_std_logic_vector(29445, 16),
38852 => conv_std_logic_vector(29596, 16),
38853 => conv_std_logic_vector(29747, 16),
38854 => conv_std_logic_vector(29898, 16),
38855 => conv_std_logic_vector(30049, 16),
38856 => conv_std_logic_vector(30200, 16),
38857 => conv_std_logic_vector(30351, 16),
38858 => conv_std_logic_vector(30502, 16),
38859 => conv_std_logic_vector(30653, 16),
38860 => conv_std_logic_vector(30804, 16),
38861 => conv_std_logic_vector(30955, 16),
38862 => conv_std_logic_vector(31106, 16),
38863 => conv_std_logic_vector(31257, 16),
38864 => conv_std_logic_vector(31408, 16),
38865 => conv_std_logic_vector(31559, 16),
38866 => conv_std_logic_vector(31710, 16),
38867 => conv_std_logic_vector(31861, 16),
38868 => conv_std_logic_vector(32012, 16),
38869 => conv_std_logic_vector(32163, 16),
38870 => conv_std_logic_vector(32314, 16),
38871 => conv_std_logic_vector(32465, 16),
38872 => conv_std_logic_vector(32616, 16),
38873 => conv_std_logic_vector(32767, 16),
38874 => conv_std_logic_vector(32918, 16),
38875 => conv_std_logic_vector(33069, 16),
38876 => conv_std_logic_vector(33220, 16),
38877 => conv_std_logic_vector(33371, 16),
38878 => conv_std_logic_vector(33522, 16),
38879 => conv_std_logic_vector(33673, 16),
38880 => conv_std_logic_vector(33824, 16),
38881 => conv_std_logic_vector(33975, 16),
38882 => conv_std_logic_vector(34126, 16),
38883 => conv_std_logic_vector(34277, 16),
38884 => conv_std_logic_vector(34428, 16),
38885 => conv_std_logic_vector(34579, 16),
38886 => conv_std_logic_vector(34730, 16),
38887 => conv_std_logic_vector(34881, 16),
38888 => conv_std_logic_vector(35032, 16),
38889 => conv_std_logic_vector(35183, 16),
38890 => conv_std_logic_vector(35334, 16),
38891 => conv_std_logic_vector(35485, 16),
38892 => conv_std_logic_vector(35636, 16),
38893 => conv_std_logic_vector(35787, 16),
38894 => conv_std_logic_vector(35938, 16),
38895 => conv_std_logic_vector(36089, 16),
38896 => conv_std_logic_vector(36240, 16),
38897 => conv_std_logic_vector(36391, 16),
38898 => conv_std_logic_vector(36542, 16),
38899 => conv_std_logic_vector(36693, 16),
38900 => conv_std_logic_vector(36844, 16),
38901 => conv_std_logic_vector(36995, 16),
38902 => conv_std_logic_vector(37146, 16),
38903 => conv_std_logic_vector(37297, 16),
38904 => conv_std_logic_vector(37448, 16),
38905 => conv_std_logic_vector(37599, 16),
38906 => conv_std_logic_vector(37750, 16),
38907 => conv_std_logic_vector(37901, 16),
38908 => conv_std_logic_vector(38052, 16),
38909 => conv_std_logic_vector(38203, 16),
38910 => conv_std_logic_vector(38354, 16),
38911 => conv_std_logic_vector(38505, 16),
38912 => conv_std_logic_vector(0, 16),
38913 => conv_std_logic_vector(152, 16),
38914 => conv_std_logic_vector(304, 16),
38915 => conv_std_logic_vector(456, 16),
38916 => conv_std_logic_vector(608, 16),
38917 => conv_std_logic_vector(760, 16),
38918 => conv_std_logic_vector(912, 16),
38919 => conv_std_logic_vector(1064, 16),
38920 => conv_std_logic_vector(1216, 16),
38921 => conv_std_logic_vector(1368, 16),
38922 => conv_std_logic_vector(1520, 16),
38923 => conv_std_logic_vector(1672, 16),
38924 => conv_std_logic_vector(1824, 16),
38925 => conv_std_logic_vector(1976, 16),
38926 => conv_std_logic_vector(2128, 16),
38927 => conv_std_logic_vector(2280, 16),
38928 => conv_std_logic_vector(2432, 16),
38929 => conv_std_logic_vector(2584, 16),
38930 => conv_std_logic_vector(2736, 16),
38931 => conv_std_logic_vector(2888, 16),
38932 => conv_std_logic_vector(3040, 16),
38933 => conv_std_logic_vector(3192, 16),
38934 => conv_std_logic_vector(3344, 16),
38935 => conv_std_logic_vector(3496, 16),
38936 => conv_std_logic_vector(3648, 16),
38937 => conv_std_logic_vector(3800, 16),
38938 => conv_std_logic_vector(3952, 16),
38939 => conv_std_logic_vector(4104, 16),
38940 => conv_std_logic_vector(4256, 16),
38941 => conv_std_logic_vector(4408, 16),
38942 => conv_std_logic_vector(4560, 16),
38943 => conv_std_logic_vector(4712, 16),
38944 => conv_std_logic_vector(4864, 16),
38945 => conv_std_logic_vector(5016, 16),
38946 => conv_std_logic_vector(5168, 16),
38947 => conv_std_logic_vector(5320, 16),
38948 => conv_std_logic_vector(5472, 16),
38949 => conv_std_logic_vector(5624, 16),
38950 => conv_std_logic_vector(5776, 16),
38951 => conv_std_logic_vector(5928, 16),
38952 => conv_std_logic_vector(6080, 16),
38953 => conv_std_logic_vector(6232, 16),
38954 => conv_std_logic_vector(6384, 16),
38955 => conv_std_logic_vector(6536, 16),
38956 => conv_std_logic_vector(6688, 16),
38957 => conv_std_logic_vector(6840, 16),
38958 => conv_std_logic_vector(6992, 16),
38959 => conv_std_logic_vector(7144, 16),
38960 => conv_std_logic_vector(7296, 16),
38961 => conv_std_logic_vector(7448, 16),
38962 => conv_std_logic_vector(7600, 16),
38963 => conv_std_logic_vector(7752, 16),
38964 => conv_std_logic_vector(7904, 16),
38965 => conv_std_logic_vector(8056, 16),
38966 => conv_std_logic_vector(8208, 16),
38967 => conv_std_logic_vector(8360, 16),
38968 => conv_std_logic_vector(8512, 16),
38969 => conv_std_logic_vector(8664, 16),
38970 => conv_std_logic_vector(8816, 16),
38971 => conv_std_logic_vector(8968, 16),
38972 => conv_std_logic_vector(9120, 16),
38973 => conv_std_logic_vector(9272, 16),
38974 => conv_std_logic_vector(9424, 16),
38975 => conv_std_logic_vector(9576, 16),
38976 => conv_std_logic_vector(9728, 16),
38977 => conv_std_logic_vector(9880, 16),
38978 => conv_std_logic_vector(10032, 16),
38979 => conv_std_logic_vector(10184, 16),
38980 => conv_std_logic_vector(10336, 16),
38981 => conv_std_logic_vector(10488, 16),
38982 => conv_std_logic_vector(10640, 16),
38983 => conv_std_logic_vector(10792, 16),
38984 => conv_std_logic_vector(10944, 16),
38985 => conv_std_logic_vector(11096, 16),
38986 => conv_std_logic_vector(11248, 16),
38987 => conv_std_logic_vector(11400, 16),
38988 => conv_std_logic_vector(11552, 16),
38989 => conv_std_logic_vector(11704, 16),
38990 => conv_std_logic_vector(11856, 16),
38991 => conv_std_logic_vector(12008, 16),
38992 => conv_std_logic_vector(12160, 16),
38993 => conv_std_logic_vector(12312, 16),
38994 => conv_std_logic_vector(12464, 16),
38995 => conv_std_logic_vector(12616, 16),
38996 => conv_std_logic_vector(12768, 16),
38997 => conv_std_logic_vector(12920, 16),
38998 => conv_std_logic_vector(13072, 16),
38999 => conv_std_logic_vector(13224, 16),
39000 => conv_std_logic_vector(13376, 16),
39001 => conv_std_logic_vector(13528, 16),
39002 => conv_std_logic_vector(13680, 16),
39003 => conv_std_logic_vector(13832, 16),
39004 => conv_std_logic_vector(13984, 16),
39005 => conv_std_logic_vector(14136, 16),
39006 => conv_std_logic_vector(14288, 16),
39007 => conv_std_logic_vector(14440, 16),
39008 => conv_std_logic_vector(14592, 16),
39009 => conv_std_logic_vector(14744, 16),
39010 => conv_std_logic_vector(14896, 16),
39011 => conv_std_logic_vector(15048, 16),
39012 => conv_std_logic_vector(15200, 16),
39013 => conv_std_logic_vector(15352, 16),
39014 => conv_std_logic_vector(15504, 16),
39015 => conv_std_logic_vector(15656, 16),
39016 => conv_std_logic_vector(15808, 16),
39017 => conv_std_logic_vector(15960, 16),
39018 => conv_std_logic_vector(16112, 16),
39019 => conv_std_logic_vector(16264, 16),
39020 => conv_std_logic_vector(16416, 16),
39021 => conv_std_logic_vector(16568, 16),
39022 => conv_std_logic_vector(16720, 16),
39023 => conv_std_logic_vector(16872, 16),
39024 => conv_std_logic_vector(17024, 16),
39025 => conv_std_logic_vector(17176, 16),
39026 => conv_std_logic_vector(17328, 16),
39027 => conv_std_logic_vector(17480, 16),
39028 => conv_std_logic_vector(17632, 16),
39029 => conv_std_logic_vector(17784, 16),
39030 => conv_std_logic_vector(17936, 16),
39031 => conv_std_logic_vector(18088, 16),
39032 => conv_std_logic_vector(18240, 16),
39033 => conv_std_logic_vector(18392, 16),
39034 => conv_std_logic_vector(18544, 16),
39035 => conv_std_logic_vector(18696, 16),
39036 => conv_std_logic_vector(18848, 16),
39037 => conv_std_logic_vector(19000, 16),
39038 => conv_std_logic_vector(19152, 16),
39039 => conv_std_logic_vector(19304, 16),
39040 => conv_std_logic_vector(19456, 16),
39041 => conv_std_logic_vector(19608, 16),
39042 => conv_std_logic_vector(19760, 16),
39043 => conv_std_logic_vector(19912, 16),
39044 => conv_std_logic_vector(20064, 16),
39045 => conv_std_logic_vector(20216, 16),
39046 => conv_std_logic_vector(20368, 16),
39047 => conv_std_logic_vector(20520, 16),
39048 => conv_std_logic_vector(20672, 16),
39049 => conv_std_logic_vector(20824, 16),
39050 => conv_std_logic_vector(20976, 16),
39051 => conv_std_logic_vector(21128, 16),
39052 => conv_std_logic_vector(21280, 16),
39053 => conv_std_logic_vector(21432, 16),
39054 => conv_std_logic_vector(21584, 16),
39055 => conv_std_logic_vector(21736, 16),
39056 => conv_std_logic_vector(21888, 16),
39057 => conv_std_logic_vector(22040, 16),
39058 => conv_std_logic_vector(22192, 16),
39059 => conv_std_logic_vector(22344, 16),
39060 => conv_std_logic_vector(22496, 16),
39061 => conv_std_logic_vector(22648, 16),
39062 => conv_std_logic_vector(22800, 16),
39063 => conv_std_logic_vector(22952, 16),
39064 => conv_std_logic_vector(23104, 16),
39065 => conv_std_logic_vector(23256, 16),
39066 => conv_std_logic_vector(23408, 16),
39067 => conv_std_logic_vector(23560, 16),
39068 => conv_std_logic_vector(23712, 16),
39069 => conv_std_logic_vector(23864, 16),
39070 => conv_std_logic_vector(24016, 16),
39071 => conv_std_logic_vector(24168, 16),
39072 => conv_std_logic_vector(24320, 16),
39073 => conv_std_logic_vector(24472, 16),
39074 => conv_std_logic_vector(24624, 16),
39075 => conv_std_logic_vector(24776, 16),
39076 => conv_std_logic_vector(24928, 16),
39077 => conv_std_logic_vector(25080, 16),
39078 => conv_std_logic_vector(25232, 16),
39079 => conv_std_logic_vector(25384, 16),
39080 => conv_std_logic_vector(25536, 16),
39081 => conv_std_logic_vector(25688, 16),
39082 => conv_std_logic_vector(25840, 16),
39083 => conv_std_logic_vector(25992, 16),
39084 => conv_std_logic_vector(26144, 16),
39085 => conv_std_logic_vector(26296, 16),
39086 => conv_std_logic_vector(26448, 16),
39087 => conv_std_logic_vector(26600, 16),
39088 => conv_std_logic_vector(26752, 16),
39089 => conv_std_logic_vector(26904, 16),
39090 => conv_std_logic_vector(27056, 16),
39091 => conv_std_logic_vector(27208, 16),
39092 => conv_std_logic_vector(27360, 16),
39093 => conv_std_logic_vector(27512, 16),
39094 => conv_std_logic_vector(27664, 16),
39095 => conv_std_logic_vector(27816, 16),
39096 => conv_std_logic_vector(27968, 16),
39097 => conv_std_logic_vector(28120, 16),
39098 => conv_std_logic_vector(28272, 16),
39099 => conv_std_logic_vector(28424, 16),
39100 => conv_std_logic_vector(28576, 16),
39101 => conv_std_logic_vector(28728, 16),
39102 => conv_std_logic_vector(28880, 16),
39103 => conv_std_logic_vector(29032, 16),
39104 => conv_std_logic_vector(29184, 16),
39105 => conv_std_logic_vector(29336, 16),
39106 => conv_std_logic_vector(29488, 16),
39107 => conv_std_logic_vector(29640, 16),
39108 => conv_std_logic_vector(29792, 16),
39109 => conv_std_logic_vector(29944, 16),
39110 => conv_std_logic_vector(30096, 16),
39111 => conv_std_logic_vector(30248, 16),
39112 => conv_std_logic_vector(30400, 16),
39113 => conv_std_logic_vector(30552, 16),
39114 => conv_std_logic_vector(30704, 16),
39115 => conv_std_logic_vector(30856, 16),
39116 => conv_std_logic_vector(31008, 16),
39117 => conv_std_logic_vector(31160, 16),
39118 => conv_std_logic_vector(31312, 16),
39119 => conv_std_logic_vector(31464, 16),
39120 => conv_std_logic_vector(31616, 16),
39121 => conv_std_logic_vector(31768, 16),
39122 => conv_std_logic_vector(31920, 16),
39123 => conv_std_logic_vector(32072, 16),
39124 => conv_std_logic_vector(32224, 16),
39125 => conv_std_logic_vector(32376, 16),
39126 => conv_std_logic_vector(32528, 16),
39127 => conv_std_logic_vector(32680, 16),
39128 => conv_std_logic_vector(32832, 16),
39129 => conv_std_logic_vector(32984, 16),
39130 => conv_std_logic_vector(33136, 16),
39131 => conv_std_logic_vector(33288, 16),
39132 => conv_std_logic_vector(33440, 16),
39133 => conv_std_logic_vector(33592, 16),
39134 => conv_std_logic_vector(33744, 16),
39135 => conv_std_logic_vector(33896, 16),
39136 => conv_std_logic_vector(34048, 16),
39137 => conv_std_logic_vector(34200, 16),
39138 => conv_std_logic_vector(34352, 16),
39139 => conv_std_logic_vector(34504, 16),
39140 => conv_std_logic_vector(34656, 16),
39141 => conv_std_logic_vector(34808, 16),
39142 => conv_std_logic_vector(34960, 16),
39143 => conv_std_logic_vector(35112, 16),
39144 => conv_std_logic_vector(35264, 16),
39145 => conv_std_logic_vector(35416, 16),
39146 => conv_std_logic_vector(35568, 16),
39147 => conv_std_logic_vector(35720, 16),
39148 => conv_std_logic_vector(35872, 16),
39149 => conv_std_logic_vector(36024, 16),
39150 => conv_std_logic_vector(36176, 16),
39151 => conv_std_logic_vector(36328, 16),
39152 => conv_std_logic_vector(36480, 16),
39153 => conv_std_logic_vector(36632, 16),
39154 => conv_std_logic_vector(36784, 16),
39155 => conv_std_logic_vector(36936, 16),
39156 => conv_std_logic_vector(37088, 16),
39157 => conv_std_logic_vector(37240, 16),
39158 => conv_std_logic_vector(37392, 16),
39159 => conv_std_logic_vector(37544, 16),
39160 => conv_std_logic_vector(37696, 16),
39161 => conv_std_logic_vector(37848, 16),
39162 => conv_std_logic_vector(38000, 16),
39163 => conv_std_logic_vector(38152, 16),
39164 => conv_std_logic_vector(38304, 16),
39165 => conv_std_logic_vector(38456, 16),
39166 => conv_std_logic_vector(38608, 16),
39167 => conv_std_logic_vector(38760, 16),
39168 => conv_std_logic_vector(0, 16),
39169 => conv_std_logic_vector(153, 16),
39170 => conv_std_logic_vector(306, 16),
39171 => conv_std_logic_vector(459, 16),
39172 => conv_std_logic_vector(612, 16),
39173 => conv_std_logic_vector(765, 16),
39174 => conv_std_logic_vector(918, 16),
39175 => conv_std_logic_vector(1071, 16),
39176 => conv_std_logic_vector(1224, 16),
39177 => conv_std_logic_vector(1377, 16),
39178 => conv_std_logic_vector(1530, 16),
39179 => conv_std_logic_vector(1683, 16),
39180 => conv_std_logic_vector(1836, 16),
39181 => conv_std_logic_vector(1989, 16),
39182 => conv_std_logic_vector(2142, 16),
39183 => conv_std_logic_vector(2295, 16),
39184 => conv_std_logic_vector(2448, 16),
39185 => conv_std_logic_vector(2601, 16),
39186 => conv_std_logic_vector(2754, 16),
39187 => conv_std_logic_vector(2907, 16),
39188 => conv_std_logic_vector(3060, 16),
39189 => conv_std_logic_vector(3213, 16),
39190 => conv_std_logic_vector(3366, 16),
39191 => conv_std_logic_vector(3519, 16),
39192 => conv_std_logic_vector(3672, 16),
39193 => conv_std_logic_vector(3825, 16),
39194 => conv_std_logic_vector(3978, 16),
39195 => conv_std_logic_vector(4131, 16),
39196 => conv_std_logic_vector(4284, 16),
39197 => conv_std_logic_vector(4437, 16),
39198 => conv_std_logic_vector(4590, 16),
39199 => conv_std_logic_vector(4743, 16),
39200 => conv_std_logic_vector(4896, 16),
39201 => conv_std_logic_vector(5049, 16),
39202 => conv_std_logic_vector(5202, 16),
39203 => conv_std_logic_vector(5355, 16),
39204 => conv_std_logic_vector(5508, 16),
39205 => conv_std_logic_vector(5661, 16),
39206 => conv_std_logic_vector(5814, 16),
39207 => conv_std_logic_vector(5967, 16),
39208 => conv_std_logic_vector(6120, 16),
39209 => conv_std_logic_vector(6273, 16),
39210 => conv_std_logic_vector(6426, 16),
39211 => conv_std_logic_vector(6579, 16),
39212 => conv_std_logic_vector(6732, 16),
39213 => conv_std_logic_vector(6885, 16),
39214 => conv_std_logic_vector(7038, 16),
39215 => conv_std_logic_vector(7191, 16),
39216 => conv_std_logic_vector(7344, 16),
39217 => conv_std_logic_vector(7497, 16),
39218 => conv_std_logic_vector(7650, 16),
39219 => conv_std_logic_vector(7803, 16),
39220 => conv_std_logic_vector(7956, 16),
39221 => conv_std_logic_vector(8109, 16),
39222 => conv_std_logic_vector(8262, 16),
39223 => conv_std_logic_vector(8415, 16),
39224 => conv_std_logic_vector(8568, 16),
39225 => conv_std_logic_vector(8721, 16),
39226 => conv_std_logic_vector(8874, 16),
39227 => conv_std_logic_vector(9027, 16),
39228 => conv_std_logic_vector(9180, 16),
39229 => conv_std_logic_vector(9333, 16),
39230 => conv_std_logic_vector(9486, 16),
39231 => conv_std_logic_vector(9639, 16),
39232 => conv_std_logic_vector(9792, 16),
39233 => conv_std_logic_vector(9945, 16),
39234 => conv_std_logic_vector(10098, 16),
39235 => conv_std_logic_vector(10251, 16),
39236 => conv_std_logic_vector(10404, 16),
39237 => conv_std_logic_vector(10557, 16),
39238 => conv_std_logic_vector(10710, 16),
39239 => conv_std_logic_vector(10863, 16),
39240 => conv_std_logic_vector(11016, 16),
39241 => conv_std_logic_vector(11169, 16),
39242 => conv_std_logic_vector(11322, 16),
39243 => conv_std_logic_vector(11475, 16),
39244 => conv_std_logic_vector(11628, 16),
39245 => conv_std_logic_vector(11781, 16),
39246 => conv_std_logic_vector(11934, 16),
39247 => conv_std_logic_vector(12087, 16),
39248 => conv_std_logic_vector(12240, 16),
39249 => conv_std_logic_vector(12393, 16),
39250 => conv_std_logic_vector(12546, 16),
39251 => conv_std_logic_vector(12699, 16),
39252 => conv_std_logic_vector(12852, 16),
39253 => conv_std_logic_vector(13005, 16),
39254 => conv_std_logic_vector(13158, 16),
39255 => conv_std_logic_vector(13311, 16),
39256 => conv_std_logic_vector(13464, 16),
39257 => conv_std_logic_vector(13617, 16),
39258 => conv_std_logic_vector(13770, 16),
39259 => conv_std_logic_vector(13923, 16),
39260 => conv_std_logic_vector(14076, 16),
39261 => conv_std_logic_vector(14229, 16),
39262 => conv_std_logic_vector(14382, 16),
39263 => conv_std_logic_vector(14535, 16),
39264 => conv_std_logic_vector(14688, 16),
39265 => conv_std_logic_vector(14841, 16),
39266 => conv_std_logic_vector(14994, 16),
39267 => conv_std_logic_vector(15147, 16),
39268 => conv_std_logic_vector(15300, 16),
39269 => conv_std_logic_vector(15453, 16),
39270 => conv_std_logic_vector(15606, 16),
39271 => conv_std_logic_vector(15759, 16),
39272 => conv_std_logic_vector(15912, 16),
39273 => conv_std_logic_vector(16065, 16),
39274 => conv_std_logic_vector(16218, 16),
39275 => conv_std_logic_vector(16371, 16),
39276 => conv_std_logic_vector(16524, 16),
39277 => conv_std_logic_vector(16677, 16),
39278 => conv_std_logic_vector(16830, 16),
39279 => conv_std_logic_vector(16983, 16),
39280 => conv_std_logic_vector(17136, 16),
39281 => conv_std_logic_vector(17289, 16),
39282 => conv_std_logic_vector(17442, 16),
39283 => conv_std_logic_vector(17595, 16),
39284 => conv_std_logic_vector(17748, 16),
39285 => conv_std_logic_vector(17901, 16),
39286 => conv_std_logic_vector(18054, 16),
39287 => conv_std_logic_vector(18207, 16),
39288 => conv_std_logic_vector(18360, 16),
39289 => conv_std_logic_vector(18513, 16),
39290 => conv_std_logic_vector(18666, 16),
39291 => conv_std_logic_vector(18819, 16),
39292 => conv_std_logic_vector(18972, 16),
39293 => conv_std_logic_vector(19125, 16),
39294 => conv_std_logic_vector(19278, 16),
39295 => conv_std_logic_vector(19431, 16),
39296 => conv_std_logic_vector(19584, 16),
39297 => conv_std_logic_vector(19737, 16),
39298 => conv_std_logic_vector(19890, 16),
39299 => conv_std_logic_vector(20043, 16),
39300 => conv_std_logic_vector(20196, 16),
39301 => conv_std_logic_vector(20349, 16),
39302 => conv_std_logic_vector(20502, 16),
39303 => conv_std_logic_vector(20655, 16),
39304 => conv_std_logic_vector(20808, 16),
39305 => conv_std_logic_vector(20961, 16),
39306 => conv_std_logic_vector(21114, 16),
39307 => conv_std_logic_vector(21267, 16),
39308 => conv_std_logic_vector(21420, 16),
39309 => conv_std_logic_vector(21573, 16),
39310 => conv_std_logic_vector(21726, 16),
39311 => conv_std_logic_vector(21879, 16),
39312 => conv_std_logic_vector(22032, 16),
39313 => conv_std_logic_vector(22185, 16),
39314 => conv_std_logic_vector(22338, 16),
39315 => conv_std_logic_vector(22491, 16),
39316 => conv_std_logic_vector(22644, 16),
39317 => conv_std_logic_vector(22797, 16),
39318 => conv_std_logic_vector(22950, 16),
39319 => conv_std_logic_vector(23103, 16),
39320 => conv_std_logic_vector(23256, 16),
39321 => conv_std_logic_vector(23409, 16),
39322 => conv_std_logic_vector(23562, 16),
39323 => conv_std_logic_vector(23715, 16),
39324 => conv_std_logic_vector(23868, 16),
39325 => conv_std_logic_vector(24021, 16),
39326 => conv_std_logic_vector(24174, 16),
39327 => conv_std_logic_vector(24327, 16),
39328 => conv_std_logic_vector(24480, 16),
39329 => conv_std_logic_vector(24633, 16),
39330 => conv_std_logic_vector(24786, 16),
39331 => conv_std_logic_vector(24939, 16),
39332 => conv_std_logic_vector(25092, 16),
39333 => conv_std_logic_vector(25245, 16),
39334 => conv_std_logic_vector(25398, 16),
39335 => conv_std_logic_vector(25551, 16),
39336 => conv_std_logic_vector(25704, 16),
39337 => conv_std_logic_vector(25857, 16),
39338 => conv_std_logic_vector(26010, 16),
39339 => conv_std_logic_vector(26163, 16),
39340 => conv_std_logic_vector(26316, 16),
39341 => conv_std_logic_vector(26469, 16),
39342 => conv_std_logic_vector(26622, 16),
39343 => conv_std_logic_vector(26775, 16),
39344 => conv_std_logic_vector(26928, 16),
39345 => conv_std_logic_vector(27081, 16),
39346 => conv_std_logic_vector(27234, 16),
39347 => conv_std_logic_vector(27387, 16),
39348 => conv_std_logic_vector(27540, 16),
39349 => conv_std_logic_vector(27693, 16),
39350 => conv_std_logic_vector(27846, 16),
39351 => conv_std_logic_vector(27999, 16),
39352 => conv_std_logic_vector(28152, 16),
39353 => conv_std_logic_vector(28305, 16),
39354 => conv_std_logic_vector(28458, 16),
39355 => conv_std_logic_vector(28611, 16),
39356 => conv_std_logic_vector(28764, 16),
39357 => conv_std_logic_vector(28917, 16),
39358 => conv_std_logic_vector(29070, 16),
39359 => conv_std_logic_vector(29223, 16),
39360 => conv_std_logic_vector(29376, 16),
39361 => conv_std_logic_vector(29529, 16),
39362 => conv_std_logic_vector(29682, 16),
39363 => conv_std_logic_vector(29835, 16),
39364 => conv_std_logic_vector(29988, 16),
39365 => conv_std_logic_vector(30141, 16),
39366 => conv_std_logic_vector(30294, 16),
39367 => conv_std_logic_vector(30447, 16),
39368 => conv_std_logic_vector(30600, 16),
39369 => conv_std_logic_vector(30753, 16),
39370 => conv_std_logic_vector(30906, 16),
39371 => conv_std_logic_vector(31059, 16),
39372 => conv_std_logic_vector(31212, 16),
39373 => conv_std_logic_vector(31365, 16),
39374 => conv_std_logic_vector(31518, 16),
39375 => conv_std_logic_vector(31671, 16),
39376 => conv_std_logic_vector(31824, 16),
39377 => conv_std_logic_vector(31977, 16),
39378 => conv_std_logic_vector(32130, 16),
39379 => conv_std_logic_vector(32283, 16),
39380 => conv_std_logic_vector(32436, 16),
39381 => conv_std_logic_vector(32589, 16),
39382 => conv_std_logic_vector(32742, 16),
39383 => conv_std_logic_vector(32895, 16),
39384 => conv_std_logic_vector(33048, 16),
39385 => conv_std_logic_vector(33201, 16),
39386 => conv_std_logic_vector(33354, 16),
39387 => conv_std_logic_vector(33507, 16),
39388 => conv_std_logic_vector(33660, 16),
39389 => conv_std_logic_vector(33813, 16),
39390 => conv_std_logic_vector(33966, 16),
39391 => conv_std_logic_vector(34119, 16),
39392 => conv_std_logic_vector(34272, 16),
39393 => conv_std_logic_vector(34425, 16),
39394 => conv_std_logic_vector(34578, 16),
39395 => conv_std_logic_vector(34731, 16),
39396 => conv_std_logic_vector(34884, 16),
39397 => conv_std_logic_vector(35037, 16),
39398 => conv_std_logic_vector(35190, 16),
39399 => conv_std_logic_vector(35343, 16),
39400 => conv_std_logic_vector(35496, 16),
39401 => conv_std_logic_vector(35649, 16),
39402 => conv_std_logic_vector(35802, 16),
39403 => conv_std_logic_vector(35955, 16),
39404 => conv_std_logic_vector(36108, 16),
39405 => conv_std_logic_vector(36261, 16),
39406 => conv_std_logic_vector(36414, 16),
39407 => conv_std_logic_vector(36567, 16),
39408 => conv_std_logic_vector(36720, 16),
39409 => conv_std_logic_vector(36873, 16),
39410 => conv_std_logic_vector(37026, 16),
39411 => conv_std_logic_vector(37179, 16),
39412 => conv_std_logic_vector(37332, 16),
39413 => conv_std_logic_vector(37485, 16),
39414 => conv_std_logic_vector(37638, 16),
39415 => conv_std_logic_vector(37791, 16),
39416 => conv_std_logic_vector(37944, 16),
39417 => conv_std_logic_vector(38097, 16),
39418 => conv_std_logic_vector(38250, 16),
39419 => conv_std_logic_vector(38403, 16),
39420 => conv_std_logic_vector(38556, 16),
39421 => conv_std_logic_vector(38709, 16),
39422 => conv_std_logic_vector(38862, 16),
39423 => conv_std_logic_vector(39015, 16),
39424 => conv_std_logic_vector(0, 16),
39425 => conv_std_logic_vector(154, 16),
39426 => conv_std_logic_vector(308, 16),
39427 => conv_std_logic_vector(462, 16),
39428 => conv_std_logic_vector(616, 16),
39429 => conv_std_logic_vector(770, 16),
39430 => conv_std_logic_vector(924, 16),
39431 => conv_std_logic_vector(1078, 16),
39432 => conv_std_logic_vector(1232, 16),
39433 => conv_std_logic_vector(1386, 16),
39434 => conv_std_logic_vector(1540, 16),
39435 => conv_std_logic_vector(1694, 16),
39436 => conv_std_logic_vector(1848, 16),
39437 => conv_std_logic_vector(2002, 16),
39438 => conv_std_logic_vector(2156, 16),
39439 => conv_std_logic_vector(2310, 16),
39440 => conv_std_logic_vector(2464, 16),
39441 => conv_std_logic_vector(2618, 16),
39442 => conv_std_logic_vector(2772, 16),
39443 => conv_std_logic_vector(2926, 16),
39444 => conv_std_logic_vector(3080, 16),
39445 => conv_std_logic_vector(3234, 16),
39446 => conv_std_logic_vector(3388, 16),
39447 => conv_std_logic_vector(3542, 16),
39448 => conv_std_logic_vector(3696, 16),
39449 => conv_std_logic_vector(3850, 16),
39450 => conv_std_logic_vector(4004, 16),
39451 => conv_std_logic_vector(4158, 16),
39452 => conv_std_logic_vector(4312, 16),
39453 => conv_std_logic_vector(4466, 16),
39454 => conv_std_logic_vector(4620, 16),
39455 => conv_std_logic_vector(4774, 16),
39456 => conv_std_logic_vector(4928, 16),
39457 => conv_std_logic_vector(5082, 16),
39458 => conv_std_logic_vector(5236, 16),
39459 => conv_std_logic_vector(5390, 16),
39460 => conv_std_logic_vector(5544, 16),
39461 => conv_std_logic_vector(5698, 16),
39462 => conv_std_logic_vector(5852, 16),
39463 => conv_std_logic_vector(6006, 16),
39464 => conv_std_logic_vector(6160, 16),
39465 => conv_std_logic_vector(6314, 16),
39466 => conv_std_logic_vector(6468, 16),
39467 => conv_std_logic_vector(6622, 16),
39468 => conv_std_logic_vector(6776, 16),
39469 => conv_std_logic_vector(6930, 16),
39470 => conv_std_logic_vector(7084, 16),
39471 => conv_std_logic_vector(7238, 16),
39472 => conv_std_logic_vector(7392, 16),
39473 => conv_std_logic_vector(7546, 16),
39474 => conv_std_logic_vector(7700, 16),
39475 => conv_std_logic_vector(7854, 16),
39476 => conv_std_logic_vector(8008, 16),
39477 => conv_std_logic_vector(8162, 16),
39478 => conv_std_logic_vector(8316, 16),
39479 => conv_std_logic_vector(8470, 16),
39480 => conv_std_logic_vector(8624, 16),
39481 => conv_std_logic_vector(8778, 16),
39482 => conv_std_logic_vector(8932, 16),
39483 => conv_std_logic_vector(9086, 16),
39484 => conv_std_logic_vector(9240, 16),
39485 => conv_std_logic_vector(9394, 16),
39486 => conv_std_logic_vector(9548, 16),
39487 => conv_std_logic_vector(9702, 16),
39488 => conv_std_logic_vector(9856, 16),
39489 => conv_std_logic_vector(10010, 16),
39490 => conv_std_logic_vector(10164, 16),
39491 => conv_std_logic_vector(10318, 16),
39492 => conv_std_logic_vector(10472, 16),
39493 => conv_std_logic_vector(10626, 16),
39494 => conv_std_logic_vector(10780, 16),
39495 => conv_std_logic_vector(10934, 16),
39496 => conv_std_logic_vector(11088, 16),
39497 => conv_std_logic_vector(11242, 16),
39498 => conv_std_logic_vector(11396, 16),
39499 => conv_std_logic_vector(11550, 16),
39500 => conv_std_logic_vector(11704, 16),
39501 => conv_std_logic_vector(11858, 16),
39502 => conv_std_logic_vector(12012, 16),
39503 => conv_std_logic_vector(12166, 16),
39504 => conv_std_logic_vector(12320, 16),
39505 => conv_std_logic_vector(12474, 16),
39506 => conv_std_logic_vector(12628, 16),
39507 => conv_std_logic_vector(12782, 16),
39508 => conv_std_logic_vector(12936, 16),
39509 => conv_std_logic_vector(13090, 16),
39510 => conv_std_logic_vector(13244, 16),
39511 => conv_std_logic_vector(13398, 16),
39512 => conv_std_logic_vector(13552, 16),
39513 => conv_std_logic_vector(13706, 16),
39514 => conv_std_logic_vector(13860, 16),
39515 => conv_std_logic_vector(14014, 16),
39516 => conv_std_logic_vector(14168, 16),
39517 => conv_std_logic_vector(14322, 16),
39518 => conv_std_logic_vector(14476, 16),
39519 => conv_std_logic_vector(14630, 16),
39520 => conv_std_logic_vector(14784, 16),
39521 => conv_std_logic_vector(14938, 16),
39522 => conv_std_logic_vector(15092, 16),
39523 => conv_std_logic_vector(15246, 16),
39524 => conv_std_logic_vector(15400, 16),
39525 => conv_std_logic_vector(15554, 16),
39526 => conv_std_logic_vector(15708, 16),
39527 => conv_std_logic_vector(15862, 16),
39528 => conv_std_logic_vector(16016, 16),
39529 => conv_std_logic_vector(16170, 16),
39530 => conv_std_logic_vector(16324, 16),
39531 => conv_std_logic_vector(16478, 16),
39532 => conv_std_logic_vector(16632, 16),
39533 => conv_std_logic_vector(16786, 16),
39534 => conv_std_logic_vector(16940, 16),
39535 => conv_std_logic_vector(17094, 16),
39536 => conv_std_logic_vector(17248, 16),
39537 => conv_std_logic_vector(17402, 16),
39538 => conv_std_logic_vector(17556, 16),
39539 => conv_std_logic_vector(17710, 16),
39540 => conv_std_logic_vector(17864, 16),
39541 => conv_std_logic_vector(18018, 16),
39542 => conv_std_logic_vector(18172, 16),
39543 => conv_std_logic_vector(18326, 16),
39544 => conv_std_logic_vector(18480, 16),
39545 => conv_std_logic_vector(18634, 16),
39546 => conv_std_logic_vector(18788, 16),
39547 => conv_std_logic_vector(18942, 16),
39548 => conv_std_logic_vector(19096, 16),
39549 => conv_std_logic_vector(19250, 16),
39550 => conv_std_logic_vector(19404, 16),
39551 => conv_std_logic_vector(19558, 16),
39552 => conv_std_logic_vector(19712, 16),
39553 => conv_std_logic_vector(19866, 16),
39554 => conv_std_logic_vector(20020, 16),
39555 => conv_std_logic_vector(20174, 16),
39556 => conv_std_logic_vector(20328, 16),
39557 => conv_std_logic_vector(20482, 16),
39558 => conv_std_logic_vector(20636, 16),
39559 => conv_std_logic_vector(20790, 16),
39560 => conv_std_logic_vector(20944, 16),
39561 => conv_std_logic_vector(21098, 16),
39562 => conv_std_logic_vector(21252, 16),
39563 => conv_std_logic_vector(21406, 16),
39564 => conv_std_logic_vector(21560, 16),
39565 => conv_std_logic_vector(21714, 16),
39566 => conv_std_logic_vector(21868, 16),
39567 => conv_std_logic_vector(22022, 16),
39568 => conv_std_logic_vector(22176, 16),
39569 => conv_std_logic_vector(22330, 16),
39570 => conv_std_logic_vector(22484, 16),
39571 => conv_std_logic_vector(22638, 16),
39572 => conv_std_logic_vector(22792, 16),
39573 => conv_std_logic_vector(22946, 16),
39574 => conv_std_logic_vector(23100, 16),
39575 => conv_std_logic_vector(23254, 16),
39576 => conv_std_logic_vector(23408, 16),
39577 => conv_std_logic_vector(23562, 16),
39578 => conv_std_logic_vector(23716, 16),
39579 => conv_std_logic_vector(23870, 16),
39580 => conv_std_logic_vector(24024, 16),
39581 => conv_std_logic_vector(24178, 16),
39582 => conv_std_logic_vector(24332, 16),
39583 => conv_std_logic_vector(24486, 16),
39584 => conv_std_logic_vector(24640, 16),
39585 => conv_std_logic_vector(24794, 16),
39586 => conv_std_logic_vector(24948, 16),
39587 => conv_std_logic_vector(25102, 16),
39588 => conv_std_logic_vector(25256, 16),
39589 => conv_std_logic_vector(25410, 16),
39590 => conv_std_logic_vector(25564, 16),
39591 => conv_std_logic_vector(25718, 16),
39592 => conv_std_logic_vector(25872, 16),
39593 => conv_std_logic_vector(26026, 16),
39594 => conv_std_logic_vector(26180, 16),
39595 => conv_std_logic_vector(26334, 16),
39596 => conv_std_logic_vector(26488, 16),
39597 => conv_std_logic_vector(26642, 16),
39598 => conv_std_logic_vector(26796, 16),
39599 => conv_std_logic_vector(26950, 16),
39600 => conv_std_logic_vector(27104, 16),
39601 => conv_std_logic_vector(27258, 16),
39602 => conv_std_logic_vector(27412, 16),
39603 => conv_std_logic_vector(27566, 16),
39604 => conv_std_logic_vector(27720, 16),
39605 => conv_std_logic_vector(27874, 16),
39606 => conv_std_logic_vector(28028, 16),
39607 => conv_std_logic_vector(28182, 16),
39608 => conv_std_logic_vector(28336, 16),
39609 => conv_std_logic_vector(28490, 16),
39610 => conv_std_logic_vector(28644, 16),
39611 => conv_std_logic_vector(28798, 16),
39612 => conv_std_logic_vector(28952, 16),
39613 => conv_std_logic_vector(29106, 16),
39614 => conv_std_logic_vector(29260, 16),
39615 => conv_std_logic_vector(29414, 16),
39616 => conv_std_logic_vector(29568, 16),
39617 => conv_std_logic_vector(29722, 16),
39618 => conv_std_logic_vector(29876, 16),
39619 => conv_std_logic_vector(30030, 16),
39620 => conv_std_logic_vector(30184, 16),
39621 => conv_std_logic_vector(30338, 16),
39622 => conv_std_logic_vector(30492, 16),
39623 => conv_std_logic_vector(30646, 16),
39624 => conv_std_logic_vector(30800, 16),
39625 => conv_std_logic_vector(30954, 16),
39626 => conv_std_logic_vector(31108, 16),
39627 => conv_std_logic_vector(31262, 16),
39628 => conv_std_logic_vector(31416, 16),
39629 => conv_std_logic_vector(31570, 16),
39630 => conv_std_logic_vector(31724, 16),
39631 => conv_std_logic_vector(31878, 16),
39632 => conv_std_logic_vector(32032, 16),
39633 => conv_std_logic_vector(32186, 16),
39634 => conv_std_logic_vector(32340, 16),
39635 => conv_std_logic_vector(32494, 16),
39636 => conv_std_logic_vector(32648, 16),
39637 => conv_std_logic_vector(32802, 16),
39638 => conv_std_logic_vector(32956, 16),
39639 => conv_std_logic_vector(33110, 16),
39640 => conv_std_logic_vector(33264, 16),
39641 => conv_std_logic_vector(33418, 16),
39642 => conv_std_logic_vector(33572, 16),
39643 => conv_std_logic_vector(33726, 16),
39644 => conv_std_logic_vector(33880, 16),
39645 => conv_std_logic_vector(34034, 16),
39646 => conv_std_logic_vector(34188, 16),
39647 => conv_std_logic_vector(34342, 16),
39648 => conv_std_logic_vector(34496, 16),
39649 => conv_std_logic_vector(34650, 16),
39650 => conv_std_logic_vector(34804, 16),
39651 => conv_std_logic_vector(34958, 16),
39652 => conv_std_logic_vector(35112, 16),
39653 => conv_std_logic_vector(35266, 16),
39654 => conv_std_logic_vector(35420, 16),
39655 => conv_std_logic_vector(35574, 16),
39656 => conv_std_logic_vector(35728, 16),
39657 => conv_std_logic_vector(35882, 16),
39658 => conv_std_logic_vector(36036, 16),
39659 => conv_std_logic_vector(36190, 16),
39660 => conv_std_logic_vector(36344, 16),
39661 => conv_std_logic_vector(36498, 16),
39662 => conv_std_logic_vector(36652, 16),
39663 => conv_std_logic_vector(36806, 16),
39664 => conv_std_logic_vector(36960, 16),
39665 => conv_std_logic_vector(37114, 16),
39666 => conv_std_logic_vector(37268, 16),
39667 => conv_std_logic_vector(37422, 16),
39668 => conv_std_logic_vector(37576, 16),
39669 => conv_std_logic_vector(37730, 16),
39670 => conv_std_logic_vector(37884, 16),
39671 => conv_std_logic_vector(38038, 16),
39672 => conv_std_logic_vector(38192, 16),
39673 => conv_std_logic_vector(38346, 16),
39674 => conv_std_logic_vector(38500, 16),
39675 => conv_std_logic_vector(38654, 16),
39676 => conv_std_logic_vector(38808, 16),
39677 => conv_std_logic_vector(38962, 16),
39678 => conv_std_logic_vector(39116, 16),
39679 => conv_std_logic_vector(39270, 16),
39680 => conv_std_logic_vector(0, 16),
39681 => conv_std_logic_vector(155, 16),
39682 => conv_std_logic_vector(310, 16),
39683 => conv_std_logic_vector(465, 16),
39684 => conv_std_logic_vector(620, 16),
39685 => conv_std_logic_vector(775, 16),
39686 => conv_std_logic_vector(930, 16),
39687 => conv_std_logic_vector(1085, 16),
39688 => conv_std_logic_vector(1240, 16),
39689 => conv_std_logic_vector(1395, 16),
39690 => conv_std_logic_vector(1550, 16),
39691 => conv_std_logic_vector(1705, 16),
39692 => conv_std_logic_vector(1860, 16),
39693 => conv_std_logic_vector(2015, 16),
39694 => conv_std_logic_vector(2170, 16),
39695 => conv_std_logic_vector(2325, 16),
39696 => conv_std_logic_vector(2480, 16),
39697 => conv_std_logic_vector(2635, 16),
39698 => conv_std_logic_vector(2790, 16),
39699 => conv_std_logic_vector(2945, 16),
39700 => conv_std_logic_vector(3100, 16),
39701 => conv_std_logic_vector(3255, 16),
39702 => conv_std_logic_vector(3410, 16),
39703 => conv_std_logic_vector(3565, 16),
39704 => conv_std_logic_vector(3720, 16),
39705 => conv_std_logic_vector(3875, 16),
39706 => conv_std_logic_vector(4030, 16),
39707 => conv_std_logic_vector(4185, 16),
39708 => conv_std_logic_vector(4340, 16),
39709 => conv_std_logic_vector(4495, 16),
39710 => conv_std_logic_vector(4650, 16),
39711 => conv_std_logic_vector(4805, 16),
39712 => conv_std_logic_vector(4960, 16),
39713 => conv_std_logic_vector(5115, 16),
39714 => conv_std_logic_vector(5270, 16),
39715 => conv_std_logic_vector(5425, 16),
39716 => conv_std_logic_vector(5580, 16),
39717 => conv_std_logic_vector(5735, 16),
39718 => conv_std_logic_vector(5890, 16),
39719 => conv_std_logic_vector(6045, 16),
39720 => conv_std_logic_vector(6200, 16),
39721 => conv_std_logic_vector(6355, 16),
39722 => conv_std_logic_vector(6510, 16),
39723 => conv_std_logic_vector(6665, 16),
39724 => conv_std_logic_vector(6820, 16),
39725 => conv_std_logic_vector(6975, 16),
39726 => conv_std_logic_vector(7130, 16),
39727 => conv_std_logic_vector(7285, 16),
39728 => conv_std_logic_vector(7440, 16),
39729 => conv_std_logic_vector(7595, 16),
39730 => conv_std_logic_vector(7750, 16),
39731 => conv_std_logic_vector(7905, 16),
39732 => conv_std_logic_vector(8060, 16),
39733 => conv_std_logic_vector(8215, 16),
39734 => conv_std_logic_vector(8370, 16),
39735 => conv_std_logic_vector(8525, 16),
39736 => conv_std_logic_vector(8680, 16),
39737 => conv_std_logic_vector(8835, 16),
39738 => conv_std_logic_vector(8990, 16),
39739 => conv_std_logic_vector(9145, 16),
39740 => conv_std_logic_vector(9300, 16),
39741 => conv_std_logic_vector(9455, 16),
39742 => conv_std_logic_vector(9610, 16),
39743 => conv_std_logic_vector(9765, 16),
39744 => conv_std_logic_vector(9920, 16),
39745 => conv_std_logic_vector(10075, 16),
39746 => conv_std_logic_vector(10230, 16),
39747 => conv_std_logic_vector(10385, 16),
39748 => conv_std_logic_vector(10540, 16),
39749 => conv_std_logic_vector(10695, 16),
39750 => conv_std_logic_vector(10850, 16),
39751 => conv_std_logic_vector(11005, 16),
39752 => conv_std_logic_vector(11160, 16),
39753 => conv_std_logic_vector(11315, 16),
39754 => conv_std_logic_vector(11470, 16),
39755 => conv_std_logic_vector(11625, 16),
39756 => conv_std_logic_vector(11780, 16),
39757 => conv_std_logic_vector(11935, 16),
39758 => conv_std_logic_vector(12090, 16),
39759 => conv_std_logic_vector(12245, 16),
39760 => conv_std_logic_vector(12400, 16),
39761 => conv_std_logic_vector(12555, 16),
39762 => conv_std_logic_vector(12710, 16),
39763 => conv_std_logic_vector(12865, 16),
39764 => conv_std_logic_vector(13020, 16),
39765 => conv_std_logic_vector(13175, 16),
39766 => conv_std_logic_vector(13330, 16),
39767 => conv_std_logic_vector(13485, 16),
39768 => conv_std_logic_vector(13640, 16),
39769 => conv_std_logic_vector(13795, 16),
39770 => conv_std_logic_vector(13950, 16),
39771 => conv_std_logic_vector(14105, 16),
39772 => conv_std_logic_vector(14260, 16),
39773 => conv_std_logic_vector(14415, 16),
39774 => conv_std_logic_vector(14570, 16),
39775 => conv_std_logic_vector(14725, 16),
39776 => conv_std_logic_vector(14880, 16),
39777 => conv_std_logic_vector(15035, 16),
39778 => conv_std_logic_vector(15190, 16),
39779 => conv_std_logic_vector(15345, 16),
39780 => conv_std_logic_vector(15500, 16),
39781 => conv_std_logic_vector(15655, 16),
39782 => conv_std_logic_vector(15810, 16),
39783 => conv_std_logic_vector(15965, 16),
39784 => conv_std_logic_vector(16120, 16),
39785 => conv_std_logic_vector(16275, 16),
39786 => conv_std_logic_vector(16430, 16),
39787 => conv_std_logic_vector(16585, 16),
39788 => conv_std_logic_vector(16740, 16),
39789 => conv_std_logic_vector(16895, 16),
39790 => conv_std_logic_vector(17050, 16),
39791 => conv_std_logic_vector(17205, 16),
39792 => conv_std_logic_vector(17360, 16),
39793 => conv_std_logic_vector(17515, 16),
39794 => conv_std_logic_vector(17670, 16),
39795 => conv_std_logic_vector(17825, 16),
39796 => conv_std_logic_vector(17980, 16),
39797 => conv_std_logic_vector(18135, 16),
39798 => conv_std_logic_vector(18290, 16),
39799 => conv_std_logic_vector(18445, 16),
39800 => conv_std_logic_vector(18600, 16),
39801 => conv_std_logic_vector(18755, 16),
39802 => conv_std_logic_vector(18910, 16),
39803 => conv_std_logic_vector(19065, 16),
39804 => conv_std_logic_vector(19220, 16),
39805 => conv_std_logic_vector(19375, 16),
39806 => conv_std_logic_vector(19530, 16),
39807 => conv_std_logic_vector(19685, 16),
39808 => conv_std_logic_vector(19840, 16),
39809 => conv_std_logic_vector(19995, 16),
39810 => conv_std_logic_vector(20150, 16),
39811 => conv_std_logic_vector(20305, 16),
39812 => conv_std_logic_vector(20460, 16),
39813 => conv_std_logic_vector(20615, 16),
39814 => conv_std_logic_vector(20770, 16),
39815 => conv_std_logic_vector(20925, 16),
39816 => conv_std_logic_vector(21080, 16),
39817 => conv_std_logic_vector(21235, 16),
39818 => conv_std_logic_vector(21390, 16),
39819 => conv_std_logic_vector(21545, 16),
39820 => conv_std_logic_vector(21700, 16),
39821 => conv_std_logic_vector(21855, 16),
39822 => conv_std_logic_vector(22010, 16),
39823 => conv_std_logic_vector(22165, 16),
39824 => conv_std_logic_vector(22320, 16),
39825 => conv_std_logic_vector(22475, 16),
39826 => conv_std_logic_vector(22630, 16),
39827 => conv_std_logic_vector(22785, 16),
39828 => conv_std_logic_vector(22940, 16),
39829 => conv_std_logic_vector(23095, 16),
39830 => conv_std_logic_vector(23250, 16),
39831 => conv_std_logic_vector(23405, 16),
39832 => conv_std_logic_vector(23560, 16),
39833 => conv_std_logic_vector(23715, 16),
39834 => conv_std_logic_vector(23870, 16),
39835 => conv_std_logic_vector(24025, 16),
39836 => conv_std_logic_vector(24180, 16),
39837 => conv_std_logic_vector(24335, 16),
39838 => conv_std_logic_vector(24490, 16),
39839 => conv_std_logic_vector(24645, 16),
39840 => conv_std_logic_vector(24800, 16),
39841 => conv_std_logic_vector(24955, 16),
39842 => conv_std_logic_vector(25110, 16),
39843 => conv_std_logic_vector(25265, 16),
39844 => conv_std_logic_vector(25420, 16),
39845 => conv_std_logic_vector(25575, 16),
39846 => conv_std_logic_vector(25730, 16),
39847 => conv_std_logic_vector(25885, 16),
39848 => conv_std_logic_vector(26040, 16),
39849 => conv_std_logic_vector(26195, 16),
39850 => conv_std_logic_vector(26350, 16),
39851 => conv_std_logic_vector(26505, 16),
39852 => conv_std_logic_vector(26660, 16),
39853 => conv_std_logic_vector(26815, 16),
39854 => conv_std_logic_vector(26970, 16),
39855 => conv_std_logic_vector(27125, 16),
39856 => conv_std_logic_vector(27280, 16),
39857 => conv_std_logic_vector(27435, 16),
39858 => conv_std_logic_vector(27590, 16),
39859 => conv_std_logic_vector(27745, 16),
39860 => conv_std_logic_vector(27900, 16),
39861 => conv_std_logic_vector(28055, 16),
39862 => conv_std_logic_vector(28210, 16),
39863 => conv_std_logic_vector(28365, 16),
39864 => conv_std_logic_vector(28520, 16),
39865 => conv_std_logic_vector(28675, 16),
39866 => conv_std_logic_vector(28830, 16),
39867 => conv_std_logic_vector(28985, 16),
39868 => conv_std_logic_vector(29140, 16),
39869 => conv_std_logic_vector(29295, 16),
39870 => conv_std_logic_vector(29450, 16),
39871 => conv_std_logic_vector(29605, 16),
39872 => conv_std_logic_vector(29760, 16),
39873 => conv_std_logic_vector(29915, 16),
39874 => conv_std_logic_vector(30070, 16),
39875 => conv_std_logic_vector(30225, 16),
39876 => conv_std_logic_vector(30380, 16),
39877 => conv_std_logic_vector(30535, 16),
39878 => conv_std_logic_vector(30690, 16),
39879 => conv_std_logic_vector(30845, 16),
39880 => conv_std_logic_vector(31000, 16),
39881 => conv_std_logic_vector(31155, 16),
39882 => conv_std_logic_vector(31310, 16),
39883 => conv_std_logic_vector(31465, 16),
39884 => conv_std_logic_vector(31620, 16),
39885 => conv_std_logic_vector(31775, 16),
39886 => conv_std_logic_vector(31930, 16),
39887 => conv_std_logic_vector(32085, 16),
39888 => conv_std_logic_vector(32240, 16),
39889 => conv_std_logic_vector(32395, 16),
39890 => conv_std_logic_vector(32550, 16),
39891 => conv_std_logic_vector(32705, 16),
39892 => conv_std_logic_vector(32860, 16),
39893 => conv_std_logic_vector(33015, 16),
39894 => conv_std_logic_vector(33170, 16),
39895 => conv_std_logic_vector(33325, 16),
39896 => conv_std_logic_vector(33480, 16),
39897 => conv_std_logic_vector(33635, 16),
39898 => conv_std_logic_vector(33790, 16),
39899 => conv_std_logic_vector(33945, 16),
39900 => conv_std_logic_vector(34100, 16),
39901 => conv_std_logic_vector(34255, 16),
39902 => conv_std_logic_vector(34410, 16),
39903 => conv_std_logic_vector(34565, 16),
39904 => conv_std_logic_vector(34720, 16),
39905 => conv_std_logic_vector(34875, 16),
39906 => conv_std_logic_vector(35030, 16),
39907 => conv_std_logic_vector(35185, 16),
39908 => conv_std_logic_vector(35340, 16),
39909 => conv_std_logic_vector(35495, 16),
39910 => conv_std_logic_vector(35650, 16),
39911 => conv_std_logic_vector(35805, 16),
39912 => conv_std_logic_vector(35960, 16),
39913 => conv_std_logic_vector(36115, 16),
39914 => conv_std_logic_vector(36270, 16),
39915 => conv_std_logic_vector(36425, 16),
39916 => conv_std_logic_vector(36580, 16),
39917 => conv_std_logic_vector(36735, 16),
39918 => conv_std_logic_vector(36890, 16),
39919 => conv_std_logic_vector(37045, 16),
39920 => conv_std_logic_vector(37200, 16),
39921 => conv_std_logic_vector(37355, 16),
39922 => conv_std_logic_vector(37510, 16),
39923 => conv_std_logic_vector(37665, 16),
39924 => conv_std_logic_vector(37820, 16),
39925 => conv_std_logic_vector(37975, 16),
39926 => conv_std_logic_vector(38130, 16),
39927 => conv_std_logic_vector(38285, 16),
39928 => conv_std_logic_vector(38440, 16),
39929 => conv_std_logic_vector(38595, 16),
39930 => conv_std_logic_vector(38750, 16),
39931 => conv_std_logic_vector(38905, 16),
39932 => conv_std_logic_vector(39060, 16),
39933 => conv_std_logic_vector(39215, 16),
39934 => conv_std_logic_vector(39370, 16),
39935 => conv_std_logic_vector(39525, 16),
39936 => conv_std_logic_vector(0, 16),
39937 => conv_std_logic_vector(156, 16),
39938 => conv_std_logic_vector(312, 16),
39939 => conv_std_logic_vector(468, 16),
39940 => conv_std_logic_vector(624, 16),
39941 => conv_std_logic_vector(780, 16),
39942 => conv_std_logic_vector(936, 16),
39943 => conv_std_logic_vector(1092, 16),
39944 => conv_std_logic_vector(1248, 16),
39945 => conv_std_logic_vector(1404, 16),
39946 => conv_std_logic_vector(1560, 16),
39947 => conv_std_logic_vector(1716, 16),
39948 => conv_std_logic_vector(1872, 16),
39949 => conv_std_logic_vector(2028, 16),
39950 => conv_std_logic_vector(2184, 16),
39951 => conv_std_logic_vector(2340, 16),
39952 => conv_std_logic_vector(2496, 16),
39953 => conv_std_logic_vector(2652, 16),
39954 => conv_std_logic_vector(2808, 16),
39955 => conv_std_logic_vector(2964, 16),
39956 => conv_std_logic_vector(3120, 16),
39957 => conv_std_logic_vector(3276, 16),
39958 => conv_std_logic_vector(3432, 16),
39959 => conv_std_logic_vector(3588, 16),
39960 => conv_std_logic_vector(3744, 16),
39961 => conv_std_logic_vector(3900, 16),
39962 => conv_std_logic_vector(4056, 16),
39963 => conv_std_logic_vector(4212, 16),
39964 => conv_std_logic_vector(4368, 16),
39965 => conv_std_logic_vector(4524, 16),
39966 => conv_std_logic_vector(4680, 16),
39967 => conv_std_logic_vector(4836, 16),
39968 => conv_std_logic_vector(4992, 16),
39969 => conv_std_logic_vector(5148, 16),
39970 => conv_std_logic_vector(5304, 16),
39971 => conv_std_logic_vector(5460, 16),
39972 => conv_std_logic_vector(5616, 16),
39973 => conv_std_logic_vector(5772, 16),
39974 => conv_std_logic_vector(5928, 16),
39975 => conv_std_logic_vector(6084, 16),
39976 => conv_std_logic_vector(6240, 16),
39977 => conv_std_logic_vector(6396, 16),
39978 => conv_std_logic_vector(6552, 16),
39979 => conv_std_logic_vector(6708, 16),
39980 => conv_std_logic_vector(6864, 16),
39981 => conv_std_logic_vector(7020, 16),
39982 => conv_std_logic_vector(7176, 16),
39983 => conv_std_logic_vector(7332, 16),
39984 => conv_std_logic_vector(7488, 16),
39985 => conv_std_logic_vector(7644, 16),
39986 => conv_std_logic_vector(7800, 16),
39987 => conv_std_logic_vector(7956, 16),
39988 => conv_std_logic_vector(8112, 16),
39989 => conv_std_logic_vector(8268, 16),
39990 => conv_std_logic_vector(8424, 16),
39991 => conv_std_logic_vector(8580, 16),
39992 => conv_std_logic_vector(8736, 16),
39993 => conv_std_logic_vector(8892, 16),
39994 => conv_std_logic_vector(9048, 16),
39995 => conv_std_logic_vector(9204, 16),
39996 => conv_std_logic_vector(9360, 16),
39997 => conv_std_logic_vector(9516, 16),
39998 => conv_std_logic_vector(9672, 16),
39999 => conv_std_logic_vector(9828, 16),
40000 => conv_std_logic_vector(9984, 16),
40001 => conv_std_logic_vector(10140, 16),
40002 => conv_std_logic_vector(10296, 16),
40003 => conv_std_logic_vector(10452, 16),
40004 => conv_std_logic_vector(10608, 16),
40005 => conv_std_logic_vector(10764, 16),
40006 => conv_std_logic_vector(10920, 16),
40007 => conv_std_logic_vector(11076, 16),
40008 => conv_std_logic_vector(11232, 16),
40009 => conv_std_logic_vector(11388, 16),
40010 => conv_std_logic_vector(11544, 16),
40011 => conv_std_logic_vector(11700, 16),
40012 => conv_std_logic_vector(11856, 16),
40013 => conv_std_logic_vector(12012, 16),
40014 => conv_std_logic_vector(12168, 16),
40015 => conv_std_logic_vector(12324, 16),
40016 => conv_std_logic_vector(12480, 16),
40017 => conv_std_logic_vector(12636, 16),
40018 => conv_std_logic_vector(12792, 16),
40019 => conv_std_logic_vector(12948, 16),
40020 => conv_std_logic_vector(13104, 16),
40021 => conv_std_logic_vector(13260, 16),
40022 => conv_std_logic_vector(13416, 16),
40023 => conv_std_logic_vector(13572, 16),
40024 => conv_std_logic_vector(13728, 16),
40025 => conv_std_logic_vector(13884, 16),
40026 => conv_std_logic_vector(14040, 16),
40027 => conv_std_logic_vector(14196, 16),
40028 => conv_std_logic_vector(14352, 16),
40029 => conv_std_logic_vector(14508, 16),
40030 => conv_std_logic_vector(14664, 16),
40031 => conv_std_logic_vector(14820, 16),
40032 => conv_std_logic_vector(14976, 16),
40033 => conv_std_logic_vector(15132, 16),
40034 => conv_std_logic_vector(15288, 16),
40035 => conv_std_logic_vector(15444, 16),
40036 => conv_std_logic_vector(15600, 16),
40037 => conv_std_logic_vector(15756, 16),
40038 => conv_std_logic_vector(15912, 16),
40039 => conv_std_logic_vector(16068, 16),
40040 => conv_std_logic_vector(16224, 16),
40041 => conv_std_logic_vector(16380, 16),
40042 => conv_std_logic_vector(16536, 16),
40043 => conv_std_logic_vector(16692, 16),
40044 => conv_std_logic_vector(16848, 16),
40045 => conv_std_logic_vector(17004, 16),
40046 => conv_std_logic_vector(17160, 16),
40047 => conv_std_logic_vector(17316, 16),
40048 => conv_std_logic_vector(17472, 16),
40049 => conv_std_logic_vector(17628, 16),
40050 => conv_std_logic_vector(17784, 16),
40051 => conv_std_logic_vector(17940, 16),
40052 => conv_std_logic_vector(18096, 16),
40053 => conv_std_logic_vector(18252, 16),
40054 => conv_std_logic_vector(18408, 16),
40055 => conv_std_logic_vector(18564, 16),
40056 => conv_std_logic_vector(18720, 16),
40057 => conv_std_logic_vector(18876, 16),
40058 => conv_std_logic_vector(19032, 16),
40059 => conv_std_logic_vector(19188, 16),
40060 => conv_std_logic_vector(19344, 16),
40061 => conv_std_logic_vector(19500, 16),
40062 => conv_std_logic_vector(19656, 16),
40063 => conv_std_logic_vector(19812, 16),
40064 => conv_std_logic_vector(19968, 16),
40065 => conv_std_logic_vector(20124, 16),
40066 => conv_std_logic_vector(20280, 16),
40067 => conv_std_logic_vector(20436, 16),
40068 => conv_std_logic_vector(20592, 16),
40069 => conv_std_logic_vector(20748, 16),
40070 => conv_std_logic_vector(20904, 16),
40071 => conv_std_logic_vector(21060, 16),
40072 => conv_std_logic_vector(21216, 16),
40073 => conv_std_logic_vector(21372, 16),
40074 => conv_std_logic_vector(21528, 16),
40075 => conv_std_logic_vector(21684, 16),
40076 => conv_std_logic_vector(21840, 16),
40077 => conv_std_logic_vector(21996, 16),
40078 => conv_std_logic_vector(22152, 16),
40079 => conv_std_logic_vector(22308, 16),
40080 => conv_std_logic_vector(22464, 16),
40081 => conv_std_logic_vector(22620, 16),
40082 => conv_std_logic_vector(22776, 16),
40083 => conv_std_logic_vector(22932, 16),
40084 => conv_std_logic_vector(23088, 16),
40085 => conv_std_logic_vector(23244, 16),
40086 => conv_std_logic_vector(23400, 16),
40087 => conv_std_logic_vector(23556, 16),
40088 => conv_std_logic_vector(23712, 16),
40089 => conv_std_logic_vector(23868, 16),
40090 => conv_std_logic_vector(24024, 16),
40091 => conv_std_logic_vector(24180, 16),
40092 => conv_std_logic_vector(24336, 16),
40093 => conv_std_logic_vector(24492, 16),
40094 => conv_std_logic_vector(24648, 16),
40095 => conv_std_logic_vector(24804, 16),
40096 => conv_std_logic_vector(24960, 16),
40097 => conv_std_logic_vector(25116, 16),
40098 => conv_std_logic_vector(25272, 16),
40099 => conv_std_logic_vector(25428, 16),
40100 => conv_std_logic_vector(25584, 16),
40101 => conv_std_logic_vector(25740, 16),
40102 => conv_std_logic_vector(25896, 16),
40103 => conv_std_logic_vector(26052, 16),
40104 => conv_std_logic_vector(26208, 16),
40105 => conv_std_logic_vector(26364, 16),
40106 => conv_std_logic_vector(26520, 16),
40107 => conv_std_logic_vector(26676, 16),
40108 => conv_std_logic_vector(26832, 16),
40109 => conv_std_logic_vector(26988, 16),
40110 => conv_std_logic_vector(27144, 16),
40111 => conv_std_logic_vector(27300, 16),
40112 => conv_std_logic_vector(27456, 16),
40113 => conv_std_logic_vector(27612, 16),
40114 => conv_std_logic_vector(27768, 16),
40115 => conv_std_logic_vector(27924, 16),
40116 => conv_std_logic_vector(28080, 16),
40117 => conv_std_logic_vector(28236, 16),
40118 => conv_std_logic_vector(28392, 16),
40119 => conv_std_logic_vector(28548, 16),
40120 => conv_std_logic_vector(28704, 16),
40121 => conv_std_logic_vector(28860, 16),
40122 => conv_std_logic_vector(29016, 16),
40123 => conv_std_logic_vector(29172, 16),
40124 => conv_std_logic_vector(29328, 16),
40125 => conv_std_logic_vector(29484, 16),
40126 => conv_std_logic_vector(29640, 16),
40127 => conv_std_logic_vector(29796, 16),
40128 => conv_std_logic_vector(29952, 16),
40129 => conv_std_logic_vector(30108, 16),
40130 => conv_std_logic_vector(30264, 16),
40131 => conv_std_logic_vector(30420, 16),
40132 => conv_std_logic_vector(30576, 16),
40133 => conv_std_logic_vector(30732, 16),
40134 => conv_std_logic_vector(30888, 16),
40135 => conv_std_logic_vector(31044, 16),
40136 => conv_std_logic_vector(31200, 16),
40137 => conv_std_logic_vector(31356, 16),
40138 => conv_std_logic_vector(31512, 16),
40139 => conv_std_logic_vector(31668, 16),
40140 => conv_std_logic_vector(31824, 16),
40141 => conv_std_logic_vector(31980, 16),
40142 => conv_std_logic_vector(32136, 16),
40143 => conv_std_logic_vector(32292, 16),
40144 => conv_std_logic_vector(32448, 16),
40145 => conv_std_logic_vector(32604, 16),
40146 => conv_std_logic_vector(32760, 16),
40147 => conv_std_logic_vector(32916, 16),
40148 => conv_std_logic_vector(33072, 16),
40149 => conv_std_logic_vector(33228, 16),
40150 => conv_std_logic_vector(33384, 16),
40151 => conv_std_logic_vector(33540, 16),
40152 => conv_std_logic_vector(33696, 16),
40153 => conv_std_logic_vector(33852, 16),
40154 => conv_std_logic_vector(34008, 16),
40155 => conv_std_logic_vector(34164, 16),
40156 => conv_std_logic_vector(34320, 16),
40157 => conv_std_logic_vector(34476, 16),
40158 => conv_std_logic_vector(34632, 16),
40159 => conv_std_logic_vector(34788, 16),
40160 => conv_std_logic_vector(34944, 16),
40161 => conv_std_logic_vector(35100, 16),
40162 => conv_std_logic_vector(35256, 16),
40163 => conv_std_logic_vector(35412, 16),
40164 => conv_std_logic_vector(35568, 16),
40165 => conv_std_logic_vector(35724, 16),
40166 => conv_std_logic_vector(35880, 16),
40167 => conv_std_logic_vector(36036, 16),
40168 => conv_std_logic_vector(36192, 16),
40169 => conv_std_logic_vector(36348, 16),
40170 => conv_std_logic_vector(36504, 16),
40171 => conv_std_logic_vector(36660, 16),
40172 => conv_std_logic_vector(36816, 16),
40173 => conv_std_logic_vector(36972, 16),
40174 => conv_std_logic_vector(37128, 16),
40175 => conv_std_logic_vector(37284, 16),
40176 => conv_std_logic_vector(37440, 16),
40177 => conv_std_logic_vector(37596, 16),
40178 => conv_std_logic_vector(37752, 16),
40179 => conv_std_logic_vector(37908, 16),
40180 => conv_std_logic_vector(38064, 16),
40181 => conv_std_logic_vector(38220, 16),
40182 => conv_std_logic_vector(38376, 16),
40183 => conv_std_logic_vector(38532, 16),
40184 => conv_std_logic_vector(38688, 16),
40185 => conv_std_logic_vector(38844, 16),
40186 => conv_std_logic_vector(39000, 16),
40187 => conv_std_logic_vector(39156, 16),
40188 => conv_std_logic_vector(39312, 16),
40189 => conv_std_logic_vector(39468, 16),
40190 => conv_std_logic_vector(39624, 16),
40191 => conv_std_logic_vector(39780, 16),
40192 => conv_std_logic_vector(0, 16),
40193 => conv_std_logic_vector(157, 16),
40194 => conv_std_logic_vector(314, 16),
40195 => conv_std_logic_vector(471, 16),
40196 => conv_std_logic_vector(628, 16),
40197 => conv_std_logic_vector(785, 16),
40198 => conv_std_logic_vector(942, 16),
40199 => conv_std_logic_vector(1099, 16),
40200 => conv_std_logic_vector(1256, 16),
40201 => conv_std_logic_vector(1413, 16),
40202 => conv_std_logic_vector(1570, 16),
40203 => conv_std_logic_vector(1727, 16),
40204 => conv_std_logic_vector(1884, 16),
40205 => conv_std_logic_vector(2041, 16),
40206 => conv_std_logic_vector(2198, 16),
40207 => conv_std_logic_vector(2355, 16),
40208 => conv_std_logic_vector(2512, 16),
40209 => conv_std_logic_vector(2669, 16),
40210 => conv_std_logic_vector(2826, 16),
40211 => conv_std_logic_vector(2983, 16),
40212 => conv_std_logic_vector(3140, 16),
40213 => conv_std_logic_vector(3297, 16),
40214 => conv_std_logic_vector(3454, 16),
40215 => conv_std_logic_vector(3611, 16),
40216 => conv_std_logic_vector(3768, 16),
40217 => conv_std_logic_vector(3925, 16),
40218 => conv_std_logic_vector(4082, 16),
40219 => conv_std_logic_vector(4239, 16),
40220 => conv_std_logic_vector(4396, 16),
40221 => conv_std_logic_vector(4553, 16),
40222 => conv_std_logic_vector(4710, 16),
40223 => conv_std_logic_vector(4867, 16),
40224 => conv_std_logic_vector(5024, 16),
40225 => conv_std_logic_vector(5181, 16),
40226 => conv_std_logic_vector(5338, 16),
40227 => conv_std_logic_vector(5495, 16),
40228 => conv_std_logic_vector(5652, 16),
40229 => conv_std_logic_vector(5809, 16),
40230 => conv_std_logic_vector(5966, 16),
40231 => conv_std_logic_vector(6123, 16),
40232 => conv_std_logic_vector(6280, 16),
40233 => conv_std_logic_vector(6437, 16),
40234 => conv_std_logic_vector(6594, 16),
40235 => conv_std_logic_vector(6751, 16),
40236 => conv_std_logic_vector(6908, 16),
40237 => conv_std_logic_vector(7065, 16),
40238 => conv_std_logic_vector(7222, 16),
40239 => conv_std_logic_vector(7379, 16),
40240 => conv_std_logic_vector(7536, 16),
40241 => conv_std_logic_vector(7693, 16),
40242 => conv_std_logic_vector(7850, 16),
40243 => conv_std_logic_vector(8007, 16),
40244 => conv_std_logic_vector(8164, 16),
40245 => conv_std_logic_vector(8321, 16),
40246 => conv_std_logic_vector(8478, 16),
40247 => conv_std_logic_vector(8635, 16),
40248 => conv_std_logic_vector(8792, 16),
40249 => conv_std_logic_vector(8949, 16),
40250 => conv_std_logic_vector(9106, 16),
40251 => conv_std_logic_vector(9263, 16),
40252 => conv_std_logic_vector(9420, 16),
40253 => conv_std_logic_vector(9577, 16),
40254 => conv_std_logic_vector(9734, 16),
40255 => conv_std_logic_vector(9891, 16),
40256 => conv_std_logic_vector(10048, 16),
40257 => conv_std_logic_vector(10205, 16),
40258 => conv_std_logic_vector(10362, 16),
40259 => conv_std_logic_vector(10519, 16),
40260 => conv_std_logic_vector(10676, 16),
40261 => conv_std_logic_vector(10833, 16),
40262 => conv_std_logic_vector(10990, 16),
40263 => conv_std_logic_vector(11147, 16),
40264 => conv_std_logic_vector(11304, 16),
40265 => conv_std_logic_vector(11461, 16),
40266 => conv_std_logic_vector(11618, 16),
40267 => conv_std_logic_vector(11775, 16),
40268 => conv_std_logic_vector(11932, 16),
40269 => conv_std_logic_vector(12089, 16),
40270 => conv_std_logic_vector(12246, 16),
40271 => conv_std_logic_vector(12403, 16),
40272 => conv_std_logic_vector(12560, 16),
40273 => conv_std_logic_vector(12717, 16),
40274 => conv_std_logic_vector(12874, 16),
40275 => conv_std_logic_vector(13031, 16),
40276 => conv_std_logic_vector(13188, 16),
40277 => conv_std_logic_vector(13345, 16),
40278 => conv_std_logic_vector(13502, 16),
40279 => conv_std_logic_vector(13659, 16),
40280 => conv_std_logic_vector(13816, 16),
40281 => conv_std_logic_vector(13973, 16),
40282 => conv_std_logic_vector(14130, 16),
40283 => conv_std_logic_vector(14287, 16),
40284 => conv_std_logic_vector(14444, 16),
40285 => conv_std_logic_vector(14601, 16),
40286 => conv_std_logic_vector(14758, 16),
40287 => conv_std_logic_vector(14915, 16),
40288 => conv_std_logic_vector(15072, 16),
40289 => conv_std_logic_vector(15229, 16),
40290 => conv_std_logic_vector(15386, 16),
40291 => conv_std_logic_vector(15543, 16),
40292 => conv_std_logic_vector(15700, 16),
40293 => conv_std_logic_vector(15857, 16),
40294 => conv_std_logic_vector(16014, 16),
40295 => conv_std_logic_vector(16171, 16),
40296 => conv_std_logic_vector(16328, 16),
40297 => conv_std_logic_vector(16485, 16),
40298 => conv_std_logic_vector(16642, 16),
40299 => conv_std_logic_vector(16799, 16),
40300 => conv_std_logic_vector(16956, 16),
40301 => conv_std_logic_vector(17113, 16),
40302 => conv_std_logic_vector(17270, 16),
40303 => conv_std_logic_vector(17427, 16),
40304 => conv_std_logic_vector(17584, 16),
40305 => conv_std_logic_vector(17741, 16),
40306 => conv_std_logic_vector(17898, 16),
40307 => conv_std_logic_vector(18055, 16),
40308 => conv_std_logic_vector(18212, 16),
40309 => conv_std_logic_vector(18369, 16),
40310 => conv_std_logic_vector(18526, 16),
40311 => conv_std_logic_vector(18683, 16),
40312 => conv_std_logic_vector(18840, 16),
40313 => conv_std_logic_vector(18997, 16),
40314 => conv_std_logic_vector(19154, 16),
40315 => conv_std_logic_vector(19311, 16),
40316 => conv_std_logic_vector(19468, 16),
40317 => conv_std_logic_vector(19625, 16),
40318 => conv_std_logic_vector(19782, 16),
40319 => conv_std_logic_vector(19939, 16),
40320 => conv_std_logic_vector(20096, 16),
40321 => conv_std_logic_vector(20253, 16),
40322 => conv_std_logic_vector(20410, 16),
40323 => conv_std_logic_vector(20567, 16),
40324 => conv_std_logic_vector(20724, 16),
40325 => conv_std_logic_vector(20881, 16),
40326 => conv_std_logic_vector(21038, 16),
40327 => conv_std_logic_vector(21195, 16),
40328 => conv_std_logic_vector(21352, 16),
40329 => conv_std_logic_vector(21509, 16),
40330 => conv_std_logic_vector(21666, 16),
40331 => conv_std_logic_vector(21823, 16),
40332 => conv_std_logic_vector(21980, 16),
40333 => conv_std_logic_vector(22137, 16),
40334 => conv_std_logic_vector(22294, 16),
40335 => conv_std_logic_vector(22451, 16),
40336 => conv_std_logic_vector(22608, 16),
40337 => conv_std_logic_vector(22765, 16),
40338 => conv_std_logic_vector(22922, 16),
40339 => conv_std_logic_vector(23079, 16),
40340 => conv_std_logic_vector(23236, 16),
40341 => conv_std_logic_vector(23393, 16),
40342 => conv_std_logic_vector(23550, 16),
40343 => conv_std_logic_vector(23707, 16),
40344 => conv_std_logic_vector(23864, 16),
40345 => conv_std_logic_vector(24021, 16),
40346 => conv_std_logic_vector(24178, 16),
40347 => conv_std_logic_vector(24335, 16),
40348 => conv_std_logic_vector(24492, 16),
40349 => conv_std_logic_vector(24649, 16),
40350 => conv_std_logic_vector(24806, 16),
40351 => conv_std_logic_vector(24963, 16),
40352 => conv_std_logic_vector(25120, 16),
40353 => conv_std_logic_vector(25277, 16),
40354 => conv_std_logic_vector(25434, 16),
40355 => conv_std_logic_vector(25591, 16),
40356 => conv_std_logic_vector(25748, 16),
40357 => conv_std_logic_vector(25905, 16),
40358 => conv_std_logic_vector(26062, 16),
40359 => conv_std_logic_vector(26219, 16),
40360 => conv_std_logic_vector(26376, 16),
40361 => conv_std_logic_vector(26533, 16),
40362 => conv_std_logic_vector(26690, 16),
40363 => conv_std_logic_vector(26847, 16),
40364 => conv_std_logic_vector(27004, 16),
40365 => conv_std_logic_vector(27161, 16),
40366 => conv_std_logic_vector(27318, 16),
40367 => conv_std_logic_vector(27475, 16),
40368 => conv_std_logic_vector(27632, 16),
40369 => conv_std_logic_vector(27789, 16),
40370 => conv_std_logic_vector(27946, 16),
40371 => conv_std_logic_vector(28103, 16),
40372 => conv_std_logic_vector(28260, 16),
40373 => conv_std_logic_vector(28417, 16),
40374 => conv_std_logic_vector(28574, 16),
40375 => conv_std_logic_vector(28731, 16),
40376 => conv_std_logic_vector(28888, 16),
40377 => conv_std_logic_vector(29045, 16),
40378 => conv_std_logic_vector(29202, 16),
40379 => conv_std_logic_vector(29359, 16),
40380 => conv_std_logic_vector(29516, 16),
40381 => conv_std_logic_vector(29673, 16),
40382 => conv_std_logic_vector(29830, 16),
40383 => conv_std_logic_vector(29987, 16),
40384 => conv_std_logic_vector(30144, 16),
40385 => conv_std_logic_vector(30301, 16),
40386 => conv_std_logic_vector(30458, 16),
40387 => conv_std_logic_vector(30615, 16),
40388 => conv_std_logic_vector(30772, 16),
40389 => conv_std_logic_vector(30929, 16),
40390 => conv_std_logic_vector(31086, 16),
40391 => conv_std_logic_vector(31243, 16),
40392 => conv_std_logic_vector(31400, 16),
40393 => conv_std_logic_vector(31557, 16),
40394 => conv_std_logic_vector(31714, 16),
40395 => conv_std_logic_vector(31871, 16),
40396 => conv_std_logic_vector(32028, 16),
40397 => conv_std_logic_vector(32185, 16),
40398 => conv_std_logic_vector(32342, 16),
40399 => conv_std_logic_vector(32499, 16),
40400 => conv_std_logic_vector(32656, 16),
40401 => conv_std_logic_vector(32813, 16),
40402 => conv_std_logic_vector(32970, 16),
40403 => conv_std_logic_vector(33127, 16),
40404 => conv_std_logic_vector(33284, 16),
40405 => conv_std_logic_vector(33441, 16),
40406 => conv_std_logic_vector(33598, 16),
40407 => conv_std_logic_vector(33755, 16),
40408 => conv_std_logic_vector(33912, 16),
40409 => conv_std_logic_vector(34069, 16),
40410 => conv_std_logic_vector(34226, 16),
40411 => conv_std_logic_vector(34383, 16),
40412 => conv_std_logic_vector(34540, 16),
40413 => conv_std_logic_vector(34697, 16),
40414 => conv_std_logic_vector(34854, 16),
40415 => conv_std_logic_vector(35011, 16),
40416 => conv_std_logic_vector(35168, 16),
40417 => conv_std_logic_vector(35325, 16),
40418 => conv_std_logic_vector(35482, 16),
40419 => conv_std_logic_vector(35639, 16),
40420 => conv_std_logic_vector(35796, 16),
40421 => conv_std_logic_vector(35953, 16),
40422 => conv_std_logic_vector(36110, 16),
40423 => conv_std_logic_vector(36267, 16),
40424 => conv_std_logic_vector(36424, 16),
40425 => conv_std_logic_vector(36581, 16),
40426 => conv_std_logic_vector(36738, 16),
40427 => conv_std_logic_vector(36895, 16),
40428 => conv_std_logic_vector(37052, 16),
40429 => conv_std_logic_vector(37209, 16),
40430 => conv_std_logic_vector(37366, 16),
40431 => conv_std_logic_vector(37523, 16),
40432 => conv_std_logic_vector(37680, 16),
40433 => conv_std_logic_vector(37837, 16),
40434 => conv_std_logic_vector(37994, 16),
40435 => conv_std_logic_vector(38151, 16),
40436 => conv_std_logic_vector(38308, 16),
40437 => conv_std_logic_vector(38465, 16),
40438 => conv_std_logic_vector(38622, 16),
40439 => conv_std_logic_vector(38779, 16),
40440 => conv_std_logic_vector(38936, 16),
40441 => conv_std_logic_vector(39093, 16),
40442 => conv_std_logic_vector(39250, 16),
40443 => conv_std_logic_vector(39407, 16),
40444 => conv_std_logic_vector(39564, 16),
40445 => conv_std_logic_vector(39721, 16),
40446 => conv_std_logic_vector(39878, 16),
40447 => conv_std_logic_vector(40035, 16),
40448 => conv_std_logic_vector(0, 16),
40449 => conv_std_logic_vector(158, 16),
40450 => conv_std_logic_vector(316, 16),
40451 => conv_std_logic_vector(474, 16),
40452 => conv_std_logic_vector(632, 16),
40453 => conv_std_logic_vector(790, 16),
40454 => conv_std_logic_vector(948, 16),
40455 => conv_std_logic_vector(1106, 16),
40456 => conv_std_logic_vector(1264, 16),
40457 => conv_std_logic_vector(1422, 16),
40458 => conv_std_logic_vector(1580, 16),
40459 => conv_std_logic_vector(1738, 16),
40460 => conv_std_logic_vector(1896, 16),
40461 => conv_std_logic_vector(2054, 16),
40462 => conv_std_logic_vector(2212, 16),
40463 => conv_std_logic_vector(2370, 16),
40464 => conv_std_logic_vector(2528, 16),
40465 => conv_std_logic_vector(2686, 16),
40466 => conv_std_logic_vector(2844, 16),
40467 => conv_std_logic_vector(3002, 16),
40468 => conv_std_logic_vector(3160, 16),
40469 => conv_std_logic_vector(3318, 16),
40470 => conv_std_logic_vector(3476, 16),
40471 => conv_std_logic_vector(3634, 16),
40472 => conv_std_logic_vector(3792, 16),
40473 => conv_std_logic_vector(3950, 16),
40474 => conv_std_logic_vector(4108, 16),
40475 => conv_std_logic_vector(4266, 16),
40476 => conv_std_logic_vector(4424, 16),
40477 => conv_std_logic_vector(4582, 16),
40478 => conv_std_logic_vector(4740, 16),
40479 => conv_std_logic_vector(4898, 16),
40480 => conv_std_logic_vector(5056, 16),
40481 => conv_std_logic_vector(5214, 16),
40482 => conv_std_logic_vector(5372, 16),
40483 => conv_std_logic_vector(5530, 16),
40484 => conv_std_logic_vector(5688, 16),
40485 => conv_std_logic_vector(5846, 16),
40486 => conv_std_logic_vector(6004, 16),
40487 => conv_std_logic_vector(6162, 16),
40488 => conv_std_logic_vector(6320, 16),
40489 => conv_std_logic_vector(6478, 16),
40490 => conv_std_logic_vector(6636, 16),
40491 => conv_std_logic_vector(6794, 16),
40492 => conv_std_logic_vector(6952, 16),
40493 => conv_std_logic_vector(7110, 16),
40494 => conv_std_logic_vector(7268, 16),
40495 => conv_std_logic_vector(7426, 16),
40496 => conv_std_logic_vector(7584, 16),
40497 => conv_std_logic_vector(7742, 16),
40498 => conv_std_logic_vector(7900, 16),
40499 => conv_std_logic_vector(8058, 16),
40500 => conv_std_logic_vector(8216, 16),
40501 => conv_std_logic_vector(8374, 16),
40502 => conv_std_logic_vector(8532, 16),
40503 => conv_std_logic_vector(8690, 16),
40504 => conv_std_logic_vector(8848, 16),
40505 => conv_std_logic_vector(9006, 16),
40506 => conv_std_logic_vector(9164, 16),
40507 => conv_std_logic_vector(9322, 16),
40508 => conv_std_logic_vector(9480, 16),
40509 => conv_std_logic_vector(9638, 16),
40510 => conv_std_logic_vector(9796, 16),
40511 => conv_std_logic_vector(9954, 16),
40512 => conv_std_logic_vector(10112, 16),
40513 => conv_std_logic_vector(10270, 16),
40514 => conv_std_logic_vector(10428, 16),
40515 => conv_std_logic_vector(10586, 16),
40516 => conv_std_logic_vector(10744, 16),
40517 => conv_std_logic_vector(10902, 16),
40518 => conv_std_logic_vector(11060, 16),
40519 => conv_std_logic_vector(11218, 16),
40520 => conv_std_logic_vector(11376, 16),
40521 => conv_std_logic_vector(11534, 16),
40522 => conv_std_logic_vector(11692, 16),
40523 => conv_std_logic_vector(11850, 16),
40524 => conv_std_logic_vector(12008, 16),
40525 => conv_std_logic_vector(12166, 16),
40526 => conv_std_logic_vector(12324, 16),
40527 => conv_std_logic_vector(12482, 16),
40528 => conv_std_logic_vector(12640, 16),
40529 => conv_std_logic_vector(12798, 16),
40530 => conv_std_logic_vector(12956, 16),
40531 => conv_std_logic_vector(13114, 16),
40532 => conv_std_logic_vector(13272, 16),
40533 => conv_std_logic_vector(13430, 16),
40534 => conv_std_logic_vector(13588, 16),
40535 => conv_std_logic_vector(13746, 16),
40536 => conv_std_logic_vector(13904, 16),
40537 => conv_std_logic_vector(14062, 16),
40538 => conv_std_logic_vector(14220, 16),
40539 => conv_std_logic_vector(14378, 16),
40540 => conv_std_logic_vector(14536, 16),
40541 => conv_std_logic_vector(14694, 16),
40542 => conv_std_logic_vector(14852, 16),
40543 => conv_std_logic_vector(15010, 16),
40544 => conv_std_logic_vector(15168, 16),
40545 => conv_std_logic_vector(15326, 16),
40546 => conv_std_logic_vector(15484, 16),
40547 => conv_std_logic_vector(15642, 16),
40548 => conv_std_logic_vector(15800, 16),
40549 => conv_std_logic_vector(15958, 16),
40550 => conv_std_logic_vector(16116, 16),
40551 => conv_std_logic_vector(16274, 16),
40552 => conv_std_logic_vector(16432, 16),
40553 => conv_std_logic_vector(16590, 16),
40554 => conv_std_logic_vector(16748, 16),
40555 => conv_std_logic_vector(16906, 16),
40556 => conv_std_logic_vector(17064, 16),
40557 => conv_std_logic_vector(17222, 16),
40558 => conv_std_logic_vector(17380, 16),
40559 => conv_std_logic_vector(17538, 16),
40560 => conv_std_logic_vector(17696, 16),
40561 => conv_std_logic_vector(17854, 16),
40562 => conv_std_logic_vector(18012, 16),
40563 => conv_std_logic_vector(18170, 16),
40564 => conv_std_logic_vector(18328, 16),
40565 => conv_std_logic_vector(18486, 16),
40566 => conv_std_logic_vector(18644, 16),
40567 => conv_std_logic_vector(18802, 16),
40568 => conv_std_logic_vector(18960, 16),
40569 => conv_std_logic_vector(19118, 16),
40570 => conv_std_logic_vector(19276, 16),
40571 => conv_std_logic_vector(19434, 16),
40572 => conv_std_logic_vector(19592, 16),
40573 => conv_std_logic_vector(19750, 16),
40574 => conv_std_logic_vector(19908, 16),
40575 => conv_std_logic_vector(20066, 16),
40576 => conv_std_logic_vector(20224, 16),
40577 => conv_std_logic_vector(20382, 16),
40578 => conv_std_logic_vector(20540, 16),
40579 => conv_std_logic_vector(20698, 16),
40580 => conv_std_logic_vector(20856, 16),
40581 => conv_std_logic_vector(21014, 16),
40582 => conv_std_logic_vector(21172, 16),
40583 => conv_std_logic_vector(21330, 16),
40584 => conv_std_logic_vector(21488, 16),
40585 => conv_std_logic_vector(21646, 16),
40586 => conv_std_logic_vector(21804, 16),
40587 => conv_std_logic_vector(21962, 16),
40588 => conv_std_logic_vector(22120, 16),
40589 => conv_std_logic_vector(22278, 16),
40590 => conv_std_logic_vector(22436, 16),
40591 => conv_std_logic_vector(22594, 16),
40592 => conv_std_logic_vector(22752, 16),
40593 => conv_std_logic_vector(22910, 16),
40594 => conv_std_logic_vector(23068, 16),
40595 => conv_std_logic_vector(23226, 16),
40596 => conv_std_logic_vector(23384, 16),
40597 => conv_std_logic_vector(23542, 16),
40598 => conv_std_logic_vector(23700, 16),
40599 => conv_std_logic_vector(23858, 16),
40600 => conv_std_logic_vector(24016, 16),
40601 => conv_std_logic_vector(24174, 16),
40602 => conv_std_logic_vector(24332, 16),
40603 => conv_std_logic_vector(24490, 16),
40604 => conv_std_logic_vector(24648, 16),
40605 => conv_std_logic_vector(24806, 16),
40606 => conv_std_logic_vector(24964, 16),
40607 => conv_std_logic_vector(25122, 16),
40608 => conv_std_logic_vector(25280, 16),
40609 => conv_std_logic_vector(25438, 16),
40610 => conv_std_logic_vector(25596, 16),
40611 => conv_std_logic_vector(25754, 16),
40612 => conv_std_logic_vector(25912, 16),
40613 => conv_std_logic_vector(26070, 16),
40614 => conv_std_logic_vector(26228, 16),
40615 => conv_std_logic_vector(26386, 16),
40616 => conv_std_logic_vector(26544, 16),
40617 => conv_std_logic_vector(26702, 16),
40618 => conv_std_logic_vector(26860, 16),
40619 => conv_std_logic_vector(27018, 16),
40620 => conv_std_logic_vector(27176, 16),
40621 => conv_std_logic_vector(27334, 16),
40622 => conv_std_logic_vector(27492, 16),
40623 => conv_std_logic_vector(27650, 16),
40624 => conv_std_logic_vector(27808, 16),
40625 => conv_std_logic_vector(27966, 16),
40626 => conv_std_logic_vector(28124, 16),
40627 => conv_std_logic_vector(28282, 16),
40628 => conv_std_logic_vector(28440, 16),
40629 => conv_std_logic_vector(28598, 16),
40630 => conv_std_logic_vector(28756, 16),
40631 => conv_std_logic_vector(28914, 16),
40632 => conv_std_logic_vector(29072, 16),
40633 => conv_std_logic_vector(29230, 16),
40634 => conv_std_logic_vector(29388, 16),
40635 => conv_std_logic_vector(29546, 16),
40636 => conv_std_logic_vector(29704, 16),
40637 => conv_std_logic_vector(29862, 16),
40638 => conv_std_logic_vector(30020, 16),
40639 => conv_std_logic_vector(30178, 16),
40640 => conv_std_logic_vector(30336, 16),
40641 => conv_std_logic_vector(30494, 16),
40642 => conv_std_logic_vector(30652, 16),
40643 => conv_std_logic_vector(30810, 16),
40644 => conv_std_logic_vector(30968, 16),
40645 => conv_std_logic_vector(31126, 16),
40646 => conv_std_logic_vector(31284, 16),
40647 => conv_std_logic_vector(31442, 16),
40648 => conv_std_logic_vector(31600, 16),
40649 => conv_std_logic_vector(31758, 16),
40650 => conv_std_logic_vector(31916, 16),
40651 => conv_std_logic_vector(32074, 16),
40652 => conv_std_logic_vector(32232, 16),
40653 => conv_std_logic_vector(32390, 16),
40654 => conv_std_logic_vector(32548, 16),
40655 => conv_std_logic_vector(32706, 16),
40656 => conv_std_logic_vector(32864, 16),
40657 => conv_std_logic_vector(33022, 16),
40658 => conv_std_logic_vector(33180, 16),
40659 => conv_std_logic_vector(33338, 16),
40660 => conv_std_logic_vector(33496, 16),
40661 => conv_std_logic_vector(33654, 16),
40662 => conv_std_logic_vector(33812, 16),
40663 => conv_std_logic_vector(33970, 16),
40664 => conv_std_logic_vector(34128, 16),
40665 => conv_std_logic_vector(34286, 16),
40666 => conv_std_logic_vector(34444, 16),
40667 => conv_std_logic_vector(34602, 16),
40668 => conv_std_logic_vector(34760, 16),
40669 => conv_std_logic_vector(34918, 16),
40670 => conv_std_logic_vector(35076, 16),
40671 => conv_std_logic_vector(35234, 16),
40672 => conv_std_logic_vector(35392, 16),
40673 => conv_std_logic_vector(35550, 16),
40674 => conv_std_logic_vector(35708, 16),
40675 => conv_std_logic_vector(35866, 16),
40676 => conv_std_logic_vector(36024, 16),
40677 => conv_std_logic_vector(36182, 16),
40678 => conv_std_logic_vector(36340, 16),
40679 => conv_std_logic_vector(36498, 16),
40680 => conv_std_logic_vector(36656, 16),
40681 => conv_std_logic_vector(36814, 16),
40682 => conv_std_logic_vector(36972, 16),
40683 => conv_std_logic_vector(37130, 16),
40684 => conv_std_logic_vector(37288, 16),
40685 => conv_std_logic_vector(37446, 16),
40686 => conv_std_logic_vector(37604, 16),
40687 => conv_std_logic_vector(37762, 16),
40688 => conv_std_logic_vector(37920, 16),
40689 => conv_std_logic_vector(38078, 16),
40690 => conv_std_logic_vector(38236, 16),
40691 => conv_std_logic_vector(38394, 16),
40692 => conv_std_logic_vector(38552, 16),
40693 => conv_std_logic_vector(38710, 16),
40694 => conv_std_logic_vector(38868, 16),
40695 => conv_std_logic_vector(39026, 16),
40696 => conv_std_logic_vector(39184, 16),
40697 => conv_std_logic_vector(39342, 16),
40698 => conv_std_logic_vector(39500, 16),
40699 => conv_std_logic_vector(39658, 16),
40700 => conv_std_logic_vector(39816, 16),
40701 => conv_std_logic_vector(39974, 16),
40702 => conv_std_logic_vector(40132, 16),
40703 => conv_std_logic_vector(40290, 16),
40704 => conv_std_logic_vector(0, 16),
40705 => conv_std_logic_vector(159, 16),
40706 => conv_std_logic_vector(318, 16),
40707 => conv_std_logic_vector(477, 16),
40708 => conv_std_logic_vector(636, 16),
40709 => conv_std_logic_vector(795, 16),
40710 => conv_std_logic_vector(954, 16),
40711 => conv_std_logic_vector(1113, 16),
40712 => conv_std_logic_vector(1272, 16),
40713 => conv_std_logic_vector(1431, 16),
40714 => conv_std_logic_vector(1590, 16),
40715 => conv_std_logic_vector(1749, 16),
40716 => conv_std_logic_vector(1908, 16),
40717 => conv_std_logic_vector(2067, 16),
40718 => conv_std_logic_vector(2226, 16),
40719 => conv_std_logic_vector(2385, 16),
40720 => conv_std_logic_vector(2544, 16),
40721 => conv_std_logic_vector(2703, 16),
40722 => conv_std_logic_vector(2862, 16),
40723 => conv_std_logic_vector(3021, 16),
40724 => conv_std_logic_vector(3180, 16),
40725 => conv_std_logic_vector(3339, 16),
40726 => conv_std_logic_vector(3498, 16),
40727 => conv_std_logic_vector(3657, 16),
40728 => conv_std_logic_vector(3816, 16),
40729 => conv_std_logic_vector(3975, 16),
40730 => conv_std_logic_vector(4134, 16),
40731 => conv_std_logic_vector(4293, 16),
40732 => conv_std_logic_vector(4452, 16),
40733 => conv_std_logic_vector(4611, 16),
40734 => conv_std_logic_vector(4770, 16),
40735 => conv_std_logic_vector(4929, 16),
40736 => conv_std_logic_vector(5088, 16),
40737 => conv_std_logic_vector(5247, 16),
40738 => conv_std_logic_vector(5406, 16),
40739 => conv_std_logic_vector(5565, 16),
40740 => conv_std_logic_vector(5724, 16),
40741 => conv_std_logic_vector(5883, 16),
40742 => conv_std_logic_vector(6042, 16),
40743 => conv_std_logic_vector(6201, 16),
40744 => conv_std_logic_vector(6360, 16),
40745 => conv_std_logic_vector(6519, 16),
40746 => conv_std_logic_vector(6678, 16),
40747 => conv_std_logic_vector(6837, 16),
40748 => conv_std_logic_vector(6996, 16),
40749 => conv_std_logic_vector(7155, 16),
40750 => conv_std_logic_vector(7314, 16),
40751 => conv_std_logic_vector(7473, 16),
40752 => conv_std_logic_vector(7632, 16),
40753 => conv_std_logic_vector(7791, 16),
40754 => conv_std_logic_vector(7950, 16),
40755 => conv_std_logic_vector(8109, 16),
40756 => conv_std_logic_vector(8268, 16),
40757 => conv_std_logic_vector(8427, 16),
40758 => conv_std_logic_vector(8586, 16),
40759 => conv_std_logic_vector(8745, 16),
40760 => conv_std_logic_vector(8904, 16),
40761 => conv_std_logic_vector(9063, 16),
40762 => conv_std_logic_vector(9222, 16),
40763 => conv_std_logic_vector(9381, 16),
40764 => conv_std_logic_vector(9540, 16),
40765 => conv_std_logic_vector(9699, 16),
40766 => conv_std_logic_vector(9858, 16),
40767 => conv_std_logic_vector(10017, 16),
40768 => conv_std_logic_vector(10176, 16),
40769 => conv_std_logic_vector(10335, 16),
40770 => conv_std_logic_vector(10494, 16),
40771 => conv_std_logic_vector(10653, 16),
40772 => conv_std_logic_vector(10812, 16),
40773 => conv_std_logic_vector(10971, 16),
40774 => conv_std_logic_vector(11130, 16),
40775 => conv_std_logic_vector(11289, 16),
40776 => conv_std_logic_vector(11448, 16),
40777 => conv_std_logic_vector(11607, 16),
40778 => conv_std_logic_vector(11766, 16),
40779 => conv_std_logic_vector(11925, 16),
40780 => conv_std_logic_vector(12084, 16),
40781 => conv_std_logic_vector(12243, 16),
40782 => conv_std_logic_vector(12402, 16),
40783 => conv_std_logic_vector(12561, 16),
40784 => conv_std_logic_vector(12720, 16),
40785 => conv_std_logic_vector(12879, 16),
40786 => conv_std_logic_vector(13038, 16),
40787 => conv_std_logic_vector(13197, 16),
40788 => conv_std_logic_vector(13356, 16),
40789 => conv_std_logic_vector(13515, 16),
40790 => conv_std_logic_vector(13674, 16),
40791 => conv_std_logic_vector(13833, 16),
40792 => conv_std_logic_vector(13992, 16),
40793 => conv_std_logic_vector(14151, 16),
40794 => conv_std_logic_vector(14310, 16),
40795 => conv_std_logic_vector(14469, 16),
40796 => conv_std_logic_vector(14628, 16),
40797 => conv_std_logic_vector(14787, 16),
40798 => conv_std_logic_vector(14946, 16),
40799 => conv_std_logic_vector(15105, 16),
40800 => conv_std_logic_vector(15264, 16),
40801 => conv_std_logic_vector(15423, 16),
40802 => conv_std_logic_vector(15582, 16),
40803 => conv_std_logic_vector(15741, 16),
40804 => conv_std_logic_vector(15900, 16),
40805 => conv_std_logic_vector(16059, 16),
40806 => conv_std_logic_vector(16218, 16),
40807 => conv_std_logic_vector(16377, 16),
40808 => conv_std_logic_vector(16536, 16),
40809 => conv_std_logic_vector(16695, 16),
40810 => conv_std_logic_vector(16854, 16),
40811 => conv_std_logic_vector(17013, 16),
40812 => conv_std_logic_vector(17172, 16),
40813 => conv_std_logic_vector(17331, 16),
40814 => conv_std_logic_vector(17490, 16),
40815 => conv_std_logic_vector(17649, 16),
40816 => conv_std_logic_vector(17808, 16),
40817 => conv_std_logic_vector(17967, 16),
40818 => conv_std_logic_vector(18126, 16),
40819 => conv_std_logic_vector(18285, 16),
40820 => conv_std_logic_vector(18444, 16),
40821 => conv_std_logic_vector(18603, 16),
40822 => conv_std_logic_vector(18762, 16),
40823 => conv_std_logic_vector(18921, 16),
40824 => conv_std_logic_vector(19080, 16),
40825 => conv_std_logic_vector(19239, 16),
40826 => conv_std_logic_vector(19398, 16),
40827 => conv_std_logic_vector(19557, 16),
40828 => conv_std_logic_vector(19716, 16),
40829 => conv_std_logic_vector(19875, 16),
40830 => conv_std_logic_vector(20034, 16),
40831 => conv_std_logic_vector(20193, 16),
40832 => conv_std_logic_vector(20352, 16),
40833 => conv_std_logic_vector(20511, 16),
40834 => conv_std_logic_vector(20670, 16),
40835 => conv_std_logic_vector(20829, 16),
40836 => conv_std_logic_vector(20988, 16),
40837 => conv_std_logic_vector(21147, 16),
40838 => conv_std_logic_vector(21306, 16),
40839 => conv_std_logic_vector(21465, 16),
40840 => conv_std_logic_vector(21624, 16),
40841 => conv_std_logic_vector(21783, 16),
40842 => conv_std_logic_vector(21942, 16),
40843 => conv_std_logic_vector(22101, 16),
40844 => conv_std_logic_vector(22260, 16),
40845 => conv_std_logic_vector(22419, 16),
40846 => conv_std_logic_vector(22578, 16),
40847 => conv_std_logic_vector(22737, 16),
40848 => conv_std_logic_vector(22896, 16),
40849 => conv_std_logic_vector(23055, 16),
40850 => conv_std_logic_vector(23214, 16),
40851 => conv_std_logic_vector(23373, 16),
40852 => conv_std_logic_vector(23532, 16),
40853 => conv_std_logic_vector(23691, 16),
40854 => conv_std_logic_vector(23850, 16),
40855 => conv_std_logic_vector(24009, 16),
40856 => conv_std_logic_vector(24168, 16),
40857 => conv_std_logic_vector(24327, 16),
40858 => conv_std_logic_vector(24486, 16),
40859 => conv_std_logic_vector(24645, 16),
40860 => conv_std_logic_vector(24804, 16),
40861 => conv_std_logic_vector(24963, 16),
40862 => conv_std_logic_vector(25122, 16),
40863 => conv_std_logic_vector(25281, 16),
40864 => conv_std_logic_vector(25440, 16),
40865 => conv_std_logic_vector(25599, 16),
40866 => conv_std_logic_vector(25758, 16),
40867 => conv_std_logic_vector(25917, 16),
40868 => conv_std_logic_vector(26076, 16),
40869 => conv_std_logic_vector(26235, 16),
40870 => conv_std_logic_vector(26394, 16),
40871 => conv_std_logic_vector(26553, 16),
40872 => conv_std_logic_vector(26712, 16),
40873 => conv_std_logic_vector(26871, 16),
40874 => conv_std_logic_vector(27030, 16),
40875 => conv_std_logic_vector(27189, 16),
40876 => conv_std_logic_vector(27348, 16),
40877 => conv_std_logic_vector(27507, 16),
40878 => conv_std_logic_vector(27666, 16),
40879 => conv_std_logic_vector(27825, 16),
40880 => conv_std_logic_vector(27984, 16),
40881 => conv_std_logic_vector(28143, 16),
40882 => conv_std_logic_vector(28302, 16),
40883 => conv_std_logic_vector(28461, 16),
40884 => conv_std_logic_vector(28620, 16),
40885 => conv_std_logic_vector(28779, 16),
40886 => conv_std_logic_vector(28938, 16),
40887 => conv_std_logic_vector(29097, 16),
40888 => conv_std_logic_vector(29256, 16),
40889 => conv_std_logic_vector(29415, 16),
40890 => conv_std_logic_vector(29574, 16),
40891 => conv_std_logic_vector(29733, 16),
40892 => conv_std_logic_vector(29892, 16),
40893 => conv_std_logic_vector(30051, 16),
40894 => conv_std_logic_vector(30210, 16),
40895 => conv_std_logic_vector(30369, 16),
40896 => conv_std_logic_vector(30528, 16),
40897 => conv_std_logic_vector(30687, 16),
40898 => conv_std_logic_vector(30846, 16),
40899 => conv_std_logic_vector(31005, 16),
40900 => conv_std_logic_vector(31164, 16),
40901 => conv_std_logic_vector(31323, 16),
40902 => conv_std_logic_vector(31482, 16),
40903 => conv_std_logic_vector(31641, 16),
40904 => conv_std_logic_vector(31800, 16),
40905 => conv_std_logic_vector(31959, 16),
40906 => conv_std_logic_vector(32118, 16),
40907 => conv_std_logic_vector(32277, 16),
40908 => conv_std_logic_vector(32436, 16),
40909 => conv_std_logic_vector(32595, 16),
40910 => conv_std_logic_vector(32754, 16),
40911 => conv_std_logic_vector(32913, 16),
40912 => conv_std_logic_vector(33072, 16),
40913 => conv_std_logic_vector(33231, 16),
40914 => conv_std_logic_vector(33390, 16),
40915 => conv_std_logic_vector(33549, 16),
40916 => conv_std_logic_vector(33708, 16),
40917 => conv_std_logic_vector(33867, 16),
40918 => conv_std_logic_vector(34026, 16),
40919 => conv_std_logic_vector(34185, 16),
40920 => conv_std_logic_vector(34344, 16),
40921 => conv_std_logic_vector(34503, 16),
40922 => conv_std_logic_vector(34662, 16),
40923 => conv_std_logic_vector(34821, 16),
40924 => conv_std_logic_vector(34980, 16),
40925 => conv_std_logic_vector(35139, 16),
40926 => conv_std_logic_vector(35298, 16),
40927 => conv_std_logic_vector(35457, 16),
40928 => conv_std_logic_vector(35616, 16),
40929 => conv_std_logic_vector(35775, 16),
40930 => conv_std_logic_vector(35934, 16),
40931 => conv_std_logic_vector(36093, 16),
40932 => conv_std_logic_vector(36252, 16),
40933 => conv_std_logic_vector(36411, 16),
40934 => conv_std_logic_vector(36570, 16),
40935 => conv_std_logic_vector(36729, 16),
40936 => conv_std_logic_vector(36888, 16),
40937 => conv_std_logic_vector(37047, 16),
40938 => conv_std_logic_vector(37206, 16),
40939 => conv_std_logic_vector(37365, 16),
40940 => conv_std_logic_vector(37524, 16),
40941 => conv_std_logic_vector(37683, 16),
40942 => conv_std_logic_vector(37842, 16),
40943 => conv_std_logic_vector(38001, 16),
40944 => conv_std_logic_vector(38160, 16),
40945 => conv_std_logic_vector(38319, 16),
40946 => conv_std_logic_vector(38478, 16),
40947 => conv_std_logic_vector(38637, 16),
40948 => conv_std_logic_vector(38796, 16),
40949 => conv_std_logic_vector(38955, 16),
40950 => conv_std_logic_vector(39114, 16),
40951 => conv_std_logic_vector(39273, 16),
40952 => conv_std_logic_vector(39432, 16),
40953 => conv_std_logic_vector(39591, 16),
40954 => conv_std_logic_vector(39750, 16),
40955 => conv_std_logic_vector(39909, 16),
40956 => conv_std_logic_vector(40068, 16),
40957 => conv_std_logic_vector(40227, 16),
40958 => conv_std_logic_vector(40386, 16),
40959 => conv_std_logic_vector(40545, 16),
40960 => conv_std_logic_vector(0, 16),
40961 => conv_std_logic_vector(160, 16),
40962 => conv_std_logic_vector(320, 16),
40963 => conv_std_logic_vector(480, 16),
40964 => conv_std_logic_vector(640, 16),
40965 => conv_std_logic_vector(800, 16),
40966 => conv_std_logic_vector(960, 16),
40967 => conv_std_logic_vector(1120, 16),
40968 => conv_std_logic_vector(1280, 16),
40969 => conv_std_logic_vector(1440, 16),
40970 => conv_std_logic_vector(1600, 16),
40971 => conv_std_logic_vector(1760, 16),
40972 => conv_std_logic_vector(1920, 16),
40973 => conv_std_logic_vector(2080, 16),
40974 => conv_std_logic_vector(2240, 16),
40975 => conv_std_logic_vector(2400, 16),
40976 => conv_std_logic_vector(2560, 16),
40977 => conv_std_logic_vector(2720, 16),
40978 => conv_std_logic_vector(2880, 16),
40979 => conv_std_logic_vector(3040, 16),
40980 => conv_std_logic_vector(3200, 16),
40981 => conv_std_logic_vector(3360, 16),
40982 => conv_std_logic_vector(3520, 16),
40983 => conv_std_logic_vector(3680, 16),
40984 => conv_std_logic_vector(3840, 16),
40985 => conv_std_logic_vector(4000, 16),
40986 => conv_std_logic_vector(4160, 16),
40987 => conv_std_logic_vector(4320, 16),
40988 => conv_std_logic_vector(4480, 16),
40989 => conv_std_logic_vector(4640, 16),
40990 => conv_std_logic_vector(4800, 16),
40991 => conv_std_logic_vector(4960, 16),
40992 => conv_std_logic_vector(5120, 16),
40993 => conv_std_logic_vector(5280, 16),
40994 => conv_std_logic_vector(5440, 16),
40995 => conv_std_logic_vector(5600, 16),
40996 => conv_std_logic_vector(5760, 16),
40997 => conv_std_logic_vector(5920, 16),
40998 => conv_std_logic_vector(6080, 16),
40999 => conv_std_logic_vector(6240, 16),
41000 => conv_std_logic_vector(6400, 16),
41001 => conv_std_logic_vector(6560, 16),
41002 => conv_std_logic_vector(6720, 16),
41003 => conv_std_logic_vector(6880, 16),
41004 => conv_std_logic_vector(7040, 16),
41005 => conv_std_logic_vector(7200, 16),
41006 => conv_std_logic_vector(7360, 16),
41007 => conv_std_logic_vector(7520, 16),
41008 => conv_std_logic_vector(7680, 16),
41009 => conv_std_logic_vector(7840, 16),
41010 => conv_std_logic_vector(8000, 16),
41011 => conv_std_logic_vector(8160, 16),
41012 => conv_std_logic_vector(8320, 16),
41013 => conv_std_logic_vector(8480, 16),
41014 => conv_std_logic_vector(8640, 16),
41015 => conv_std_logic_vector(8800, 16),
41016 => conv_std_logic_vector(8960, 16),
41017 => conv_std_logic_vector(9120, 16),
41018 => conv_std_logic_vector(9280, 16),
41019 => conv_std_logic_vector(9440, 16),
41020 => conv_std_logic_vector(9600, 16),
41021 => conv_std_logic_vector(9760, 16),
41022 => conv_std_logic_vector(9920, 16),
41023 => conv_std_logic_vector(10080, 16),
41024 => conv_std_logic_vector(10240, 16),
41025 => conv_std_logic_vector(10400, 16),
41026 => conv_std_logic_vector(10560, 16),
41027 => conv_std_logic_vector(10720, 16),
41028 => conv_std_logic_vector(10880, 16),
41029 => conv_std_logic_vector(11040, 16),
41030 => conv_std_logic_vector(11200, 16),
41031 => conv_std_logic_vector(11360, 16),
41032 => conv_std_logic_vector(11520, 16),
41033 => conv_std_logic_vector(11680, 16),
41034 => conv_std_logic_vector(11840, 16),
41035 => conv_std_logic_vector(12000, 16),
41036 => conv_std_logic_vector(12160, 16),
41037 => conv_std_logic_vector(12320, 16),
41038 => conv_std_logic_vector(12480, 16),
41039 => conv_std_logic_vector(12640, 16),
41040 => conv_std_logic_vector(12800, 16),
41041 => conv_std_logic_vector(12960, 16),
41042 => conv_std_logic_vector(13120, 16),
41043 => conv_std_logic_vector(13280, 16),
41044 => conv_std_logic_vector(13440, 16),
41045 => conv_std_logic_vector(13600, 16),
41046 => conv_std_logic_vector(13760, 16),
41047 => conv_std_logic_vector(13920, 16),
41048 => conv_std_logic_vector(14080, 16),
41049 => conv_std_logic_vector(14240, 16),
41050 => conv_std_logic_vector(14400, 16),
41051 => conv_std_logic_vector(14560, 16),
41052 => conv_std_logic_vector(14720, 16),
41053 => conv_std_logic_vector(14880, 16),
41054 => conv_std_logic_vector(15040, 16),
41055 => conv_std_logic_vector(15200, 16),
41056 => conv_std_logic_vector(15360, 16),
41057 => conv_std_logic_vector(15520, 16),
41058 => conv_std_logic_vector(15680, 16),
41059 => conv_std_logic_vector(15840, 16),
41060 => conv_std_logic_vector(16000, 16),
41061 => conv_std_logic_vector(16160, 16),
41062 => conv_std_logic_vector(16320, 16),
41063 => conv_std_logic_vector(16480, 16),
41064 => conv_std_logic_vector(16640, 16),
41065 => conv_std_logic_vector(16800, 16),
41066 => conv_std_logic_vector(16960, 16),
41067 => conv_std_logic_vector(17120, 16),
41068 => conv_std_logic_vector(17280, 16),
41069 => conv_std_logic_vector(17440, 16),
41070 => conv_std_logic_vector(17600, 16),
41071 => conv_std_logic_vector(17760, 16),
41072 => conv_std_logic_vector(17920, 16),
41073 => conv_std_logic_vector(18080, 16),
41074 => conv_std_logic_vector(18240, 16),
41075 => conv_std_logic_vector(18400, 16),
41076 => conv_std_logic_vector(18560, 16),
41077 => conv_std_logic_vector(18720, 16),
41078 => conv_std_logic_vector(18880, 16),
41079 => conv_std_logic_vector(19040, 16),
41080 => conv_std_logic_vector(19200, 16),
41081 => conv_std_logic_vector(19360, 16),
41082 => conv_std_logic_vector(19520, 16),
41083 => conv_std_logic_vector(19680, 16),
41084 => conv_std_logic_vector(19840, 16),
41085 => conv_std_logic_vector(20000, 16),
41086 => conv_std_logic_vector(20160, 16),
41087 => conv_std_logic_vector(20320, 16),
41088 => conv_std_logic_vector(20480, 16),
41089 => conv_std_logic_vector(20640, 16),
41090 => conv_std_logic_vector(20800, 16),
41091 => conv_std_logic_vector(20960, 16),
41092 => conv_std_logic_vector(21120, 16),
41093 => conv_std_logic_vector(21280, 16),
41094 => conv_std_logic_vector(21440, 16),
41095 => conv_std_logic_vector(21600, 16),
41096 => conv_std_logic_vector(21760, 16),
41097 => conv_std_logic_vector(21920, 16),
41098 => conv_std_logic_vector(22080, 16),
41099 => conv_std_logic_vector(22240, 16),
41100 => conv_std_logic_vector(22400, 16),
41101 => conv_std_logic_vector(22560, 16),
41102 => conv_std_logic_vector(22720, 16),
41103 => conv_std_logic_vector(22880, 16),
41104 => conv_std_logic_vector(23040, 16),
41105 => conv_std_logic_vector(23200, 16),
41106 => conv_std_logic_vector(23360, 16),
41107 => conv_std_logic_vector(23520, 16),
41108 => conv_std_logic_vector(23680, 16),
41109 => conv_std_logic_vector(23840, 16),
41110 => conv_std_logic_vector(24000, 16),
41111 => conv_std_logic_vector(24160, 16),
41112 => conv_std_logic_vector(24320, 16),
41113 => conv_std_logic_vector(24480, 16),
41114 => conv_std_logic_vector(24640, 16),
41115 => conv_std_logic_vector(24800, 16),
41116 => conv_std_logic_vector(24960, 16),
41117 => conv_std_logic_vector(25120, 16),
41118 => conv_std_logic_vector(25280, 16),
41119 => conv_std_logic_vector(25440, 16),
41120 => conv_std_logic_vector(25600, 16),
41121 => conv_std_logic_vector(25760, 16),
41122 => conv_std_logic_vector(25920, 16),
41123 => conv_std_logic_vector(26080, 16),
41124 => conv_std_logic_vector(26240, 16),
41125 => conv_std_logic_vector(26400, 16),
41126 => conv_std_logic_vector(26560, 16),
41127 => conv_std_logic_vector(26720, 16),
41128 => conv_std_logic_vector(26880, 16),
41129 => conv_std_logic_vector(27040, 16),
41130 => conv_std_logic_vector(27200, 16),
41131 => conv_std_logic_vector(27360, 16),
41132 => conv_std_logic_vector(27520, 16),
41133 => conv_std_logic_vector(27680, 16),
41134 => conv_std_logic_vector(27840, 16),
41135 => conv_std_logic_vector(28000, 16),
41136 => conv_std_logic_vector(28160, 16),
41137 => conv_std_logic_vector(28320, 16),
41138 => conv_std_logic_vector(28480, 16),
41139 => conv_std_logic_vector(28640, 16),
41140 => conv_std_logic_vector(28800, 16),
41141 => conv_std_logic_vector(28960, 16),
41142 => conv_std_logic_vector(29120, 16),
41143 => conv_std_logic_vector(29280, 16),
41144 => conv_std_logic_vector(29440, 16),
41145 => conv_std_logic_vector(29600, 16),
41146 => conv_std_logic_vector(29760, 16),
41147 => conv_std_logic_vector(29920, 16),
41148 => conv_std_logic_vector(30080, 16),
41149 => conv_std_logic_vector(30240, 16),
41150 => conv_std_logic_vector(30400, 16),
41151 => conv_std_logic_vector(30560, 16),
41152 => conv_std_logic_vector(30720, 16),
41153 => conv_std_logic_vector(30880, 16),
41154 => conv_std_logic_vector(31040, 16),
41155 => conv_std_logic_vector(31200, 16),
41156 => conv_std_logic_vector(31360, 16),
41157 => conv_std_logic_vector(31520, 16),
41158 => conv_std_logic_vector(31680, 16),
41159 => conv_std_logic_vector(31840, 16),
41160 => conv_std_logic_vector(32000, 16),
41161 => conv_std_logic_vector(32160, 16),
41162 => conv_std_logic_vector(32320, 16),
41163 => conv_std_logic_vector(32480, 16),
41164 => conv_std_logic_vector(32640, 16),
41165 => conv_std_logic_vector(32800, 16),
41166 => conv_std_logic_vector(32960, 16),
41167 => conv_std_logic_vector(33120, 16),
41168 => conv_std_logic_vector(33280, 16),
41169 => conv_std_logic_vector(33440, 16),
41170 => conv_std_logic_vector(33600, 16),
41171 => conv_std_logic_vector(33760, 16),
41172 => conv_std_logic_vector(33920, 16),
41173 => conv_std_logic_vector(34080, 16),
41174 => conv_std_logic_vector(34240, 16),
41175 => conv_std_logic_vector(34400, 16),
41176 => conv_std_logic_vector(34560, 16),
41177 => conv_std_logic_vector(34720, 16),
41178 => conv_std_logic_vector(34880, 16),
41179 => conv_std_logic_vector(35040, 16),
41180 => conv_std_logic_vector(35200, 16),
41181 => conv_std_logic_vector(35360, 16),
41182 => conv_std_logic_vector(35520, 16),
41183 => conv_std_logic_vector(35680, 16),
41184 => conv_std_logic_vector(35840, 16),
41185 => conv_std_logic_vector(36000, 16),
41186 => conv_std_logic_vector(36160, 16),
41187 => conv_std_logic_vector(36320, 16),
41188 => conv_std_logic_vector(36480, 16),
41189 => conv_std_logic_vector(36640, 16),
41190 => conv_std_logic_vector(36800, 16),
41191 => conv_std_logic_vector(36960, 16),
41192 => conv_std_logic_vector(37120, 16),
41193 => conv_std_logic_vector(37280, 16),
41194 => conv_std_logic_vector(37440, 16),
41195 => conv_std_logic_vector(37600, 16),
41196 => conv_std_logic_vector(37760, 16),
41197 => conv_std_logic_vector(37920, 16),
41198 => conv_std_logic_vector(38080, 16),
41199 => conv_std_logic_vector(38240, 16),
41200 => conv_std_logic_vector(38400, 16),
41201 => conv_std_logic_vector(38560, 16),
41202 => conv_std_logic_vector(38720, 16),
41203 => conv_std_logic_vector(38880, 16),
41204 => conv_std_logic_vector(39040, 16),
41205 => conv_std_logic_vector(39200, 16),
41206 => conv_std_logic_vector(39360, 16),
41207 => conv_std_logic_vector(39520, 16),
41208 => conv_std_logic_vector(39680, 16),
41209 => conv_std_logic_vector(39840, 16),
41210 => conv_std_logic_vector(40000, 16),
41211 => conv_std_logic_vector(40160, 16),
41212 => conv_std_logic_vector(40320, 16),
41213 => conv_std_logic_vector(40480, 16),
41214 => conv_std_logic_vector(40640, 16),
41215 => conv_std_logic_vector(40800, 16),
41216 => conv_std_logic_vector(0, 16),
41217 => conv_std_logic_vector(161, 16),
41218 => conv_std_logic_vector(322, 16),
41219 => conv_std_logic_vector(483, 16),
41220 => conv_std_logic_vector(644, 16),
41221 => conv_std_logic_vector(805, 16),
41222 => conv_std_logic_vector(966, 16),
41223 => conv_std_logic_vector(1127, 16),
41224 => conv_std_logic_vector(1288, 16),
41225 => conv_std_logic_vector(1449, 16),
41226 => conv_std_logic_vector(1610, 16),
41227 => conv_std_logic_vector(1771, 16),
41228 => conv_std_logic_vector(1932, 16),
41229 => conv_std_logic_vector(2093, 16),
41230 => conv_std_logic_vector(2254, 16),
41231 => conv_std_logic_vector(2415, 16),
41232 => conv_std_logic_vector(2576, 16),
41233 => conv_std_logic_vector(2737, 16),
41234 => conv_std_logic_vector(2898, 16),
41235 => conv_std_logic_vector(3059, 16),
41236 => conv_std_logic_vector(3220, 16),
41237 => conv_std_logic_vector(3381, 16),
41238 => conv_std_logic_vector(3542, 16),
41239 => conv_std_logic_vector(3703, 16),
41240 => conv_std_logic_vector(3864, 16),
41241 => conv_std_logic_vector(4025, 16),
41242 => conv_std_logic_vector(4186, 16),
41243 => conv_std_logic_vector(4347, 16),
41244 => conv_std_logic_vector(4508, 16),
41245 => conv_std_logic_vector(4669, 16),
41246 => conv_std_logic_vector(4830, 16),
41247 => conv_std_logic_vector(4991, 16),
41248 => conv_std_logic_vector(5152, 16),
41249 => conv_std_logic_vector(5313, 16),
41250 => conv_std_logic_vector(5474, 16),
41251 => conv_std_logic_vector(5635, 16),
41252 => conv_std_logic_vector(5796, 16),
41253 => conv_std_logic_vector(5957, 16),
41254 => conv_std_logic_vector(6118, 16),
41255 => conv_std_logic_vector(6279, 16),
41256 => conv_std_logic_vector(6440, 16),
41257 => conv_std_logic_vector(6601, 16),
41258 => conv_std_logic_vector(6762, 16),
41259 => conv_std_logic_vector(6923, 16),
41260 => conv_std_logic_vector(7084, 16),
41261 => conv_std_logic_vector(7245, 16),
41262 => conv_std_logic_vector(7406, 16),
41263 => conv_std_logic_vector(7567, 16),
41264 => conv_std_logic_vector(7728, 16),
41265 => conv_std_logic_vector(7889, 16),
41266 => conv_std_logic_vector(8050, 16),
41267 => conv_std_logic_vector(8211, 16),
41268 => conv_std_logic_vector(8372, 16),
41269 => conv_std_logic_vector(8533, 16),
41270 => conv_std_logic_vector(8694, 16),
41271 => conv_std_logic_vector(8855, 16),
41272 => conv_std_logic_vector(9016, 16),
41273 => conv_std_logic_vector(9177, 16),
41274 => conv_std_logic_vector(9338, 16),
41275 => conv_std_logic_vector(9499, 16),
41276 => conv_std_logic_vector(9660, 16),
41277 => conv_std_logic_vector(9821, 16),
41278 => conv_std_logic_vector(9982, 16),
41279 => conv_std_logic_vector(10143, 16),
41280 => conv_std_logic_vector(10304, 16),
41281 => conv_std_logic_vector(10465, 16),
41282 => conv_std_logic_vector(10626, 16),
41283 => conv_std_logic_vector(10787, 16),
41284 => conv_std_logic_vector(10948, 16),
41285 => conv_std_logic_vector(11109, 16),
41286 => conv_std_logic_vector(11270, 16),
41287 => conv_std_logic_vector(11431, 16),
41288 => conv_std_logic_vector(11592, 16),
41289 => conv_std_logic_vector(11753, 16),
41290 => conv_std_logic_vector(11914, 16),
41291 => conv_std_logic_vector(12075, 16),
41292 => conv_std_logic_vector(12236, 16),
41293 => conv_std_logic_vector(12397, 16),
41294 => conv_std_logic_vector(12558, 16),
41295 => conv_std_logic_vector(12719, 16),
41296 => conv_std_logic_vector(12880, 16),
41297 => conv_std_logic_vector(13041, 16),
41298 => conv_std_logic_vector(13202, 16),
41299 => conv_std_logic_vector(13363, 16),
41300 => conv_std_logic_vector(13524, 16),
41301 => conv_std_logic_vector(13685, 16),
41302 => conv_std_logic_vector(13846, 16),
41303 => conv_std_logic_vector(14007, 16),
41304 => conv_std_logic_vector(14168, 16),
41305 => conv_std_logic_vector(14329, 16),
41306 => conv_std_logic_vector(14490, 16),
41307 => conv_std_logic_vector(14651, 16),
41308 => conv_std_logic_vector(14812, 16),
41309 => conv_std_logic_vector(14973, 16),
41310 => conv_std_logic_vector(15134, 16),
41311 => conv_std_logic_vector(15295, 16),
41312 => conv_std_logic_vector(15456, 16),
41313 => conv_std_logic_vector(15617, 16),
41314 => conv_std_logic_vector(15778, 16),
41315 => conv_std_logic_vector(15939, 16),
41316 => conv_std_logic_vector(16100, 16),
41317 => conv_std_logic_vector(16261, 16),
41318 => conv_std_logic_vector(16422, 16),
41319 => conv_std_logic_vector(16583, 16),
41320 => conv_std_logic_vector(16744, 16),
41321 => conv_std_logic_vector(16905, 16),
41322 => conv_std_logic_vector(17066, 16),
41323 => conv_std_logic_vector(17227, 16),
41324 => conv_std_logic_vector(17388, 16),
41325 => conv_std_logic_vector(17549, 16),
41326 => conv_std_logic_vector(17710, 16),
41327 => conv_std_logic_vector(17871, 16),
41328 => conv_std_logic_vector(18032, 16),
41329 => conv_std_logic_vector(18193, 16),
41330 => conv_std_logic_vector(18354, 16),
41331 => conv_std_logic_vector(18515, 16),
41332 => conv_std_logic_vector(18676, 16),
41333 => conv_std_logic_vector(18837, 16),
41334 => conv_std_logic_vector(18998, 16),
41335 => conv_std_logic_vector(19159, 16),
41336 => conv_std_logic_vector(19320, 16),
41337 => conv_std_logic_vector(19481, 16),
41338 => conv_std_logic_vector(19642, 16),
41339 => conv_std_logic_vector(19803, 16),
41340 => conv_std_logic_vector(19964, 16),
41341 => conv_std_logic_vector(20125, 16),
41342 => conv_std_logic_vector(20286, 16),
41343 => conv_std_logic_vector(20447, 16),
41344 => conv_std_logic_vector(20608, 16),
41345 => conv_std_logic_vector(20769, 16),
41346 => conv_std_logic_vector(20930, 16),
41347 => conv_std_logic_vector(21091, 16),
41348 => conv_std_logic_vector(21252, 16),
41349 => conv_std_logic_vector(21413, 16),
41350 => conv_std_logic_vector(21574, 16),
41351 => conv_std_logic_vector(21735, 16),
41352 => conv_std_logic_vector(21896, 16),
41353 => conv_std_logic_vector(22057, 16),
41354 => conv_std_logic_vector(22218, 16),
41355 => conv_std_logic_vector(22379, 16),
41356 => conv_std_logic_vector(22540, 16),
41357 => conv_std_logic_vector(22701, 16),
41358 => conv_std_logic_vector(22862, 16),
41359 => conv_std_logic_vector(23023, 16),
41360 => conv_std_logic_vector(23184, 16),
41361 => conv_std_logic_vector(23345, 16),
41362 => conv_std_logic_vector(23506, 16),
41363 => conv_std_logic_vector(23667, 16),
41364 => conv_std_logic_vector(23828, 16),
41365 => conv_std_logic_vector(23989, 16),
41366 => conv_std_logic_vector(24150, 16),
41367 => conv_std_logic_vector(24311, 16),
41368 => conv_std_logic_vector(24472, 16),
41369 => conv_std_logic_vector(24633, 16),
41370 => conv_std_logic_vector(24794, 16),
41371 => conv_std_logic_vector(24955, 16),
41372 => conv_std_logic_vector(25116, 16),
41373 => conv_std_logic_vector(25277, 16),
41374 => conv_std_logic_vector(25438, 16),
41375 => conv_std_logic_vector(25599, 16),
41376 => conv_std_logic_vector(25760, 16),
41377 => conv_std_logic_vector(25921, 16),
41378 => conv_std_logic_vector(26082, 16),
41379 => conv_std_logic_vector(26243, 16),
41380 => conv_std_logic_vector(26404, 16),
41381 => conv_std_logic_vector(26565, 16),
41382 => conv_std_logic_vector(26726, 16),
41383 => conv_std_logic_vector(26887, 16),
41384 => conv_std_logic_vector(27048, 16),
41385 => conv_std_logic_vector(27209, 16),
41386 => conv_std_logic_vector(27370, 16),
41387 => conv_std_logic_vector(27531, 16),
41388 => conv_std_logic_vector(27692, 16),
41389 => conv_std_logic_vector(27853, 16),
41390 => conv_std_logic_vector(28014, 16),
41391 => conv_std_logic_vector(28175, 16),
41392 => conv_std_logic_vector(28336, 16),
41393 => conv_std_logic_vector(28497, 16),
41394 => conv_std_logic_vector(28658, 16),
41395 => conv_std_logic_vector(28819, 16),
41396 => conv_std_logic_vector(28980, 16),
41397 => conv_std_logic_vector(29141, 16),
41398 => conv_std_logic_vector(29302, 16),
41399 => conv_std_logic_vector(29463, 16),
41400 => conv_std_logic_vector(29624, 16),
41401 => conv_std_logic_vector(29785, 16),
41402 => conv_std_logic_vector(29946, 16),
41403 => conv_std_logic_vector(30107, 16),
41404 => conv_std_logic_vector(30268, 16),
41405 => conv_std_logic_vector(30429, 16),
41406 => conv_std_logic_vector(30590, 16),
41407 => conv_std_logic_vector(30751, 16),
41408 => conv_std_logic_vector(30912, 16),
41409 => conv_std_logic_vector(31073, 16),
41410 => conv_std_logic_vector(31234, 16),
41411 => conv_std_logic_vector(31395, 16),
41412 => conv_std_logic_vector(31556, 16),
41413 => conv_std_logic_vector(31717, 16),
41414 => conv_std_logic_vector(31878, 16),
41415 => conv_std_logic_vector(32039, 16),
41416 => conv_std_logic_vector(32200, 16),
41417 => conv_std_logic_vector(32361, 16),
41418 => conv_std_logic_vector(32522, 16),
41419 => conv_std_logic_vector(32683, 16),
41420 => conv_std_logic_vector(32844, 16),
41421 => conv_std_logic_vector(33005, 16),
41422 => conv_std_logic_vector(33166, 16),
41423 => conv_std_logic_vector(33327, 16),
41424 => conv_std_logic_vector(33488, 16),
41425 => conv_std_logic_vector(33649, 16),
41426 => conv_std_logic_vector(33810, 16),
41427 => conv_std_logic_vector(33971, 16),
41428 => conv_std_logic_vector(34132, 16),
41429 => conv_std_logic_vector(34293, 16),
41430 => conv_std_logic_vector(34454, 16),
41431 => conv_std_logic_vector(34615, 16),
41432 => conv_std_logic_vector(34776, 16),
41433 => conv_std_logic_vector(34937, 16),
41434 => conv_std_logic_vector(35098, 16),
41435 => conv_std_logic_vector(35259, 16),
41436 => conv_std_logic_vector(35420, 16),
41437 => conv_std_logic_vector(35581, 16),
41438 => conv_std_logic_vector(35742, 16),
41439 => conv_std_logic_vector(35903, 16),
41440 => conv_std_logic_vector(36064, 16),
41441 => conv_std_logic_vector(36225, 16),
41442 => conv_std_logic_vector(36386, 16),
41443 => conv_std_logic_vector(36547, 16),
41444 => conv_std_logic_vector(36708, 16),
41445 => conv_std_logic_vector(36869, 16),
41446 => conv_std_logic_vector(37030, 16),
41447 => conv_std_logic_vector(37191, 16),
41448 => conv_std_logic_vector(37352, 16),
41449 => conv_std_logic_vector(37513, 16),
41450 => conv_std_logic_vector(37674, 16),
41451 => conv_std_logic_vector(37835, 16),
41452 => conv_std_logic_vector(37996, 16),
41453 => conv_std_logic_vector(38157, 16),
41454 => conv_std_logic_vector(38318, 16),
41455 => conv_std_logic_vector(38479, 16),
41456 => conv_std_logic_vector(38640, 16),
41457 => conv_std_logic_vector(38801, 16),
41458 => conv_std_logic_vector(38962, 16),
41459 => conv_std_logic_vector(39123, 16),
41460 => conv_std_logic_vector(39284, 16),
41461 => conv_std_logic_vector(39445, 16),
41462 => conv_std_logic_vector(39606, 16),
41463 => conv_std_logic_vector(39767, 16),
41464 => conv_std_logic_vector(39928, 16),
41465 => conv_std_logic_vector(40089, 16),
41466 => conv_std_logic_vector(40250, 16),
41467 => conv_std_logic_vector(40411, 16),
41468 => conv_std_logic_vector(40572, 16),
41469 => conv_std_logic_vector(40733, 16),
41470 => conv_std_logic_vector(40894, 16),
41471 => conv_std_logic_vector(41055, 16),
41472 => conv_std_logic_vector(0, 16),
41473 => conv_std_logic_vector(162, 16),
41474 => conv_std_logic_vector(324, 16),
41475 => conv_std_logic_vector(486, 16),
41476 => conv_std_logic_vector(648, 16),
41477 => conv_std_logic_vector(810, 16),
41478 => conv_std_logic_vector(972, 16),
41479 => conv_std_logic_vector(1134, 16),
41480 => conv_std_logic_vector(1296, 16),
41481 => conv_std_logic_vector(1458, 16),
41482 => conv_std_logic_vector(1620, 16),
41483 => conv_std_logic_vector(1782, 16),
41484 => conv_std_logic_vector(1944, 16),
41485 => conv_std_logic_vector(2106, 16),
41486 => conv_std_logic_vector(2268, 16),
41487 => conv_std_logic_vector(2430, 16),
41488 => conv_std_logic_vector(2592, 16),
41489 => conv_std_logic_vector(2754, 16),
41490 => conv_std_logic_vector(2916, 16),
41491 => conv_std_logic_vector(3078, 16),
41492 => conv_std_logic_vector(3240, 16),
41493 => conv_std_logic_vector(3402, 16),
41494 => conv_std_logic_vector(3564, 16),
41495 => conv_std_logic_vector(3726, 16),
41496 => conv_std_logic_vector(3888, 16),
41497 => conv_std_logic_vector(4050, 16),
41498 => conv_std_logic_vector(4212, 16),
41499 => conv_std_logic_vector(4374, 16),
41500 => conv_std_logic_vector(4536, 16),
41501 => conv_std_logic_vector(4698, 16),
41502 => conv_std_logic_vector(4860, 16),
41503 => conv_std_logic_vector(5022, 16),
41504 => conv_std_logic_vector(5184, 16),
41505 => conv_std_logic_vector(5346, 16),
41506 => conv_std_logic_vector(5508, 16),
41507 => conv_std_logic_vector(5670, 16),
41508 => conv_std_logic_vector(5832, 16),
41509 => conv_std_logic_vector(5994, 16),
41510 => conv_std_logic_vector(6156, 16),
41511 => conv_std_logic_vector(6318, 16),
41512 => conv_std_logic_vector(6480, 16),
41513 => conv_std_logic_vector(6642, 16),
41514 => conv_std_logic_vector(6804, 16),
41515 => conv_std_logic_vector(6966, 16),
41516 => conv_std_logic_vector(7128, 16),
41517 => conv_std_logic_vector(7290, 16),
41518 => conv_std_logic_vector(7452, 16),
41519 => conv_std_logic_vector(7614, 16),
41520 => conv_std_logic_vector(7776, 16),
41521 => conv_std_logic_vector(7938, 16),
41522 => conv_std_logic_vector(8100, 16),
41523 => conv_std_logic_vector(8262, 16),
41524 => conv_std_logic_vector(8424, 16),
41525 => conv_std_logic_vector(8586, 16),
41526 => conv_std_logic_vector(8748, 16),
41527 => conv_std_logic_vector(8910, 16),
41528 => conv_std_logic_vector(9072, 16),
41529 => conv_std_logic_vector(9234, 16),
41530 => conv_std_logic_vector(9396, 16),
41531 => conv_std_logic_vector(9558, 16),
41532 => conv_std_logic_vector(9720, 16),
41533 => conv_std_logic_vector(9882, 16),
41534 => conv_std_logic_vector(10044, 16),
41535 => conv_std_logic_vector(10206, 16),
41536 => conv_std_logic_vector(10368, 16),
41537 => conv_std_logic_vector(10530, 16),
41538 => conv_std_logic_vector(10692, 16),
41539 => conv_std_logic_vector(10854, 16),
41540 => conv_std_logic_vector(11016, 16),
41541 => conv_std_logic_vector(11178, 16),
41542 => conv_std_logic_vector(11340, 16),
41543 => conv_std_logic_vector(11502, 16),
41544 => conv_std_logic_vector(11664, 16),
41545 => conv_std_logic_vector(11826, 16),
41546 => conv_std_logic_vector(11988, 16),
41547 => conv_std_logic_vector(12150, 16),
41548 => conv_std_logic_vector(12312, 16),
41549 => conv_std_logic_vector(12474, 16),
41550 => conv_std_logic_vector(12636, 16),
41551 => conv_std_logic_vector(12798, 16),
41552 => conv_std_logic_vector(12960, 16),
41553 => conv_std_logic_vector(13122, 16),
41554 => conv_std_logic_vector(13284, 16),
41555 => conv_std_logic_vector(13446, 16),
41556 => conv_std_logic_vector(13608, 16),
41557 => conv_std_logic_vector(13770, 16),
41558 => conv_std_logic_vector(13932, 16),
41559 => conv_std_logic_vector(14094, 16),
41560 => conv_std_logic_vector(14256, 16),
41561 => conv_std_logic_vector(14418, 16),
41562 => conv_std_logic_vector(14580, 16),
41563 => conv_std_logic_vector(14742, 16),
41564 => conv_std_logic_vector(14904, 16),
41565 => conv_std_logic_vector(15066, 16),
41566 => conv_std_logic_vector(15228, 16),
41567 => conv_std_logic_vector(15390, 16),
41568 => conv_std_logic_vector(15552, 16),
41569 => conv_std_logic_vector(15714, 16),
41570 => conv_std_logic_vector(15876, 16),
41571 => conv_std_logic_vector(16038, 16),
41572 => conv_std_logic_vector(16200, 16),
41573 => conv_std_logic_vector(16362, 16),
41574 => conv_std_logic_vector(16524, 16),
41575 => conv_std_logic_vector(16686, 16),
41576 => conv_std_logic_vector(16848, 16),
41577 => conv_std_logic_vector(17010, 16),
41578 => conv_std_logic_vector(17172, 16),
41579 => conv_std_logic_vector(17334, 16),
41580 => conv_std_logic_vector(17496, 16),
41581 => conv_std_logic_vector(17658, 16),
41582 => conv_std_logic_vector(17820, 16),
41583 => conv_std_logic_vector(17982, 16),
41584 => conv_std_logic_vector(18144, 16),
41585 => conv_std_logic_vector(18306, 16),
41586 => conv_std_logic_vector(18468, 16),
41587 => conv_std_logic_vector(18630, 16),
41588 => conv_std_logic_vector(18792, 16),
41589 => conv_std_logic_vector(18954, 16),
41590 => conv_std_logic_vector(19116, 16),
41591 => conv_std_logic_vector(19278, 16),
41592 => conv_std_logic_vector(19440, 16),
41593 => conv_std_logic_vector(19602, 16),
41594 => conv_std_logic_vector(19764, 16),
41595 => conv_std_logic_vector(19926, 16),
41596 => conv_std_logic_vector(20088, 16),
41597 => conv_std_logic_vector(20250, 16),
41598 => conv_std_logic_vector(20412, 16),
41599 => conv_std_logic_vector(20574, 16),
41600 => conv_std_logic_vector(20736, 16),
41601 => conv_std_logic_vector(20898, 16),
41602 => conv_std_logic_vector(21060, 16),
41603 => conv_std_logic_vector(21222, 16),
41604 => conv_std_logic_vector(21384, 16),
41605 => conv_std_logic_vector(21546, 16),
41606 => conv_std_logic_vector(21708, 16),
41607 => conv_std_logic_vector(21870, 16),
41608 => conv_std_logic_vector(22032, 16),
41609 => conv_std_logic_vector(22194, 16),
41610 => conv_std_logic_vector(22356, 16),
41611 => conv_std_logic_vector(22518, 16),
41612 => conv_std_logic_vector(22680, 16),
41613 => conv_std_logic_vector(22842, 16),
41614 => conv_std_logic_vector(23004, 16),
41615 => conv_std_logic_vector(23166, 16),
41616 => conv_std_logic_vector(23328, 16),
41617 => conv_std_logic_vector(23490, 16),
41618 => conv_std_logic_vector(23652, 16),
41619 => conv_std_logic_vector(23814, 16),
41620 => conv_std_logic_vector(23976, 16),
41621 => conv_std_logic_vector(24138, 16),
41622 => conv_std_logic_vector(24300, 16),
41623 => conv_std_logic_vector(24462, 16),
41624 => conv_std_logic_vector(24624, 16),
41625 => conv_std_logic_vector(24786, 16),
41626 => conv_std_logic_vector(24948, 16),
41627 => conv_std_logic_vector(25110, 16),
41628 => conv_std_logic_vector(25272, 16),
41629 => conv_std_logic_vector(25434, 16),
41630 => conv_std_logic_vector(25596, 16),
41631 => conv_std_logic_vector(25758, 16),
41632 => conv_std_logic_vector(25920, 16),
41633 => conv_std_logic_vector(26082, 16),
41634 => conv_std_logic_vector(26244, 16),
41635 => conv_std_logic_vector(26406, 16),
41636 => conv_std_logic_vector(26568, 16),
41637 => conv_std_logic_vector(26730, 16),
41638 => conv_std_logic_vector(26892, 16),
41639 => conv_std_logic_vector(27054, 16),
41640 => conv_std_logic_vector(27216, 16),
41641 => conv_std_logic_vector(27378, 16),
41642 => conv_std_logic_vector(27540, 16),
41643 => conv_std_logic_vector(27702, 16),
41644 => conv_std_logic_vector(27864, 16),
41645 => conv_std_logic_vector(28026, 16),
41646 => conv_std_logic_vector(28188, 16),
41647 => conv_std_logic_vector(28350, 16),
41648 => conv_std_logic_vector(28512, 16),
41649 => conv_std_logic_vector(28674, 16),
41650 => conv_std_logic_vector(28836, 16),
41651 => conv_std_logic_vector(28998, 16),
41652 => conv_std_logic_vector(29160, 16),
41653 => conv_std_logic_vector(29322, 16),
41654 => conv_std_logic_vector(29484, 16),
41655 => conv_std_logic_vector(29646, 16),
41656 => conv_std_logic_vector(29808, 16),
41657 => conv_std_logic_vector(29970, 16),
41658 => conv_std_logic_vector(30132, 16),
41659 => conv_std_logic_vector(30294, 16),
41660 => conv_std_logic_vector(30456, 16),
41661 => conv_std_logic_vector(30618, 16),
41662 => conv_std_logic_vector(30780, 16),
41663 => conv_std_logic_vector(30942, 16),
41664 => conv_std_logic_vector(31104, 16),
41665 => conv_std_logic_vector(31266, 16),
41666 => conv_std_logic_vector(31428, 16),
41667 => conv_std_logic_vector(31590, 16),
41668 => conv_std_logic_vector(31752, 16),
41669 => conv_std_logic_vector(31914, 16),
41670 => conv_std_logic_vector(32076, 16),
41671 => conv_std_logic_vector(32238, 16),
41672 => conv_std_logic_vector(32400, 16),
41673 => conv_std_logic_vector(32562, 16),
41674 => conv_std_logic_vector(32724, 16),
41675 => conv_std_logic_vector(32886, 16),
41676 => conv_std_logic_vector(33048, 16),
41677 => conv_std_logic_vector(33210, 16),
41678 => conv_std_logic_vector(33372, 16),
41679 => conv_std_logic_vector(33534, 16),
41680 => conv_std_logic_vector(33696, 16),
41681 => conv_std_logic_vector(33858, 16),
41682 => conv_std_logic_vector(34020, 16),
41683 => conv_std_logic_vector(34182, 16),
41684 => conv_std_logic_vector(34344, 16),
41685 => conv_std_logic_vector(34506, 16),
41686 => conv_std_logic_vector(34668, 16),
41687 => conv_std_logic_vector(34830, 16),
41688 => conv_std_logic_vector(34992, 16),
41689 => conv_std_logic_vector(35154, 16),
41690 => conv_std_logic_vector(35316, 16),
41691 => conv_std_logic_vector(35478, 16),
41692 => conv_std_logic_vector(35640, 16),
41693 => conv_std_logic_vector(35802, 16),
41694 => conv_std_logic_vector(35964, 16),
41695 => conv_std_logic_vector(36126, 16),
41696 => conv_std_logic_vector(36288, 16),
41697 => conv_std_logic_vector(36450, 16),
41698 => conv_std_logic_vector(36612, 16),
41699 => conv_std_logic_vector(36774, 16),
41700 => conv_std_logic_vector(36936, 16),
41701 => conv_std_logic_vector(37098, 16),
41702 => conv_std_logic_vector(37260, 16),
41703 => conv_std_logic_vector(37422, 16),
41704 => conv_std_logic_vector(37584, 16),
41705 => conv_std_logic_vector(37746, 16),
41706 => conv_std_logic_vector(37908, 16),
41707 => conv_std_logic_vector(38070, 16),
41708 => conv_std_logic_vector(38232, 16),
41709 => conv_std_logic_vector(38394, 16),
41710 => conv_std_logic_vector(38556, 16),
41711 => conv_std_logic_vector(38718, 16),
41712 => conv_std_logic_vector(38880, 16),
41713 => conv_std_logic_vector(39042, 16),
41714 => conv_std_logic_vector(39204, 16),
41715 => conv_std_logic_vector(39366, 16),
41716 => conv_std_logic_vector(39528, 16),
41717 => conv_std_logic_vector(39690, 16),
41718 => conv_std_logic_vector(39852, 16),
41719 => conv_std_logic_vector(40014, 16),
41720 => conv_std_logic_vector(40176, 16),
41721 => conv_std_logic_vector(40338, 16),
41722 => conv_std_logic_vector(40500, 16),
41723 => conv_std_logic_vector(40662, 16),
41724 => conv_std_logic_vector(40824, 16),
41725 => conv_std_logic_vector(40986, 16),
41726 => conv_std_logic_vector(41148, 16),
41727 => conv_std_logic_vector(41310, 16),
41728 => conv_std_logic_vector(0, 16),
41729 => conv_std_logic_vector(163, 16),
41730 => conv_std_logic_vector(326, 16),
41731 => conv_std_logic_vector(489, 16),
41732 => conv_std_logic_vector(652, 16),
41733 => conv_std_logic_vector(815, 16),
41734 => conv_std_logic_vector(978, 16),
41735 => conv_std_logic_vector(1141, 16),
41736 => conv_std_logic_vector(1304, 16),
41737 => conv_std_logic_vector(1467, 16),
41738 => conv_std_logic_vector(1630, 16),
41739 => conv_std_logic_vector(1793, 16),
41740 => conv_std_logic_vector(1956, 16),
41741 => conv_std_logic_vector(2119, 16),
41742 => conv_std_logic_vector(2282, 16),
41743 => conv_std_logic_vector(2445, 16),
41744 => conv_std_logic_vector(2608, 16),
41745 => conv_std_logic_vector(2771, 16),
41746 => conv_std_logic_vector(2934, 16),
41747 => conv_std_logic_vector(3097, 16),
41748 => conv_std_logic_vector(3260, 16),
41749 => conv_std_logic_vector(3423, 16),
41750 => conv_std_logic_vector(3586, 16),
41751 => conv_std_logic_vector(3749, 16),
41752 => conv_std_logic_vector(3912, 16),
41753 => conv_std_logic_vector(4075, 16),
41754 => conv_std_logic_vector(4238, 16),
41755 => conv_std_logic_vector(4401, 16),
41756 => conv_std_logic_vector(4564, 16),
41757 => conv_std_logic_vector(4727, 16),
41758 => conv_std_logic_vector(4890, 16),
41759 => conv_std_logic_vector(5053, 16),
41760 => conv_std_logic_vector(5216, 16),
41761 => conv_std_logic_vector(5379, 16),
41762 => conv_std_logic_vector(5542, 16),
41763 => conv_std_logic_vector(5705, 16),
41764 => conv_std_logic_vector(5868, 16),
41765 => conv_std_logic_vector(6031, 16),
41766 => conv_std_logic_vector(6194, 16),
41767 => conv_std_logic_vector(6357, 16),
41768 => conv_std_logic_vector(6520, 16),
41769 => conv_std_logic_vector(6683, 16),
41770 => conv_std_logic_vector(6846, 16),
41771 => conv_std_logic_vector(7009, 16),
41772 => conv_std_logic_vector(7172, 16),
41773 => conv_std_logic_vector(7335, 16),
41774 => conv_std_logic_vector(7498, 16),
41775 => conv_std_logic_vector(7661, 16),
41776 => conv_std_logic_vector(7824, 16),
41777 => conv_std_logic_vector(7987, 16),
41778 => conv_std_logic_vector(8150, 16),
41779 => conv_std_logic_vector(8313, 16),
41780 => conv_std_logic_vector(8476, 16),
41781 => conv_std_logic_vector(8639, 16),
41782 => conv_std_logic_vector(8802, 16),
41783 => conv_std_logic_vector(8965, 16),
41784 => conv_std_logic_vector(9128, 16),
41785 => conv_std_logic_vector(9291, 16),
41786 => conv_std_logic_vector(9454, 16),
41787 => conv_std_logic_vector(9617, 16),
41788 => conv_std_logic_vector(9780, 16),
41789 => conv_std_logic_vector(9943, 16),
41790 => conv_std_logic_vector(10106, 16),
41791 => conv_std_logic_vector(10269, 16),
41792 => conv_std_logic_vector(10432, 16),
41793 => conv_std_logic_vector(10595, 16),
41794 => conv_std_logic_vector(10758, 16),
41795 => conv_std_logic_vector(10921, 16),
41796 => conv_std_logic_vector(11084, 16),
41797 => conv_std_logic_vector(11247, 16),
41798 => conv_std_logic_vector(11410, 16),
41799 => conv_std_logic_vector(11573, 16),
41800 => conv_std_logic_vector(11736, 16),
41801 => conv_std_logic_vector(11899, 16),
41802 => conv_std_logic_vector(12062, 16),
41803 => conv_std_logic_vector(12225, 16),
41804 => conv_std_logic_vector(12388, 16),
41805 => conv_std_logic_vector(12551, 16),
41806 => conv_std_logic_vector(12714, 16),
41807 => conv_std_logic_vector(12877, 16),
41808 => conv_std_logic_vector(13040, 16),
41809 => conv_std_logic_vector(13203, 16),
41810 => conv_std_logic_vector(13366, 16),
41811 => conv_std_logic_vector(13529, 16),
41812 => conv_std_logic_vector(13692, 16),
41813 => conv_std_logic_vector(13855, 16),
41814 => conv_std_logic_vector(14018, 16),
41815 => conv_std_logic_vector(14181, 16),
41816 => conv_std_logic_vector(14344, 16),
41817 => conv_std_logic_vector(14507, 16),
41818 => conv_std_logic_vector(14670, 16),
41819 => conv_std_logic_vector(14833, 16),
41820 => conv_std_logic_vector(14996, 16),
41821 => conv_std_logic_vector(15159, 16),
41822 => conv_std_logic_vector(15322, 16),
41823 => conv_std_logic_vector(15485, 16),
41824 => conv_std_logic_vector(15648, 16),
41825 => conv_std_logic_vector(15811, 16),
41826 => conv_std_logic_vector(15974, 16),
41827 => conv_std_logic_vector(16137, 16),
41828 => conv_std_logic_vector(16300, 16),
41829 => conv_std_logic_vector(16463, 16),
41830 => conv_std_logic_vector(16626, 16),
41831 => conv_std_logic_vector(16789, 16),
41832 => conv_std_logic_vector(16952, 16),
41833 => conv_std_logic_vector(17115, 16),
41834 => conv_std_logic_vector(17278, 16),
41835 => conv_std_logic_vector(17441, 16),
41836 => conv_std_logic_vector(17604, 16),
41837 => conv_std_logic_vector(17767, 16),
41838 => conv_std_logic_vector(17930, 16),
41839 => conv_std_logic_vector(18093, 16),
41840 => conv_std_logic_vector(18256, 16),
41841 => conv_std_logic_vector(18419, 16),
41842 => conv_std_logic_vector(18582, 16),
41843 => conv_std_logic_vector(18745, 16),
41844 => conv_std_logic_vector(18908, 16),
41845 => conv_std_logic_vector(19071, 16),
41846 => conv_std_logic_vector(19234, 16),
41847 => conv_std_logic_vector(19397, 16),
41848 => conv_std_logic_vector(19560, 16),
41849 => conv_std_logic_vector(19723, 16),
41850 => conv_std_logic_vector(19886, 16),
41851 => conv_std_logic_vector(20049, 16),
41852 => conv_std_logic_vector(20212, 16),
41853 => conv_std_logic_vector(20375, 16),
41854 => conv_std_logic_vector(20538, 16),
41855 => conv_std_logic_vector(20701, 16),
41856 => conv_std_logic_vector(20864, 16),
41857 => conv_std_logic_vector(21027, 16),
41858 => conv_std_logic_vector(21190, 16),
41859 => conv_std_logic_vector(21353, 16),
41860 => conv_std_logic_vector(21516, 16),
41861 => conv_std_logic_vector(21679, 16),
41862 => conv_std_logic_vector(21842, 16),
41863 => conv_std_logic_vector(22005, 16),
41864 => conv_std_logic_vector(22168, 16),
41865 => conv_std_logic_vector(22331, 16),
41866 => conv_std_logic_vector(22494, 16),
41867 => conv_std_logic_vector(22657, 16),
41868 => conv_std_logic_vector(22820, 16),
41869 => conv_std_logic_vector(22983, 16),
41870 => conv_std_logic_vector(23146, 16),
41871 => conv_std_logic_vector(23309, 16),
41872 => conv_std_logic_vector(23472, 16),
41873 => conv_std_logic_vector(23635, 16),
41874 => conv_std_logic_vector(23798, 16),
41875 => conv_std_logic_vector(23961, 16),
41876 => conv_std_logic_vector(24124, 16),
41877 => conv_std_logic_vector(24287, 16),
41878 => conv_std_logic_vector(24450, 16),
41879 => conv_std_logic_vector(24613, 16),
41880 => conv_std_logic_vector(24776, 16),
41881 => conv_std_logic_vector(24939, 16),
41882 => conv_std_logic_vector(25102, 16),
41883 => conv_std_logic_vector(25265, 16),
41884 => conv_std_logic_vector(25428, 16),
41885 => conv_std_logic_vector(25591, 16),
41886 => conv_std_logic_vector(25754, 16),
41887 => conv_std_logic_vector(25917, 16),
41888 => conv_std_logic_vector(26080, 16),
41889 => conv_std_logic_vector(26243, 16),
41890 => conv_std_logic_vector(26406, 16),
41891 => conv_std_logic_vector(26569, 16),
41892 => conv_std_logic_vector(26732, 16),
41893 => conv_std_logic_vector(26895, 16),
41894 => conv_std_logic_vector(27058, 16),
41895 => conv_std_logic_vector(27221, 16),
41896 => conv_std_logic_vector(27384, 16),
41897 => conv_std_logic_vector(27547, 16),
41898 => conv_std_logic_vector(27710, 16),
41899 => conv_std_logic_vector(27873, 16),
41900 => conv_std_logic_vector(28036, 16),
41901 => conv_std_logic_vector(28199, 16),
41902 => conv_std_logic_vector(28362, 16),
41903 => conv_std_logic_vector(28525, 16),
41904 => conv_std_logic_vector(28688, 16),
41905 => conv_std_logic_vector(28851, 16),
41906 => conv_std_logic_vector(29014, 16),
41907 => conv_std_logic_vector(29177, 16),
41908 => conv_std_logic_vector(29340, 16),
41909 => conv_std_logic_vector(29503, 16),
41910 => conv_std_logic_vector(29666, 16),
41911 => conv_std_logic_vector(29829, 16),
41912 => conv_std_logic_vector(29992, 16),
41913 => conv_std_logic_vector(30155, 16),
41914 => conv_std_logic_vector(30318, 16),
41915 => conv_std_logic_vector(30481, 16),
41916 => conv_std_logic_vector(30644, 16),
41917 => conv_std_logic_vector(30807, 16),
41918 => conv_std_logic_vector(30970, 16),
41919 => conv_std_logic_vector(31133, 16),
41920 => conv_std_logic_vector(31296, 16),
41921 => conv_std_logic_vector(31459, 16),
41922 => conv_std_logic_vector(31622, 16),
41923 => conv_std_logic_vector(31785, 16),
41924 => conv_std_logic_vector(31948, 16),
41925 => conv_std_logic_vector(32111, 16),
41926 => conv_std_logic_vector(32274, 16),
41927 => conv_std_logic_vector(32437, 16),
41928 => conv_std_logic_vector(32600, 16),
41929 => conv_std_logic_vector(32763, 16),
41930 => conv_std_logic_vector(32926, 16),
41931 => conv_std_logic_vector(33089, 16),
41932 => conv_std_logic_vector(33252, 16),
41933 => conv_std_logic_vector(33415, 16),
41934 => conv_std_logic_vector(33578, 16),
41935 => conv_std_logic_vector(33741, 16),
41936 => conv_std_logic_vector(33904, 16),
41937 => conv_std_logic_vector(34067, 16),
41938 => conv_std_logic_vector(34230, 16),
41939 => conv_std_logic_vector(34393, 16),
41940 => conv_std_logic_vector(34556, 16),
41941 => conv_std_logic_vector(34719, 16),
41942 => conv_std_logic_vector(34882, 16),
41943 => conv_std_logic_vector(35045, 16),
41944 => conv_std_logic_vector(35208, 16),
41945 => conv_std_logic_vector(35371, 16),
41946 => conv_std_logic_vector(35534, 16),
41947 => conv_std_logic_vector(35697, 16),
41948 => conv_std_logic_vector(35860, 16),
41949 => conv_std_logic_vector(36023, 16),
41950 => conv_std_logic_vector(36186, 16),
41951 => conv_std_logic_vector(36349, 16),
41952 => conv_std_logic_vector(36512, 16),
41953 => conv_std_logic_vector(36675, 16),
41954 => conv_std_logic_vector(36838, 16),
41955 => conv_std_logic_vector(37001, 16),
41956 => conv_std_logic_vector(37164, 16),
41957 => conv_std_logic_vector(37327, 16),
41958 => conv_std_logic_vector(37490, 16),
41959 => conv_std_logic_vector(37653, 16),
41960 => conv_std_logic_vector(37816, 16),
41961 => conv_std_logic_vector(37979, 16),
41962 => conv_std_logic_vector(38142, 16),
41963 => conv_std_logic_vector(38305, 16),
41964 => conv_std_logic_vector(38468, 16),
41965 => conv_std_logic_vector(38631, 16),
41966 => conv_std_logic_vector(38794, 16),
41967 => conv_std_logic_vector(38957, 16),
41968 => conv_std_logic_vector(39120, 16),
41969 => conv_std_logic_vector(39283, 16),
41970 => conv_std_logic_vector(39446, 16),
41971 => conv_std_logic_vector(39609, 16),
41972 => conv_std_logic_vector(39772, 16),
41973 => conv_std_logic_vector(39935, 16),
41974 => conv_std_logic_vector(40098, 16),
41975 => conv_std_logic_vector(40261, 16),
41976 => conv_std_logic_vector(40424, 16),
41977 => conv_std_logic_vector(40587, 16),
41978 => conv_std_logic_vector(40750, 16),
41979 => conv_std_logic_vector(40913, 16),
41980 => conv_std_logic_vector(41076, 16),
41981 => conv_std_logic_vector(41239, 16),
41982 => conv_std_logic_vector(41402, 16),
41983 => conv_std_logic_vector(41565, 16),
41984 => conv_std_logic_vector(0, 16),
41985 => conv_std_logic_vector(164, 16),
41986 => conv_std_logic_vector(328, 16),
41987 => conv_std_logic_vector(492, 16),
41988 => conv_std_logic_vector(656, 16),
41989 => conv_std_logic_vector(820, 16),
41990 => conv_std_logic_vector(984, 16),
41991 => conv_std_logic_vector(1148, 16),
41992 => conv_std_logic_vector(1312, 16),
41993 => conv_std_logic_vector(1476, 16),
41994 => conv_std_logic_vector(1640, 16),
41995 => conv_std_logic_vector(1804, 16),
41996 => conv_std_logic_vector(1968, 16),
41997 => conv_std_logic_vector(2132, 16),
41998 => conv_std_logic_vector(2296, 16),
41999 => conv_std_logic_vector(2460, 16),
42000 => conv_std_logic_vector(2624, 16),
42001 => conv_std_logic_vector(2788, 16),
42002 => conv_std_logic_vector(2952, 16),
42003 => conv_std_logic_vector(3116, 16),
42004 => conv_std_logic_vector(3280, 16),
42005 => conv_std_logic_vector(3444, 16),
42006 => conv_std_logic_vector(3608, 16),
42007 => conv_std_logic_vector(3772, 16),
42008 => conv_std_logic_vector(3936, 16),
42009 => conv_std_logic_vector(4100, 16),
42010 => conv_std_logic_vector(4264, 16),
42011 => conv_std_logic_vector(4428, 16),
42012 => conv_std_logic_vector(4592, 16),
42013 => conv_std_logic_vector(4756, 16),
42014 => conv_std_logic_vector(4920, 16),
42015 => conv_std_logic_vector(5084, 16),
42016 => conv_std_logic_vector(5248, 16),
42017 => conv_std_logic_vector(5412, 16),
42018 => conv_std_logic_vector(5576, 16),
42019 => conv_std_logic_vector(5740, 16),
42020 => conv_std_logic_vector(5904, 16),
42021 => conv_std_logic_vector(6068, 16),
42022 => conv_std_logic_vector(6232, 16),
42023 => conv_std_logic_vector(6396, 16),
42024 => conv_std_logic_vector(6560, 16),
42025 => conv_std_logic_vector(6724, 16),
42026 => conv_std_logic_vector(6888, 16),
42027 => conv_std_logic_vector(7052, 16),
42028 => conv_std_logic_vector(7216, 16),
42029 => conv_std_logic_vector(7380, 16),
42030 => conv_std_logic_vector(7544, 16),
42031 => conv_std_logic_vector(7708, 16),
42032 => conv_std_logic_vector(7872, 16),
42033 => conv_std_logic_vector(8036, 16),
42034 => conv_std_logic_vector(8200, 16),
42035 => conv_std_logic_vector(8364, 16),
42036 => conv_std_logic_vector(8528, 16),
42037 => conv_std_logic_vector(8692, 16),
42038 => conv_std_logic_vector(8856, 16),
42039 => conv_std_logic_vector(9020, 16),
42040 => conv_std_logic_vector(9184, 16),
42041 => conv_std_logic_vector(9348, 16),
42042 => conv_std_logic_vector(9512, 16),
42043 => conv_std_logic_vector(9676, 16),
42044 => conv_std_logic_vector(9840, 16),
42045 => conv_std_logic_vector(10004, 16),
42046 => conv_std_logic_vector(10168, 16),
42047 => conv_std_logic_vector(10332, 16),
42048 => conv_std_logic_vector(10496, 16),
42049 => conv_std_logic_vector(10660, 16),
42050 => conv_std_logic_vector(10824, 16),
42051 => conv_std_logic_vector(10988, 16),
42052 => conv_std_logic_vector(11152, 16),
42053 => conv_std_logic_vector(11316, 16),
42054 => conv_std_logic_vector(11480, 16),
42055 => conv_std_logic_vector(11644, 16),
42056 => conv_std_logic_vector(11808, 16),
42057 => conv_std_logic_vector(11972, 16),
42058 => conv_std_logic_vector(12136, 16),
42059 => conv_std_logic_vector(12300, 16),
42060 => conv_std_logic_vector(12464, 16),
42061 => conv_std_logic_vector(12628, 16),
42062 => conv_std_logic_vector(12792, 16),
42063 => conv_std_logic_vector(12956, 16),
42064 => conv_std_logic_vector(13120, 16),
42065 => conv_std_logic_vector(13284, 16),
42066 => conv_std_logic_vector(13448, 16),
42067 => conv_std_logic_vector(13612, 16),
42068 => conv_std_logic_vector(13776, 16),
42069 => conv_std_logic_vector(13940, 16),
42070 => conv_std_logic_vector(14104, 16),
42071 => conv_std_logic_vector(14268, 16),
42072 => conv_std_logic_vector(14432, 16),
42073 => conv_std_logic_vector(14596, 16),
42074 => conv_std_logic_vector(14760, 16),
42075 => conv_std_logic_vector(14924, 16),
42076 => conv_std_logic_vector(15088, 16),
42077 => conv_std_logic_vector(15252, 16),
42078 => conv_std_logic_vector(15416, 16),
42079 => conv_std_logic_vector(15580, 16),
42080 => conv_std_logic_vector(15744, 16),
42081 => conv_std_logic_vector(15908, 16),
42082 => conv_std_logic_vector(16072, 16),
42083 => conv_std_logic_vector(16236, 16),
42084 => conv_std_logic_vector(16400, 16),
42085 => conv_std_logic_vector(16564, 16),
42086 => conv_std_logic_vector(16728, 16),
42087 => conv_std_logic_vector(16892, 16),
42088 => conv_std_logic_vector(17056, 16),
42089 => conv_std_logic_vector(17220, 16),
42090 => conv_std_logic_vector(17384, 16),
42091 => conv_std_logic_vector(17548, 16),
42092 => conv_std_logic_vector(17712, 16),
42093 => conv_std_logic_vector(17876, 16),
42094 => conv_std_logic_vector(18040, 16),
42095 => conv_std_logic_vector(18204, 16),
42096 => conv_std_logic_vector(18368, 16),
42097 => conv_std_logic_vector(18532, 16),
42098 => conv_std_logic_vector(18696, 16),
42099 => conv_std_logic_vector(18860, 16),
42100 => conv_std_logic_vector(19024, 16),
42101 => conv_std_logic_vector(19188, 16),
42102 => conv_std_logic_vector(19352, 16),
42103 => conv_std_logic_vector(19516, 16),
42104 => conv_std_logic_vector(19680, 16),
42105 => conv_std_logic_vector(19844, 16),
42106 => conv_std_logic_vector(20008, 16),
42107 => conv_std_logic_vector(20172, 16),
42108 => conv_std_logic_vector(20336, 16),
42109 => conv_std_logic_vector(20500, 16),
42110 => conv_std_logic_vector(20664, 16),
42111 => conv_std_logic_vector(20828, 16),
42112 => conv_std_logic_vector(20992, 16),
42113 => conv_std_logic_vector(21156, 16),
42114 => conv_std_logic_vector(21320, 16),
42115 => conv_std_logic_vector(21484, 16),
42116 => conv_std_logic_vector(21648, 16),
42117 => conv_std_logic_vector(21812, 16),
42118 => conv_std_logic_vector(21976, 16),
42119 => conv_std_logic_vector(22140, 16),
42120 => conv_std_logic_vector(22304, 16),
42121 => conv_std_logic_vector(22468, 16),
42122 => conv_std_logic_vector(22632, 16),
42123 => conv_std_logic_vector(22796, 16),
42124 => conv_std_logic_vector(22960, 16),
42125 => conv_std_logic_vector(23124, 16),
42126 => conv_std_logic_vector(23288, 16),
42127 => conv_std_logic_vector(23452, 16),
42128 => conv_std_logic_vector(23616, 16),
42129 => conv_std_logic_vector(23780, 16),
42130 => conv_std_logic_vector(23944, 16),
42131 => conv_std_logic_vector(24108, 16),
42132 => conv_std_logic_vector(24272, 16),
42133 => conv_std_logic_vector(24436, 16),
42134 => conv_std_logic_vector(24600, 16),
42135 => conv_std_logic_vector(24764, 16),
42136 => conv_std_logic_vector(24928, 16),
42137 => conv_std_logic_vector(25092, 16),
42138 => conv_std_logic_vector(25256, 16),
42139 => conv_std_logic_vector(25420, 16),
42140 => conv_std_logic_vector(25584, 16),
42141 => conv_std_logic_vector(25748, 16),
42142 => conv_std_logic_vector(25912, 16),
42143 => conv_std_logic_vector(26076, 16),
42144 => conv_std_logic_vector(26240, 16),
42145 => conv_std_logic_vector(26404, 16),
42146 => conv_std_logic_vector(26568, 16),
42147 => conv_std_logic_vector(26732, 16),
42148 => conv_std_logic_vector(26896, 16),
42149 => conv_std_logic_vector(27060, 16),
42150 => conv_std_logic_vector(27224, 16),
42151 => conv_std_logic_vector(27388, 16),
42152 => conv_std_logic_vector(27552, 16),
42153 => conv_std_logic_vector(27716, 16),
42154 => conv_std_logic_vector(27880, 16),
42155 => conv_std_logic_vector(28044, 16),
42156 => conv_std_logic_vector(28208, 16),
42157 => conv_std_logic_vector(28372, 16),
42158 => conv_std_logic_vector(28536, 16),
42159 => conv_std_logic_vector(28700, 16),
42160 => conv_std_logic_vector(28864, 16),
42161 => conv_std_logic_vector(29028, 16),
42162 => conv_std_logic_vector(29192, 16),
42163 => conv_std_logic_vector(29356, 16),
42164 => conv_std_logic_vector(29520, 16),
42165 => conv_std_logic_vector(29684, 16),
42166 => conv_std_logic_vector(29848, 16),
42167 => conv_std_logic_vector(30012, 16),
42168 => conv_std_logic_vector(30176, 16),
42169 => conv_std_logic_vector(30340, 16),
42170 => conv_std_logic_vector(30504, 16),
42171 => conv_std_logic_vector(30668, 16),
42172 => conv_std_logic_vector(30832, 16),
42173 => conv_std_logic_vector(30996, 16),
42174 => conv_std_logic_vector(31160, 16),
42175 => conv_std_logic_vector(31324, 16),
42176 => conv_std_logic_vector(31488, 16),
42177 => conv_std_logic_vector(31652, 16),
42178 => conv_std_logic_vector(31816, 16),
42179 => conv_std_logic_vector(31980, 16),
42180 => conv_std_logic_vector(32144, 16),
42181 => conv_std_logic_vector(32308, 16),
42182 => conv_std_logic_vector(32472, 16),
42183 => conv_std_logic_vector(32636, 16),
42184 => conv_std_logic_vector(32800, 16),
42185 => conv_std_logic_vector(32964, 16),
42186 => conv_std_logic_vector(33128, 16),
42187 => conv_std_logic_vector(33292, 16),
42188 => conv_std_logic_vector(33456, 16),
42189 => conv_std_logic_vector(33620, 16),
42190 => conv_std_logic_vector(33784, 16),
42191 => conv_std_logic_vector(33948, 16),
42192 => conv_std_logic_vector(34112, 16),
42193 => conv_std_logic_vector(34276, 16),
42194 => conv_std_logic_vector(34440, 16),
42195 => conv_std_logic_vector(34604, 16),
42196 => conv_std_logic_vector(34768, 16),
42197 => conv_std_logic_vector(34932, 16),
42198 => conv_std_logic_vector(35096, 16),
42199 => conv_std_logic_vector(35260, 16),
42200 => conv_std_logic_vector(35424, 16),
42201 => conv_std_logic_vector(35588, 16),
42202 => conv_std_logic_vector(35752, 16),
42203 => conv_std_logic_vector(35916, 16),
42204 => conv_std_logic_vector(36080, 16),
42205 => conv_std_logic_vector(36244, 16),
42206 => conv_std_logic_vector(36408, 16),
42207 => conv_std_logic_vector(36572, 16),
42208 => conv_std_logic_vector(36736, 16),
42209 => conv_std_logic_vector(36900, 16),
42210 => conv_std_logic_vector(37064, 16),
42211 => conv_std_logic_vector(37228, 16),
42212 => conv_std_logic_vector(37392, 16),
42213 => conv_std_logic_vector(37556, 16),
42214 => conv_std_logic_vector(37720, 16),
42215 => conv_std_logic_vector(37884, 16),
42216 => conv_std_logic_vector(38048, 16),
42217 => conv_std_logic_vector(38212, 16),
42218 => conv_std_logic_vector(38376, 16),
42219 => conv_std_logic_vector(38540, 16),
42220 => conv_std_logic_vector(38704, 16),
42221 => conv_std_logic_vector(38868, 16),
42222 => conv_std_logic_vector(39032, 16),
42223 => conv_std_logic_vector(39196, 16),
42224 => conv_std_logic_vector(39360, 16),
42225 => conv_std_logic_vector(39524, 16),
42226 => conv_std_logic_vector(39688, 16),
42227 => conv_std_logic_vector(39852, 16),
42228 => conv_std_logic_vector(40016, 16),
42229 => conv_std_logic_vector(40180, 16),
42230 => conv_std_logic_vector(40344, 16),
42231 => conv_std_logic_vector(40508, 16),
42232 => conv_std_logic_vector(40672, 16),
42233 => conv_std_logic_vector(40836, 16),
42234 => conv_std_logic_vector(41000, 16),
42235 => conv_std_logic_vector(41164, 16),
42236 => conv_std_logic_vector(41328, 16),
42237 => conv_std_logic_vector(41492, 16),
42238 => conv_std_logic_vector(41656, 16),
42239 => conv_std_logic_vector(41820, 16),
42240 => conv_std_logic_vector(0, 16),
42241 => conv_std_logic_vector(165, 16),
42242 => conv_std_logic_vector(330, 16),
42243 => conv_std_logic_vector(495, 16),
42244 => conv_std_logic_vector(660, 16),
42245 => conv_std_logic_vector(825, 16),
42246 => conv_std_logic_vector(990, 16),
42247 => conv_std_logic_vector(1155, 16),
42248 => conv_std_logic_vector(1320, 16),
42249 => conv_std_logic_vector(1485, 16),
42250 => conv_std_logic_vector(1650, 16),
42251 => conv_std_logic_vector(1815, 16),
42252 => conv_std_logic_vector(1980, 16),
42253 => conv_std_logic_vector(2145, 16),
42254 => conv_std_logic_vector(2310, 16),
42255 => conv_std_logic_vector(2475, 16),
42256 => conv_std_logic_vector(2640, 16),
42257 => conv_std_logic_vector(2805, 16),
42258 => conv_std_logic_vector(2970, 16),
42259 => conv_std_logic_vector(3135, 16),
42260 => conv_std_logic_vector(3300, 16),
42261 => conv_std_logic_vector(3465, 16),
42262 => conv_std_logic_vector(3630, 16),
42263 => conv_std_logic_vector(3795, 16),
42264 => conv_std_logic_vector(3960, 16),
42265 => conv_std_logic_vector(4125, 16),
42266 => conv_std_logic_vector(4290, 16),
42267 => conv_std_logic_vector(4455, 16),
42268 => conv_std_logic_vector(4620, 16),
42269 => conv_std_logic_vector(4785, 16),
42270 => conv_std_logic_vector(4950, 16),
42271 => conv_std_logic_vector(5115, 16),
42272 => conv_std_logic_vector(5280, 16),
42273 => conv_std_logic_vector(5445, 16),
42274 => conv_std_logic_vector(5610, 16),
42275 => conv_std_logic_vector(5775, 16),
42276 => conv_std_logic_vector(5940, 16),
42277 => conv_std_logic_vector(6105, 16),
42278 => conv_std_logic_vector(6270, 16),
42279 => conv_std_logic_vector(6435, 16),
42280 => conv_std_logic_vector(6600, 16),
42281 => conv_std_logic_vector(6765, 16),
42282 => conv_std_logic_vector(6930, 16),
42283 => conv_std_logic_vector(7095, 16),
42284 => conv_std_logic_vector(7260, 16),
42285 => conv_std_logic_vector(7425, 16),
42286 => conv_std_logic_vector(7590, 16),
42287 => conv_std_logic_vector(7755, 16),
42288 => conv_std_logic_vector(7920, 16),
42289 => conv_std_logic_vector(8085, 16),
42290 => conv_std_logic_vector(8250, 16),
42291 => conv_std_logic_vector(8415, 16),
42292 => conv_std_logic_vector(8580, 16),
42293 => conv_std_logic_vector(8745, 16),
42294 => conv_std_logic_vector(8910, 16),
42295 => conv_std_logic_vector(9075, 16),
42296 => conv_std_logic_vector(9240, 16),
42297 => conv_std_logic_vector(9405, 16),
42298 => conv_std_logic_vector(9570, 16),
42299 => conv_std_logic_vector(9735, 16),
42300 => conv_std_logic_vector(9900, 16),
42301 => conv_std_logic_vector(10065, 16),
42302 => conv_std_logic_vector(10230, 16),
42303 => conv_std_logic_vector(10395, 16),
42304 => conv_std_logic_vector(10560, 16),
42305 => conv_std_logic_vector(10725, 16),
42306 => conv_std_logic_vector(10890, 16),
42307 => conv_std_logic_vector(11055, 16),
42308 => conv_std_logic_vector(11220, 16),
42309 => conv_std_logic_vector(11385, 16),
42310 => conv_std_logic_vector(11550, 16),
42311 => conv_std_logic_vector(11715, 16),
42312 => conv_std_logic_vector(11880, 16),
42313 => conv_std_logic_vector(12045, 16),
42314 => conv_std_logic_vector(12210, 16),
42315 => conv_std_logic_vector(12375, 16),
42316 => conv_std_logic_vector(12540, 16),
42317 => conv_std_logic_vector(12705, 16),
42318 => conv_std_logic_vector(12870, 16),
42319 => conv_std_logic_vector(13035, 16),
42320 => conv_std_logic_vector(13200, 16),
42321 => conv_std_logic_vector(13365, 16),
42322 => conv_std_logic_vector(13530, 16),
42323 => conv_std_logic_vector(13695, 16),
42324 => conv_std_logic_vector(13860, 16),
42325 => conv_std_logic_vector(14025, 16),
42326 => conv_std_logic_vector(14190, 16),
42327 => conv_std_logic_vector(14355, 16),
42328 => conv_std_logic_vector(14520, 16),
42329 => conv_std_logic_vector(14685, 16),
42330 => conv_std_logic_vector(14850, 16),
42331 => conv_std_logic_vector(15015, 16),
42332 => conv_std_logic_vector(15180, 16),
42333 => conv_std_logic_vector(15345, 16),
42334 => conv_std_logic_vector(15510, 16),
42335 => conv_std_logic_vector(15675, 16),
42336 => conv_std_logic_vector(15840, 16),
42337 => conv_std_logic_vector(16005, 16),
42338 => conv_std_logic_vector(16170, 16),
42339 => conv_std_logic_vector(16335, 16),
42340 => conv_std_logic_vector(16500, 16),
42341 => conv_std_logic_vector(16665, 16),
42342 => conv_std_logic_vector(16830, 16),
42343 => conv_std_logic_vector(16995, 16),
42344 => conv_std_logic_vector(17160, 16),
42345 => conv_std_logic_vector(17325, 16),
42346 => conv_std_logic_vector(17490, 16),
42347 => conv_std_logic_vector(17655, 16),
42348 => conv_std_logic_vector(17820, 16),
42349 => conv_std_logic_vector(17985, 16),
42350 => conv_std_logic_vector(18150, 16),
42351 => conv_std_logic_vector(18315, 16),
42352 => conv_std_logic_vector(18480, 16),
42353 => conv_std_logic_vector(18645, 16),
42354 => conv_std_logic_vector(18810, 16),
42355 => conv_std_logic_vector(18975, 16),
42356 => conv_std_logic_vector(19140, 16),
42357 => conv_std_logic_vector(19305, 16),
42358 => conv_std_logic_vector(19470, 16),
42359 => conv_std_logic_vector(19635, 16),
42360 => conv_std_logic_vector(19800, 16),
42361 => conv_std_logic_vector(19965, 16),
42362 => conv_std_logic_vector(20130, 16),
42363 => conv_std_logic_vector(20295, 16),
42364 => conv_std_logic_vector(20460, 16),
42365 => conv_std_logic_vector(20625, 16),
42366 => conv_std_logic_vector(20790, 16),
42367 => conv_std_logic_vector(20955, 16),
42368 => conv_std_logic_vector(21120, 16),
42369 => conv_std_logic_vector(21285, 16),
42370 => conv_std_logic_vector(21450, 16),
42371 => conv_std_logic_vector(21615, 16),
42372 => conv_std_logic_vector(21780, 16),
42373 => conv_std_logic_vector(21945, 16),
42374 => conv_std_logic_vector(22110, 16),
42375 => conv_std_logic_vector(22275, 16),
42376 => conv_std_logic_vector(22440, 16),
42377 => conv_std_logic_vector(22605, 16),
42378 => conv_std_logic_vector(22770, 16),
42379 => conv_std_logic_vector(22935, 16),
42380 => conv_std_logic_vector(23100, 16),
42381 => conv_std_logic_vector(23265, 16),
42382 => conv_std_logic_vector(23430, 16),
42383 => conv_std_logic_vector(23595, 16),
42384 => conv_std_logic_vector(23760, 16),
42385 => conv_std_logic_vector(23925, 16),
42386 => conv_std_logic_vector(24090, 16),
42387 => conv_std_logic_vector(24255, 16),
42388 => conv_std_logic_vector(24420, 16),
42389 => conv_std_logic_vector(24585, 16),
42390 => conv_std_logic_vector(24750, 16),
42391 => conv_std_logic_vector(24915, 16),
42392 => conv_std_logic_vector(25080, 16),
42393 => conv_std_logic_vector(25245, 16),
42394 => conv_std_logic_vector(25410, 16),
42395 => conv_std_logic_vector(25575, 16),
42396 => conv_std_logic_vector(25740, 16),
42397 => conv_std_logic_vector(25905, 16),
42398 => conv_std_logic_vector(26070, 16),
42399 => conv_std_logic_vector(26235, 16),
42400 => conv_std_logic_vector(26400, 16),
42401 => conv_std_logic_vector(26565, 16),
42402 => conv_std_logic_vector(26730, 16),
42403 => conv_std_logic_vector(26895, 16),
42404 => conv_std_logic_vector(27060, 16),
42405 => conv_std_logic_vector(27225, 16),
42406 => conv_std_logic_vector(27390, 16),
42407 => conv_std_logic_vector(27555, 16),
42408 => conv_std_logic_vector(27720, 16),
42409 => conv_std_logic_vector(27885, 16),
42410 => conv_std_logic_vector(28050, 16),
42411 => conv_std_logic_vector(28215, 16),
42412 => conv_std_logic_vector(28380, 16),
42413 => conv_std_logic_vector(28545, 16),
42414 => conv_std_logic_vector(28710, 16),
42415 => conv_std_logic_vector(28875, 16),
42416 => conv_std_logic_vector(29040, 16),
42417 => conv_std_logic_vector(29205, 16),
42418 => conv_std_logic_vector(29370, 16),
42419 => conv_std_logic_vector(29535, 16),
42420 => conv_std_logic_vector(29700, 16),
42421 => conv_std_logic_vector(29865, 16),
42422 => conv_std_logic_vector(30030, 16),
42423 => conv_std_logic_vector(30195, 16),
42424 => conv_std_logic_vector(30360, 16),
42425 => conv_std_logic_vector(30525, 16),
42426 => conv_std_logic_vector(30690, 16),
42427 => conv_std_logic_vector(30855, 16),
42428 => conv_std_logic_vector(31020, 16),
42429 => conv_std_logic_vector(31185, 16),
42430 => conv_std_logic_vector(31350, 16),
42431 => conv_std_logic_vector(31515, 16),
42432 => conv_std_logic_vector(31680, 16),
42433 => conv_std_logic_vector(31845, 16),
42434 => conv_std_logic_vector(32010, 16),
42435 => conv_std_logic_vector(32175, 16),
42436 => conv_std_logic_vector(32340, 16),
42437 => conv_std_logic_vector(32505, 16),
42438 => conv_std_logic_vector(32670, 16),
42439 => conv_std_logic_vector(32835, 16),
42440 => conv_std_logic_vector(33000, 16),
42441 => conv_std_logic_vector(33165, 16),
42442 => conv_std_logic_vector(33330, 16),
42443 => conv_std_logic_vector(33495, 16),
42444 => conv_std_logic_vector(33660, 16),
42445 => conv_std_logic_vector(33825, 16),
42446 => conv_std_logic_vector(33990, 16),
42447 => conv_std_logic_vector(34155, 16),
42448 => conv_std_logic_vector(34320, 16),
42449 => conv_std_logic_vector(34485, 16),
42450 => conv_std_logic_vector(34650, 16),
42451 => conv_std_logic_vector(34815, 16),
42452 => conv_std_logic_vector(34980, 16),
42453 => conv_std_logic_vector(35145, 16),
42454 => conv_std_logic_vector(35310, 16),
42455 => conv_std_logic_vector(35475, 16),
42456 => conv_std_logic_vector(35640, 16),
42457 => conv_std_logic_vector(35805, 16),
42458 => conv_std_logic_vector(35970, 16),
42459 => conv_std_logic_vector(36135, 16),
42460 => conv_std_logic_vector(36300, 16),
42461 => conv_std_logic_vector(36465, 16),
42462 => conv_std_logic_vector(36630, 16),
42463 => conv_std_logic_vector(36795, 16),
42464 => conv_std_logic_vector(36960, 16),
42465 => conv_std_logic_vector(37125, 16),
42466 => conv_std_logic_vector(37290, 16),
42467 => conv_std_logic_vector(37455, 16),
42468 => conv_std_logic_vector(37620, 16),
42469 => conv_std_logic_vector(37785, 16),
42470 => conv_std_logic_vector(37950, 16),
42471 => conv_std_logic_vector(38115, 16),
42472 => conv_std_logic_vector(38280, 16),
42473 => conv_std_logic_vector(38445, 16),
42474 => conv_std_logic_vector(38610, 16),
42475 => conv_std_logic_vector(38775, 16),
42476 => conv_std_logic_vector(38940, 16),
42477 => conv_std_logic_vector(39105, 16),
42478 => conv_std_logic_vector(39270, 16),
42479 => conv_std_logic_vector(39435, 16),
42480 => conv_std_logic_vector(39600, 16),
42481 => conv_std_logic_vector(39765, 16),
42482 => conv_std_logic_vector(39930, 16),
42483 => conv_std_logic_vector(40095, 16),
42484 => conv_std_logic_vector(40260, 16),
42485 => conv_std_logic_vector(40425, 16),
42486 => conv_std_logic_vector(40590, 16),
42487 => conv_std_logic_vector(40755, 16),
42488 => conv_std_logic_vector(40920, 16),
42489 => conv_std_logic_vector(41085, 16),
42490 => conv_std_logic_vector(41250, 16),
42491 => conv_std_logic_vector(41415, 16),
42492 => conv_std_logic_vector(41580, 16),
42493 => conv_std_logic_vector(41745, 16),
42494 => conv_std_logic_vector(41910, 16),
42495 => conv_std_logic_vector(42075, 16),
42496 => conv_std_logic_vector(0, 16),
42497 => conv_std_logic_vector(166, 16),
42498 => conv_std_logic_vector(332, 16),
42499 => conv_std_logic_vector(498, 16),
42500 => conv_std_logic_vector(664, 16),
42501 => conv_std_logic_vector(830, 16),
42502 => conv_std_logic_vector(996, 16),
42503 => conv_std_logic_vector(1162, 16),
42504 => conv_std_logic_vector(1328, 16),
42505 => conv_std_logic_vector(1494, 16),
42506 => conv_std_logic_vector(1660, 16),
42507 => conv_std_logic_vector(1826, 16),
42508 => conv_std_logic_vector(1992, 16),
42509 => conv_std_logic_vector(2158, 16),
42510 => conv_std_logic_vector(2324, 16),
42511 => conv_std_logic_vector(2490, 16),
42512 => conv_std_logic_vector(2656, 16),
42513 => conv_std_logic_vector(2822, 16),
42514 => conv_std_logic_vector(2988, 16),
42515 => conv_std_logic_vector(3154, 16),
42516 => conv_std_logic_vector(3320, 16),
42517 => conv_std_logic_vector(3486, 16),
42518 => conv_std_logic_vector(3652, 16),
42519 => conv_std_logic_vector(3818, 16),
42520 => conv_std_logic_vector(3984, 16),
42521 => conv_std_logic_vector(4150, 16),
42522 => conv_std_logic_vector(4316, 16),
42523 => conv_std_logic_vector(4482, 16),
42524 => conv_std_logic_vector(4648, 16),
42525 => conv_std_logic_vector(4814, 16),
42526 => conv_std_logic_vector(4980, 16),
42527 => conv_std_logic_vector(5146, 16),
42528 => conv_std_logic_vector(5312, 16),
42529 => conv_std_logic_vector(5478, 16),
42530 => conv_std_logic_vector(5644, 16),
42531 => conv_std_logic_vector(5810, 16),
42532 => conv_std_logic_vector(5976, 16),
42533 => conv_std_logic_vector(6142, 16),
42534 => conv_std_logic_vector(6308, 16),
42535 => conv_std_logic_vector(6474, 16),
42536 => conv_std_logic_vector(6640, 16),
42537 => conv_std_logic_vector(6806, 16),
42538 => conv_std_logic_vector(6972, 16),
42539 => conv_std_logic_vector(7138, 16),
42540 => conv_std_logic_vector(7304, 16),
42541 => conv_std_logic_vector(7470, 16),
42542 => conv_std_logic_vector(7636, 16),
42543 => conv_std_logic_vector(7802, 16),
42544 => conv_std_logic_vector(7968, 16),
42545 => conv_std_logic_vector(8134, 16),
42546 => conv_std_logic_vector(8300, 16),
42547 => conv_std_logic_vector(8466, 16),
42548 => conv_std_logic_vector(8632, 16),
42549 => conv_std_logic_vector(8798, 16),
42550 => conv_std_logic_vector(8964, 16),
42551 => conv_std_logic_vector(9130, 16),
42552 => conv_std_logic_vector(9296, 16),
42553 => conv_std_logic_vector(9462, 16),
42554 => conv_std_logic_vector(9628, 16),
42555 => conv_std_logic_vector(9794, 16),
42556 => conv_std_logic_vector(9960, 16),
42557 => conv_std_logic_vector(10126, 16),
42558 => conv_std_logic_vector(10292, 16),
42559 => conv_std_logic_vector(10458, 16),
42560 => conv_std_logic_vector(10624, 16),
42561 => conv_std_logic_vector(10790, 16),
42562 => conv_std_logic_vector(10956, 16),
42563 => conv_std_logic_vector(11122, 16),
42564 => conv_std_logic_vector(11288, 16),
42565 => conv_std_logic_vector(11454, 16),
42566 => conv_std_logic_vector(11620, 16),
42567 => conv_std_logic_vector(11786, 16),
42568 => conv_std_logic_vector(11952, 16),
42569 => conv_std_logic_vector(12118, 16),
42570 => conv_std_logic_vector(12284, 16),
42571 => conv_std_logic_vector(12450, 16),
42572 => conv_std_logic_vector(12616, 16),
42573 => conv_std_logic_vector(12782, 16),
42574 => conv_std_logic_vector(12948, 16),
42575 => conv_std_logic_vector(13114, 16),
42576 => conv_std_logic_vector(13280, 16),
42577 => conv_std_logic_vector(13446, 16),
42578 => conv_std_logic_vector(13612, 16),
42579 => conv_std_logic_vector(13778, 16),
42580 => conv_std_logic_vector(13944, 16),
42581 => conv_std_logic_vector(14110, 16),
42582 => conv_std_logic_vector(14276, 16),
42583 => conv_std_logic_vector(14442, 16),
42584 => conv_std_logic_vector(14608, 16),
42585 => conv_std_logic_vector(14774, 16),
42586 => conv_std_logic_vector(14940, 16),
42587 => conv_std_logic_vector(15106, 16),
42588 => conv_std_logic_vector(15272, 16),
42589 => conv_std_logic_vector(15438, 16),
42590 => conv_std_logic_vector(15604, 16),
42591 => conv_std_logic_vector(15770, 16),
42592 => conv_std_logic_vector(15936, 16),
42593 => conv_std_logic_vector(16102, 16),
42594 => conv_std_logic_vector(16268, 16),
42595 => conv_std_logic_vector(16434, 16),
42596 => conv_std_logic_vector(16600, 16),
42597 => conv_std_logic_vector(16766, 16),
42598 => conv_std_logic_vector(16932, 16),
42599 => conv_std_logic_vector(17098, 16),
42600 => conv_std_logic_vector(17264, 16),
42601 => conv_std_logic_vector(17430, 16),
42602 => conv_std_logic_vector(17596, 16),
42603 => conv_std_logic_vector(17762, 16),
42604 => conv_std_logic_vector(17928, 16),
42605 => conv_std_logic_vector(18094, 16),
42606 => conv_std_logic_vector(18260, 16),
42607 => conv_std_logic_vector(18426, 16),
42608 => conv_std_logic_vector(18592, 16),
42609 => conv_std_logic_vector(18758, 16),
42610 => conv_std_logic_vector(18924, 16),
42611 => conv_std_logic_vector(19090, 16),
42612 => conv_std_logic_vector(19256, 16),
42613 => conv_std_logic_vector(19422, 16),
42614 => conv_std_logic_vector(19588, 16),
42615 => conv_std_logic_vector(19754, 16),
42616 => conv_std_logic_vector(19920, 16),
42617 => conv_std_logic_vector(20086, 16),
42618 => conv_std_logic_vector(20252, 16),
42619 => conv_std_logic_vector(20418, 16),
42620 => conv_std_logic_vector(20584, 16),
42621 => conv_std_logic_vector(20750, 16),
42622 => conv_std_logic_vector(20916, 16),
42623 => conv_std_logic_vector(21082, 16),
42624 => conv_std_logic_vector(21248, 16),
42625 => conv_std_logic_vector(21414, 16),
42626 => conv_std_logic_vector(21580, 16),
42627 => conv_std_logic_vector(21746, 16),
42628 => conv_std_logic_vector(21912, 16),
42629 => conv_std_logic_vector(22078, 16),
42630 => conv_std_logic_vector(22244, 16),
42631 => conv_std_logic_vector(22410, 16),
42632 => conv_std_logic_vector(22576, 16),
42633 => conv_std_logic_vector(22742, 16),
42634 => conv_std_logic_vector(22908, 16),
42635 => conv_std_logic_vector(23074, 16),
42636 => conv_std_logic_vector(23240, 16),
42637 => conv_std_logic_vector(23406, 16),
42638 => conv_std_logic_vector(23572, 16),
42639 => conv_std_logic_vector(23738, 16),
42640 => conv_std_logic_vector(23904, 16),
42641 => conv_std_logic_vector(24070, 16),
42642 => conv_std_logic_vector(24236, 16),
42643 => conv_std_logic_vector(24402, 16),
42644 => conv_std_logic_vector(24568, 16),
42645 => conv_std_logic_vector(24734, 16),
42646 => conv_std_logic_vector(24900, 16),
42647 => conv_std_logic_vector(25066, 16),
42648 => conv_std_logic_vector(25232, 16),
42649 => conv_std_logic_vector(25398, 16),
42650 => conv_std_logic_vector(25564, 16),
42651 => conv_std_logic_vector(25730, 16),
42652 => conv_std_logic_vector(25896, 16),
42653 => conv_std_logic_vector(26062, 16),
42654 => conv_std_logic_vector(26228, 16),
42655 => conv_std_logic_vector(26394, 16),
42656 => conv_std_logic_vector(26560, 16),
42657 => conv_std_logic_vector(26726, 16),
42658 => conv_std_logic_vector(26892, 16),
42659 => conv_std_logic_vector(27058, 16),
42660 => conv_std_logic_vector(27224, 16),
42661 => conv_std_logic_vector(27390, 16),
42662 => conv_std_logic_vector(27556, 16),
42663 => conv_std_logic_vector(27722, 16),
42664 => conv_std_logic_vector(27888, 16),
42665 => conv_std_logic_vector(28054, 16),
42666 => conv_std_logic_vector(28220, 16),
42667 => conv_std_logic_vector(28386, 16),
42668 => conv_std_logic_vector(28552, 16),
42669 => conv_std_logic_vector(28718, 16),
42670 => conv_std_logic_vector(28884, 16),
42671 => conv_std_logic_vector(29050, 16),
42672 => conv_std_logic_vector(29216, 16),
42673 => conv_std_logic_vector(29382, 16),
42674 => conv_std_logic_vector(29548, 16),
42675 => conv_std_logic_vector(29714, 16),
42676 => conv_std_logic_vector(29880, 16),
42677 => conv_std_logic_vector(30046, 16),
42678 => conv_std_logic_vector(30212, 16),
42679 => conv_std_logic_vector(30378, 16),
42680 => conv_std_logic_vector(30544, 16),
42681 => conv_std_logic_vector(30710, 16),
42682 => conv_std_logic_vector(30876, 16),
42683 => conv_std_logic_vector(31042, 16),
42684 => conv_std_logic_vector(31208, 16),
42685 => conv_std_logic_vector(31374, 16),
42686 => conv_std_logic_vector(31540, 16),
42687 => conv_std_logic_vector(31706, 16),
42688 => conv_std_logic_vector(31872, 16),
42689 => conv_std_logic_vector(32038, 16),
42690 => conv_std_logic_vector(32204, 16),
42691 => conv_std_logic_vector(32370, 16),
42692 => conv_std_logic_vector(32536, 16),
42693 => conv_std_logic_vector(32702, 16),
42694 => conv_std_logic_vector(32868, 16),
42695 => conv_std_logic_vector(33034, 16),
42696 => conv_std_logic_vector(33200, 16),
42697 => conv_std_logic_vector(33366, 16),
42698 => conv_std_logic_vector(33532, 16),
42699 => conv_std_logic_vector(33698, 16),
42700 => conv_std_logic_vector(33864, 16),
42701 => conv_std_logic_vector(34030, 16),
42702 => conv_std_logic_vector(34196, 16),
42703 => conv_std_logic_vector(34362, 16),
42704 => conv_std_logic_vector(34528, 16),
42705 => conv_std_logic_vector(34694, 16),
42706 => conv_std_logic_vector(34860, 16),
42707 => conv_std_logic_vector(35026, 16),
42708 => conv_std_logic_vector(35192, 16),
42709 => conv_std_logic_vector(35358, 16),
42710 => conv_std_logic_vector(35524, 16),
42711 => conv_std_logic_vector(35690, 16),
42712 => conv_std_logic_vector(35856, 16),
42713 => conv_std_logic_vector(36022, 16),
42714 => conv_std_logic_vector(36188, 16),
42715 => conv_std_logic_vector(36354, 16),
42716 => conv_std_logic_vector(36520, 16),
42717 => conv_std_logic_vector(36686, 16),
42718 => conv_std_logic_vector(36852, 16),
42719 => conv_std_logic_vector(37018, 16),
42720 => conv_std_logic_vector(37184, 16),
42721 => conv_std_logic_vector(37350, 16),
42722 => conv_std_logic_vector(37516, 16),
42723 => conv_std_logic_vector(37682, 16),
42724 => conv_std_logic_vector(37848, 16),
42725 => conv_std_logic_vector(38014, 16),
42726 => conv_std_logic_vector(38180, 16),
42727 => conv_std_logic_vector(38346, 16),
42728 => conv_std_logic_vector(38512, 16),
42729 => conv_std_logic_vector(38678, 16),
42730 => conv_std_logic_vector(38844, 16),
42731 => conv_std_logic_vector(39010, 16),
42732 => conv_std_logic_vector(39176, 16),
42733 => conv_std_logic_vector(39342, 16),
42734 => conv_std_logic_vector(39508, 16),
42735 => conv_std_logic_vector(39674, 16),
42736 => conv_std_logic_vector(39840, 16),
42737 => conv_std_logic_vector(40006, 16),
42738 => conv_std_logic_vector(40172, 16),
42739 => conv_std_logic_vector(40338, 16),
42740 => conv_std_logic_vector(40504, 16),
42741 => conv_std_logic_vector(40670, 16),
42742 => conv_std_logic_vector(40836, 16),
42743 => conv_std_logic_vector(41002, 16),
42744 => conv_std_logic_vector(41168, 16),
42745 => conv_std_logic_vector(41334, 16),
42746 => conv_std_logic_vector(41500, 16),
42747 => conv_std_logic_vector(41666, 16),
42748 => conv_std_logic_vector(41832, 16),
42749 => conv_std_logic_vector(41998, 16),
42750 => conv_std_logic_vector(42164, 16),
42751 => conv_std_logic_vector(42330, 16),
42752 => conv_std_logic_vector(0, 16),
42753 => conv_std_logic_vector(167, 16),
42754 => conv_std_logic_vector(334, 16),
42755 => conv_std_logic_vector(501, 16),
42756 => conv_std_logic_vector(668, 16),
42757 => conv_std_logic_vector(835, 16),
42758 => conv_std_logic_vector(1002, 16),
42759 => conv_std_logic_vector(1169, 16),
42760 => conv_std_logic_vector(1336, 16),
42761 => conv_std_logic_vector(1503, 16),
42762 => conv_std_logic_vector(1670, 16),
42763 => conv_std_logic_vector(1837, 16),
42764 => conv_std_logic_vector(2004, 16),
42765 => conv_std_logic_vector(2171, 16),
42766 => conv_std_logic_vector(2338, 16),
42767 => conv_std_logic_vector(2505, 16),
42768 => conv_std_logic_vector(2672, 16),
42769 => conv_std_logic_vector(2839, 16),
42770 => conv_std_logic_vector(3006, 16),
42771 => conv_std_logic_vector(3173, 16),
42772 => conv_std_logic_vector(3340, 16),
42773 => conv_std_logic_vector(3507, 16),
42774 => conv_std_logic_vector(3674, 16),
42775 => conv_std_logic_vector(3841, 16),
42776 => conv_std_logic_vector(4008, 16),
42777 => conv_std_logic_vector(4175, 16),
42778 => conv_std_logic_vector(4342, 16),
42779 => conv_std_logic_vector(4509, 16),
42780 => conv_std_logic_vector(4676, 16),
42781 => conv_std_logic_vector(4843, 16),
42782 => conv_std_logic_vector(5010, 16),
42783 => conv_std_logic_vector(5177, 16),
42784 => conv_std_logic_vector(5344, 16),
42785 => conv_std_logic_vector(5511, 16),
42786 => conv_std_logic_vector(5678, 16),
42787 => conv_std_logic_vector(5845, 16),
42788 => conv_std_logic_vector(6012, 16),
42789 => conv_std_logic_vector(6179, 16),
42790 => conv_std_logic_vector(6346, 16),
42791 => conv_std_logic_vector(6513, 16),
42792 => conv_std_logic_vector(6680, 16),
42793 => conv_std_logic_vector(6847, 16),
42794 => conv_std_logic_vector(7014, 16),
42795 => conv_std_logic_vector(7181, 16),
42796 => conv_std_logic_vector(7348, 16),
42797 => conv_std_logic_vector(7515, 16),
42798 => conv_std_logic_vector(7682, 16),
42799 => conv_std_logic_vector(7849, 16),
42800 => conv_std_logic_vector(8016, 16),
42801 => conv_std_logic_vector(8183, 16),
42802 => conv_std_logic_vector(8350, 16),
42803 => conv_std_logic_vector(8517, 16),
42804 => conv_std_logic_vector(8684, 16),
42805 => conv_std_logic_vector(8851, 16),
42806 => conv_std_logic_vector(9018, 16),
42807 => conv_std_logic_vector(9185, 16),
42808 => conv_std_logic_vector(9352, 16),
42809 => conv_std_logic_vector(9519, 16),
42810 => conv_std_logic_vector(9686, 16),
42811 => conv_std_logic_vector(9853, 16),
42812 => conv_std_logic_vector(10020, 16),
42813 => conv_std_logic_vector(10187, 16),
42814 => conv_std_logic_vector(10354, 16),
42815 => conv_std_logic_vector(10521, 16),
42816 => conv_std_logic_vector(10688, 16),
42817 => conv_std_logic_vector(10855, 16),
42818 => conv_std_logic_vector(11022, 16),
42819 => conv_std_logic_vector(11189, 16),
42820 => conv_std_logic_vector(11356, 16),
42821 => conv_std_logic_vector(11523, 16),
42822 => conv_std_logic_vector(11690, 16),
42823 => conv_std_logic_vector(11857, 16),
42824 => conv_std_logic_vector(12024, 16),
42825 => conv_std_logic_vector(12191, 16),
42826 => conv_std_logic_vector(12358, 16),
42827 => conv_std_logic_vector(12525, 16),
42828 => conv_std_logic_vector(12692, 16),
42829 => conv_std_logic_vector(12859, 16),
42830 => conv_std_logic_vector(13026, 16),
42831 => conv_std_logic_vector(13193, 16),
42832 => conv_std_logic_vector(13360, 16),
42833 => conv_std_logic_vector(13527, 16),
42834 => conv_std_logic_vector(13694, 16),
42835 => conv_std_logic_vector(13861, 16),
42836 => conv_std_logic_vector(14028, 16),
42837 => conv_std_logic_vector(14195, 16),
42838 => conv_std_logic_vector(14362, 16),
42839 => conv_std_logic_vector(14529, 16),
42840 => conv_std_logic_vector(14696, 16),
42841 => conv_std_logic_vector(14863, 16),
42842 => conv_std_logic_vector(15030, 16),
42843 => conv_std_logic_vector(15197, 16),
42844 => conv_std_logic_vector(15364, 16),
42845 => conv_std_logic_vector(15531, 16),
42846 => conv_std_logic_vector(15698, 16),
42847 => conv_std_logic_vector(15865, 16),
42848 => conv_std_logic_vector(16032, 16),
42849 => conv_std_logic_vector(16199, 16),
42850 => conv_std_logic_vector(16366, 16),
42851 => conv_std_logic_vector(16533, 16),
42852 => conv_std_logic_vector(16700, 16),
42853 => conv_std_logic_vector(16867, 16),
42854 => conv_std_logic_vector(17034, 16),
42855 => conv_std_logic_vector(17201, 16),
42856 => conv_std_logic_vector(17368, 16),
42857 => conv_std_logic_vector(17535, 16),
42858 => conv_std_logic_vector(17702, 16),
42859 => conv_std_logic_vector(17869, 16),
42860 => conv_std_logic_vector(18036, 16),
42861 => conv_std_logic_vector(18203, 16),
42862 => conv_std_logic_vector(18370, 16),
42863 => conv_std_logic_vector(18537, 16),
42864 => conv_std_logic_vector(18704, 16),
42865 => conv_std_logic_vector(18871, 16),
42866 => conv_std_logic_vector(19038, 16),
42867 => conv_std_logic_vector(19205, 16),
42868 => conv_std_logic_vector(19372, 16),
42869 => conv_std_logic_vector(19539, 16),
42870 => conv_std_logic_vector(19706, 16),
42871 => conv_std_logic_vector(19873, 16),
42872 => conv_std_logic_vector(20040, 16),
42873 => conv_std_logic_vector(20207, 16),
42874 => conv_std_logic_vector(20374, 16),
42875 => conv_std_logic_vector(20541, 16),
42876 => conv_std_logic_vector(20708, 16),
42877 => conv_std_logic_vector(20875, 16),
42878 => conv_std_logic_vector(21042, 16),
42879 => conv_std_logic_vector(21209, 16),
42880 => conv_std_logic_vector(21376, 16),
42881 => conv_std_logic_vector(21543, 16),
42882 => conv_std_logic_vector(21710, 16),
42883 => conv_std_logic_vector(21877, 16),
42884 => conv_std_logic_vector(22044, 16),
42885 => conv_std_logic_vector(22211, 16),
42886 => conv_std_logic_vector(22378, 16),
42887 => conv_std_logic_vector(22545, 16),
42888 => conv_std_logic_vector(22712, 16),
42889 => conv_std_logic_vector(22879, 16),
42890 => conv_std_logic_vector(23046, 16),
42891 => conv_std_logic_vector(23213, 16),
42892 => conv_std_logic_vector(23380, 16),
42893 => conv_std_logic_vector(23547, 16),
42894 => conv_std_logic_vector(23714, 16),
42895 => conv_std_logic_vector(23881, 16),
42896 => conv_std_logic_vector(24048, 16),
42897 => conv_std_logic_vector(24215, 16),
42898 => conv_std_logic_vector(24382, 16),
42899 => conv_std_logic_vector(24549, 16),
42900 => conv_std_logic_vector(24716, 16),
42901 => conv_std_logic_vector(24883, 16),
42902 => conv_std_logic_vector(25050, 16),
42903 => conv_std_logic_vector(25217, 16),
42904 => conv_std_logic_vector(25384, 16),
42905 => conv_std_logic_vector(25551, 16),
42906 => conv_std_logic_vector(25718, 16),
42907 => conv_std_logic_vector(25885, 16),
42908 => conv_std_logic_vector(26052, 16),
42909 => conv_std_logic_vector(26219, 16),
42910 => conv_std_logic_vector(26386, 16),
42911 => conv_std_logic_vector(26553, 16),
42912 => conv_std_logic_vector(26720, 16),
42913 => conv_std_logic_vector(26887, 16),
42914 => conv_std_logic_vector(27054, 16),
42915 => conv_std_logic_vector(27221, 16),
42916 => conv_std_logic_vector(27388, 16),
42917 => conv_std_logic_vector(27555, 16),
42918 => conv_std_logic_vector(27722, 16),
42919 => conv_std_logic_vector(27889, 16),
42920 => conv_std_logic_vector(28056, 16),
42921 => conv_std_logic_vector(28223, 16),
42922 => conv_std_logic_vector(28390, 16),
42923 => conv_std_logic_vector(28557, 16),
42924 => conv_std_logic_vector(28724, 16),
42925 => conv_std_logic_vector(28891, 16),
42926 => conv_std_logic_vector(29058, 16),
42927 => conv_std_logic_vector(29225, 16),
42928 => conv_std_logic_vector(29392, 16),
42929 => conv_std_logic_vector(29559, 16),
42930 => conv_std_logic_vector(29726, 16),
42931 => conv_std_logic_vector(29893, 16),
42932 => conv_std_logic_vector(30060, 16),
42933 => conv_std_logic_vector(30227, 16),
42934 => conv_std_logic_vector(30394, 16),
42935 => conv_std_logic_vector(30561, 16),
42936 => conv_std_logic_vector(30728, 16),
42937 => conv_std_logic_vector(30895, 16),
42938 => conv_std_logic_vector(31062, 16),
42939 => conv_std_logic_vector(31229, 16),
42940 => conv_std_logic_vector(31396, 16),
42941 => conv_std_logic_vector(31563, 16),
42942 => conv_std_logic_vector(31730, 16),
42943 => conv_std_logic_vector(31897, 16),
42944 => conv_std_logic_vector(32064, 16),
42945 => conv_std_logic_vector(32231, 16),
42946 => conv_std_logic_vector(32398, 16),
42947 => conv_std_logic_vector(32565, 16),
42948 => conv_std_logic_vector(32732, 16),
42949 => conv_std_logic_vector(32899, 16),
42950 => conv_std_logic_vector(33066, 16),
42951 => conv_std_logic_vector(33233, 16),
42952 => conv_std_logic_vector(33400, 16),
42953 => conv_std_logic_vector(33567, 16),
42954 => conv_std_logic_vector(33734, 16),
42955 => conv_std_logic_vector(33901, 16),
42956 => conv_std_logic_vector(34068, 16),
42957 => conv_std_logic_vector(34235, 16),
42958 => conv_std_logic_vector(34402, 16),
42959 => conv_std_logic_vector(34569, 16),
42960 => conv_std_logic_vector(34736, 16),
42961 => conv_std_logic_vector(34903, 16),
42962 => conv_std_logic_vector(35070, 16),
42963 => conv_std_logic_vector(35237, 16),
42964 => conv_std_logic_vector(35404, 16),
42965 => conv_std_logic_vector(35571, 16),
42966 => conv_std_logic_vector(35738, 16),
42967 => conv_std_logic_vector(35905, 16),
42968 => conv_std_logic_vector(36072, 16),
42969 => conv_std_logic_vector(36239, 16),
42970 => conv_std_logic_vector(36406, 16),
42971 => conv_std_logic_vector(36573, 16),
42972 => conv_std_logic_vector(36740, 16),
42973 => conv_std_logic_vector(36907, 16),
42974 => conv_std_logic_vector(37074, 16),
42975 => conv_std_logic_vector(37241, 16),
42976 => conv_std_logic_vector(37408, 16),
42977 => conv_std_logic_vector(37575, 16),
42978 => conv_std_logic_vector(37742, 16),
42979 => conv_std_logic_vector(37909, 16),
42980 => conv_std_logic_vector(38076, 16),
42981 => conv_std_logic_vector(38243, 16),
42982 => conv_std_logic_vector(38410, 16),
42983 => conv_std_logic_vector(38577, 16),
42984 => conv_std_logic_vector(38744, 16),
42985 => conv_std_logic_vector(38911, 16),
42986 => conv_std_logic_vector(39078, 16),
42987 => conv_std_logic_vector(39245, 16),
42988 => conv_std_logic_vector(39412, 16),
42989 => conv_std_logic_vector(39579, 16),
42990 => conv_std_logic_vector(39746, 16),
42991 => conv_std_logic_vector(39913, 16),
42992 => conv_std_logic_vector(40080, 16),
42993 => conv_std_logic_vector(40247, 16),
42994 => conv_std_logic_vector(40414, 16),
42995 => conv_std_logic_vector(40581, 16),
42996 => conv_std_logic_vector(40748, 16),
42997 => conv_std_logic_vector(40915, 16),
42998 => conv_std_logic_vector(41082, 16),
42999 => conv_std_logic_vector(41249, 16),
43000 => conv_std_logic_vector(41416, 16),
43001 => conv_std_logic_vector(41583, 16),
43002 => conv_std_logic_vector(41750, 16),
43003 => conv_std_logic_vector(41917, 16),
43004 => conv_std_logic_vector(42084, 16),
43005 => conv_std_logic_vector(42251, 16),
43006 => conv_std_logic_vector(42418, 16),
43007 => conv_std_logic_vector(42585, 16),
43008 => conv_std_logic_vector(0, 16),
43009 => conv_std_logic_vector(168, 16),
43010 => conv_std_logic_vector(336, 16),
43011 => conv_std_logic_vector(504, 16),
43012 => conv_std_logic_vector(672, 16),
43013 => conv_std_logic_vector(840, 16),
43014 => conv_std_logic_vector(1008, 16),
43015 => conv_std_logic_vector(1176, 16),
43016 => conv_std_logic_vector(1344, 16),
43017 => conv_std_logic_vector(1512, 16),
43018 => conv_std_logic_vector(1680, 16),
43019 => conv_std_logic_vector(1848, 16),
43020 => conv_std_logic_vector(2016, 16),
43021 => conv_std_logic_vector(2184, 16),
43022 => conv_std_logic_vector(2352, 16),
43023 => conv_std_logic_vector(2520, 16),
43024 => conv_std_logic_vector(2688, 16),
43025 => conv_std_logic_vector(2856, 16),
43026 => conv_std_logic_vector(3024, 16),
43027 => conv_std_logic_vector(3192, 16),
43028 => conv_std_logic_vector(3360, 16),
43029 => conv_std_logic_vector(3528, 16),
43030 => conv_std_logic_vector(3696, 16),
43031 => conv_std_logic_vector(3864, 16),
43032 => conv_std_logic_vector(4032, 16),
43033 => conv_std_logic_vector(4200, 16),
43034 => conv_std_logic_vector(4368, 16),
43035 => conv_std_logic_vector(4536, 16),
43036 => conv_std_logic_vector(4704, 16),
43037 => conv_std_logic_vector(4872, 16),
43038 => conv_std_logic_vector(5040, 16),
43039 => conv_std_logic_vector(5208, 16),
43040 => conv_std_logic_vector(5376, 16),
43041 => conv_std_logic_vector(5544, 16),
43042 => conv_std_logic_vector(5712, 16),
43043 => conv_std_logic_vector(5880, 16),
43044 => conv_std_logic_vector(6048, 16),
43045 => conv_std_logic_vector(6216, 16),
43046 => conv_std_logic_vector(6384, 16),
43047 => conv_std_logic_vector(6552, 16),
43048 => conv_std_logic_vector(6720, 16),
43049 => conv_std_logic_vector(6888, 16),
43050 => conv_std_logic_vector(7056, 16),
43051 => conv_std_logic_vector(7224, 16),
43052 => conv_std_logic_vector(7392, 16),
43053 => conv_std_logic_vector(7560, 16),
43054 => conv_std_logic_vector(7728, 16),
43055 => conv_std_logic_vector(7896, 16),
43056 => conv_std_logic_vector(8064, 16),
43057 => conv_std_logic_vector(8232, 16),
43058 => conv_std_logic_vector(8400, 16),
43059 => conv_std_logic_vector(8568, 16),
43060 => conv_std_logic_vector(8736, 16),
43061 => conv_std_logic_vector(8904, 16),
43062 => conv_std_logic_vector(9072, 16),
43063 => conv_std_logic_vector(9240, 16),
43064 => conv_std_logic_vector(9408, 16),
43065 => conv_std_logic_vector(9576, 16),
43066 => conv_std_logic_vector(9744, 16),
43067 => conv_std_logic_vector(9912, 16),
43068 => conv_std_logic_vector(10080, 16),
43069 => conv_std_logic_vector(10248, 16),
43070 => conv_std_logic_vector(10416, 16),
43071 => conv_std_logic_vector(10584, 16),
43072 => conv_std_logic_vector(10752, 16),
43073 => conv_std_logic_vector(10920, 16),
43074 => conv_std_logic_vector(11088, 16),
43075 => conv_std_logic_vector(11256, 16),
43076 => conv_std_logic_vector(11424, 16),
43077 => conv_std_logic_vector(11592, 16),
43078 => conv_std_logic_vector(11760, 16),
43079 => conv_std_logic_vector(11928, 16),
43080 => conv_std_logic_vector(12096, 16),
43081 => conv_std_logic_vector(12264, 16),
43082 => conv_std_logic_vector(12432, 16),
43083 => conv_std_logic_vector(12600, 16),
43084 => conv_std_logic_vector(12768, 16),
43085 => conv_std_logic_vector(12936, 16),
43086 => conv_std_logic_vector(13104, 16),
43087 => conv_std_logic_vector(13272, 16),
43088 => conv_std_logic_vector(13440, 16),
43089 => conv_std_logic_vector(13608, 16),
43090 => conv_std_logic_vector(13776, 16),
43091 => conv_std_logic_vector(13944, 16),
43092 => conv_std_logic_vector(14112, 16),
43093 => conv_std_logic_vector(14280, 16),
43094 => conv_std_logic_vector(14448, 16),
43095 => conv_std_logic_vector(14616, 16),
43096 => conv_std_logic_vector(14784, 16),
43097 => conv_std_logic_vector(14952, 16),
43098 => conv_std_logic_vector(15120, 16),
43099 => conv_std_logic_vector(15288, 16),
43100 => conv_std_logic_vector(15456, 16),
43101 => conv_std_logic_vector(15624, 16),
43102 => conv_std_logic_vector(15792, 16),
43103 => conv_std_logic_vector(15960, 16),
43104 => conv_std_logic_vector(16128, 16),
43105 => conv_std_logic_vector(16296, 16),
43106 => conv_std_logic_vector(16464, 16),
43107 => conv_std_logic_vector(16632, 16),
43108 => conv_std_logic_vector(16800, 16),
43109 => conv_std_logic_vector(16968, 16),
43110 => conv_std_logic_vector(17136, 16),
43111 => conv_std_logic_vector(17304, 16),
43112 => conv_std_logic_vector(17472, 16),
43113 => conv_std_logic_vector(17640, 16),
43114 => conv_std_logic_vector(17808, 16),
43115 => conv_std_logic_vector(17976, 16),
43116 => conv_std_logic_vector(18144, 16),
43117 => conv_std_logic_vector(18312, 16),
43118 => conv_std_logic_vector(18480, 16),
43119 => conv_std_logic_vector(18648, 16),
43120 => conv_std_logic_vector(18816, 16),
43121 => conv_std_logic_vector(18984, 16),
43122 => conv_std_logic_vector(19152, 16),
43123 => conv_std_logic_vector(19320, 16),
43124 => conv_std_logic_vector(19488, 16),
43125 => conv_std_logic_vector(19656, 16),
43126 => conv_std_logic_vector(19824, 16),
43127 => conv_std_logic_vector(19992, 16),
43128 => conv_std_logic_vector(20160, 16),
43129 => conv_std_logic_vector(20328, 16),
43130 => conv_std_logic_vector(20496, 16),
43131 => conv_std_logic_vector(20664, 16),
43132 => conv_std_logic_vector(20832, 16),
43133 => conv_std_logic_vector(21000, 16),
43134 => conv_std_logic_vector(21168, 16),
43135 => conv_std_logic_vector(21336, 16),
43136 => conv_std_logic_vector(21504, 16),
43137 => conv_std_logic_vector(21672, 16),
43138 => conv_std_logic_vector(21840, 16),
43139 => conv_std_logic_vector(22008, 16),
43140 => conv_std_logic_vector(22176, 16),
43141 => conv_std_logic_vector(22344, 16),
43142 => conv_std_logic_vector(22512, 16),
43143 => conv_std_logic_vector(22680, 16),
43144 => conv_std_logic_vector(22848, 16),
43145 => conv_std_logic_vector(23016, 16),
43146 => conv_std_logic_vector(23184, 16),
43147 => conv_std_logic_vector(23352, 16),
43148 => conv_std_logic_vector(23520, 16),
43149 => conv_std_logic_vector(23688, 16),
43150 => conv_std_logic_vector(23856, 16),
43151 => conv_std_logic_vector(24024, 16),
43152 => conv_std_logic_vector(24192, 16),
43153 => conv_std_logic_vector(24360, 16),
43154 => conv_std_logic_vector(24528, 16),
43155 => conv_std_logic_vector(24696, 16),
43156 => conv_std_logic_vector(24864, 16),
43157 => conv_std_logic_vector(25032, 16),
43158 => conv_std_logic_vector(25200, 16),
43159 => conv_std_logic_vector(25368, 16),
43160 => conv_std_logic_vector(25536, 16),
43161 => conv_std_logic_vector(25704, 16),
43162 => conv_std_logic_vector(25872, 16),
43163 => conv_std_logic_vector(26040, 16),
43164 => conv_std_logic_vector(26208, 16),
43165 => conv_std_logic_vector(26376, 16),
43166 => conv_std_logic_vector(26544, 16),
43167 => conv_std_logic_vector(26712, 16),
43168 => conv_std_logic_vector(26880, 16),
43169 => conv_std_logic_vector(27048, 16),
43170 => conv_std_logic_vector(27216, 16),
43171 => conv_std_logic_vector(27384, 16),
43172 => conv_std_logic_vector(27552, 16),
43173 => conv_std_logic_vector(27720, 16),
43174 => conv_std_logic_vector(27888, 16),
43175 => conv_std_logic_vector(28056, 16),
43176 => conv_std_logic_vector(28224, 16),
43177 => conv_std_logic_vector(28392, 16),
43178 => conv_std_logic_vector(28560, 16),
43179 => conv_std_logic_vector(28728, 16),
43180 => conv_std_logic_vector(28896, 16),
43181 => conv_std_logic_vector(29064, 16),
43182 => conv_std_logic_vector(29232, 16),
43183 => conv_std_logic_vector(29400, 16),
43184 => conv_std_logic_vector(29568, 16),
43185 => conv_std_logic_vector(29736, 16),
43186 => conv_std_logic_vector(29904, 16),
43187 => conv_std_logic_vector(30072, 16),
43188 => conv_std_logic_vector(30240, 16),
43189 => conv_std_logic_vector(30408, 16),
43190 => conv_std_logic_vector(30576, 16),
43191 => conv_std_logic_vector(30744, 16),
43192 => conv_std_logic_vector(30912, 16),
43193 => conv_std_logic_vector(31080, 16),
43194 => conv_std_logic_vector(31248, 16),
43195 => conv_std_logic_vector(31416, 16),
43196 => conv_std_logic_vector(31584, 16),
43197 => conv_std_logic_vector(31752, 16),
43198 => conv_std_logic_vector(31920, 16),
43199 => conv_std_logic_vector(32088, 16),
43200 => conv_std_logic_vector(32256, 16),
43201 => conv_std_logic_vector(32424, 16),
43202 => conv_std_logic_vector(32592, 16),
43203 => conv_std_logic_vector(32760, 16),
43204 => conv_std_logic_vector(32928, 16),
43205 => conv_std_logic_vector(33096, 16),
43206 => conv_std_logic_vector(33264, 16),
43207 => conv_std_logic_vector(33432, 16),
43208 => conv_std_logic_vector(33600, 16),
43209 => conv_std_logic_vector(33768, 16),
43210 => conv_std_logic_vector(33936, 16),
43211 => conv_std_logic_vector(34104, 16),
43212 => conv_std_logic_vector(34272, 16),
43213 => conv_std_logic_vector(34440, 16),
43214 => conv_std_logic_vector(34608, 16),
43215 => conv_std_logic_vector(34776, 16),
43216 => conv_std_logic_vector(34944, 16),
43217 => conv_std_logic_vector(35112, 16),
43218 => conv_std_logic_vector(35280, 16),
43219 => conv_std_logic_vector(35448, 16),
43220 => conv_std_logic_vector(35616, 16),
43221 => conv_std_logic_vector(35784, 16),
43222 => conv_std_logic_vector(35952, 16),
43223 => conv_std_logic_vector(36120, 16),
43224 => conv_std_logic_vector(36288, 16),
43225 => conv_std_logic_vector(36456, 16),
43226 => conv_std_logic_vector(36624, 16),
43227 => conv_std_logic_vector(36792, 16),
43228 => conv_std_logic_vector(36960, 16),
43229 => conv_std_logic_vector(37128, 16),
43230 => conv_std_logic_vector(37296, 16),
43231 => conv_std_logic_vector(37464, 16),
43232 => conv_std_logic_vector(37632, 16),
43233 => conv_std_logic_vector(37800, 16),
43234 => conv_std_logic_vector(37968, 16),
43235 => conv_std_logic_vector(38136, 16),
43236 => conv_std_logic_vector(38304, 16),
43237 => conv_std_logic_vector(38472, 16),
43238 => conv_std_logic_vector(38640, 16),
43239 => conv_std_logic_vector(38808, 16),
43240 => conv_std_logic_vector(38976, 16),
43241 => conv_std_logic_vector(39144, 16),
43242 => conv_std_logic_vector(39312, 16),
43243 => conv_std_logic_vector(39480, 16),
43244 => conv_std_logic_vector(39648, 16),
43245 => conv_std_logic_vector(39816, 16),
43246 => conv_std_logic_vector(39984, 16),
43247 => conv_std_logic_vector(40152, 16),
43248 => conv_std_logic_vector(40320, 16),
43249 => conv_std_logic_vector(40488, 16),
43250 => conv_std_logic_vector(40656, 16),
43251 => conv_std_logic_vector(40824, 16),
43252 => conv_std_logic_vector(40992, 16),
43253 => conv_std_logic_vector(41160, 16),
43254 => conv_std_logic_vector(41328, 16),
43255 => conv_std_logic_vector(41496, 16),
43256 => conv_std_logic_vector(41664, 16),
43257 => conv_std_logic_vector(41832, 16),
43258 => conv_std_logic_vector(42000, 16),
43259 => conv_std_logic_vector(42168, 16),
43260 => conv_std_logic_vector(42336, 16),
43261 => conv_std_logic_vector(42504, 16),
43262 => conv_std_logic_vector(42672, 16),
43263 => conv_std_logic_vector(42840, 16),
43264 => conv_std_logic_vector(0, 16),
43265 => conv_std_logic_vector(169, 16),
43266 => conv_std_logic_vector(338, 16),
43267 => conv_std_logic_vector(507, 16),
43268 => conv_std_logic_vector(676, 16),
43269 => conv_std_logic_vector(845, 16),
43270 => conv_std_logic_vector(1014, 16),
43271 => conv_std_logic_vector(1183, 16),
43272 => conv_std_logic_vector(1352, 16),
43273 => conv_std_logic_vector(1521, 16),
43274 => conv_std_logic_vector(1690, 16),
43275 => conv_std_logic_vector(1859, 16),
43276 => conv_std_logic_vector(2028, 16),
43277 => conv_std_logic_vector(2197, 16),
43278 => conv_std_logic_vector(2366, 16),
43279 => conv_std_logic_vector(2535, 16),
43280 => conv_std_logic_vector(2704, 16),
43281 => conv_std_logic_vector(2873, 16),
43282 => conv_std_logic_vector(3042, 16),
43283 => conv_std_logic_vector(3211, 16),
43284 => conv_std_logic_vector(3380, 16),
43285 => conv_std_logic_vector(3549, 16),
43286 => conv_std_logic_vector(3718, 16),
43287 => conv_std_logic_vector(3887, 16),
43288 => conv_std_logic_vector(4056, 16),
43289 => conv_std_logic_vector(4225, 16),
43290 => conv_std_logic_vector(4394, 16),
43291 => conv_std_logic_vector(4563, 16),
43292 => conv_std_logic_vector(4732, 16),
43293 => conv_std_logic_vector(4901, 16),
43294 => conv_std_logic_vector(5070, 16),
43295 => conv_std_logic_vector(5239, 16),
43296 => conv_std_logic_vector(5408, 16),
43297 => conv_std_logic_vector(5577, 16),
43298 => conv_std_logic_vector(5746, 16),
43299 => conv_std_logic_vector(5915, 16),
43300 => conv_std_logic_vector(6084, 16),
43301 => conv_std_logic_vector(6253, 16),
43302 => conv_std_logic_vector(6422, 16),
43303 => conv_std_logic_vector(6591, 16),
43304 => conv_std_logic_vector(6760, 16),
43305 => conv_std_logic_vector(6929, 16),
43306 => conv_std_logic_vector(7098, 16),
43307 => conv_std_logic_vector(7267, 16),
43308 => conv_std_logic_vector(7436, 16),
43309 => conv_std_logic_vector(7605, 16),
43310 => conv_std_logic_vector(7774, 16),
43311 => conv_std_logic_vector(7943, 16),
43312 => conv_std_logic_vector(8112, 16),
43313 => conv_std_logic_vector(8281, 16),
43314 => conv_std_logic_vector(8450, 16),
43315 => conv_std_logic_vector(8619, 16),
43316 => conv_std_logic_vector(8788, 16),
43317 => conv_std_logic_vector(8957, 16),
43318 => conv_std_logic_vector(9126, 16),
43319 => conv_std_logic_vector(9295, 16),
43320 => conv_std_logic_vector(9464, 16),
43321 => conv_std_logic_vector(9633, 16),
43322 => conv_std_logic_vector(9802, 16),
43323 => conv_std_logic_vector(9971, 16),
43324 => conv_std_logic_vector(10140, 16),
43325 => conv_std_logic_vector(10309, 16),
43326 => conv_std_logic_vector(10478, 16),
43327 => conv_std_logic_vector(10647, 16),
43328 => conv_std_logic_vector(10816, 16),
43329 => conv_std_logic_vector(10985, 16),
43330 => conv_std_logic_vector(11154, 16),
43331 => conv_std_logic_vector(11323, 16),
43332 => conv_std_logic_vector(11492, 16),
43333 => conv_std_logic_vector(11661, 16),
43334 => conv_std_logic_vector(11830, 16),
43335 => conv_std_logic_vector(11999, 16),
43336 => conv_std_logic_vector(12168, 16),
43337 => conv_std_logic_vector(12337, 16),
43338 => conv_std_logic_vector(12506, 16),
43339 => conv_std_logic_vector(12675, 16),
43340 => conv_std_logic_vector(12844, 16),
43341 => conv_std_logic_vector(13013, 16),
43342 => conv_std_logic_vector(13182, 16),
43343 => conv_std_logic_vector(13351, 16),
43344 => conv_std_logic_vector(13520, 16),
43345 => conv_std_logic_vector(13689, 16),
43346 => conv_std_logic_vector(13858, 16),
43347 => conv_std_logic_vector(14027, 16),
43348 => conv_std_logic_vector(14196, 16),
43349 => conv_std_logic_vector(14365, 16),
43350 => conv_std_logic_vector(14534, 16),
43351 => conv_std_logic_vector(14703, 16),
43352 => conv_std_logic_vector(14872, 16),
43353 => conv_std_logic_vector(15041, 16),
43354 => conv_std_logic_vector(15210, 16),
43355 => conv_std_logic_vector(15379, 16),
43356 => conv_std_logic_vector(15548, 16),
43357 => conv_std_logic_vector(15717, 16),
43358 => conv_std_logic_vector(15886, 16),
43359 => conv_std_logic_vector(16055, 16),
43360 => conv_std_logic_vector(16224, 16),
43361 => conv_std_logic_vector(16393, 16),
43362 => conv_std_logic_vector(16562, 16),
43363 => conv_std_logic_vector(16731, 16),
43364 => conv_std_logic_vector(16900, 16),
43365 => conv_std_logic_vector(17069, 16),
43366 => conv_std_logic_vector(17238, 16),
43367 => conv_std_logic_vector(17407, 16),
43368 => conv_std_logic_vector(17576, 16),
43369 => conv_std_logic_vector(17745, 16),
43370 => conv_std_logic_vector(17914, 16),
43371 => conv_std_logic_vector(18083, 16),
43372 => conv_std_logic_vector(18252, 16),
43373 => conv_std_logic_vector(18421, 16),
43374 => conv_std_logic_vector(18590, 16),
43375 => conv_std_logic_vector(18759, 16),
43376 => conv_std_logic_vector(18928, 16),
43377 => conv_std_logic_vector(19097, 16),
43378 => conv_std_logic_vector(19266, 16),
43379 => conv_std_logic_vector(19435, 16),
43380 => conv_std_logic_vector(19604, 16),
43381 => conv_std_logic_vector(19773, 16),
43382 => conv_std_logic_vector(19942, 16),
43383 => conv_std_logic_vector(20111, 16),
43384 => conv_std_logic_vector(20280, 16),
43385 => conv_std_logic_vector(20449, 16),
43386 => conv_std_logic_vector(20618, 16),
43387 => conv_std_logic_vector(20787, 16),
43388 => conv_std_logic_vector(20956, 16),
43389 => conv_std_logic_vector(21125, 16),
43390 => conv_std_logic_vector(21294, 16),
43391 => conv_std_logic_vector(21463, 16),
43392 => conv_std_logic_vector(21632, 16),
43393 => conv_std_logic_vector(21801, 16),
43394 => conv_std_logic_vector(21970, 16),
43395 => conv_std_logic_vector(22139, 16),
43396 => conv_std_logic_vector(22308, 16),
43397 => conv_std_logic_vector(22477, 16),
43398 => conv_std_logic_vector(22646, 16),
43399 => conv_std_logic_vector(22815, 16),
43400 => conv_std_logic_vector(22984, 16),
43401 => conv_std_logic_vector(23153, 16),
43402 => conv_std_logic_vector(23322, 16),
43403 => conv_std_logic_vector(23491, 16),
43404 => conv_std_logic_vector(23660, 16),
43405 => conv_std_logic_vector(23829, 16),
43406 => conv_std_logic_vector(23998, 16),
43407 => conv_std_logic_vector(24167, 16),
43408 => conv_std_logic_vector(24336, 16),
43409 => conv_std_logic_vector(24505, 16),
43410 => conv_std_logic_vector(24674, 16),
43411 => conv_std_logic_vector(24843, 16),
43412 => conv_std_logic_vector(25012, 16),
43413 => conv_std_logic_vector(25181, 16),
43414 => conv_std_logic_vector(25350, 16),
43415 => conv_std_logic_vector(25519, 16),
43416 => conv_std_logic_vector(25688, 16),
43417 => conv_std_logic_vector(25857, 16),
43418 => conv_std_logic_vector(26026, 16),
43419 => conv_std_logic_vector(26195, 16),
43420 => conv_std_logic_vector(26364, 16),
43421 => conv_std_logic_vector(26533, 16),
43422 => conv_std_logic_vector(26702, 16),
43423 => conv_std_logic_vector(26871, 16),
43424 => conv_std_logic_vector(27040, 16),
43425 => conv_std_logic_vector(27209, 16),
43426 => conv_std_logic_vector(27378, 16),
43427 => conv_std_logic_vector(27547, 16),
43428 => conv_std_logic_vector(27716, 16),
43429 => conv_std_logic_vector(27885, 16),
43430 => conv_std_logic_vector(28054, 16),
43431 => conv_std_logic_vector(28223, 16),
43432 => conv_std_logic_vector(28392, 16),
43433 => conv_std_logic_vector(28561, 16),
43434 => conv_std_logic_vector(28730, 16),
43435 => conv_std_logic_vector(28899, 16),
43436 => conv_std_logic_vector(29068, 16),
43437 => conv_std_logic_vector(29237, 16),
43438 => conv_std_logic_vector(29406, 16),
43439 => conv_std_logic_vector(29575, 16),
43440 => conv_std_logic_vector(29744, 16),
43441 => conv_std_logic_vector(29913, 16),
43442 => conv_std_logic_vector(30082, 16),
43443 => conv_std_logic_vector(30251, 16),
43444 => conv_std_logic_vector(30420, 16),
43445 => conv_std_logic_vector(30589, 16),
43446 => conv_std_logic_vector(30758, 16),
43447 => conv_std_logic_vector(30927, 16),
43448 => conv_std_logic_vector(31096, 16),
43449 => conv_std_logic_vector(31265, 16),
43450 => conv_std_logic_vector(31434, 16),
43451 => conv_std_logic_vector(31603, 16),
43452 => conv_std_logic_vector(31772, 16),
43453 => conv_std_logic_vector(31941, 16),
43454 => conv_std_logic_vector(32110, 16),
43455 => conv_std_logic_vector(32279, 16),
43456 => conv_std_logic_vector(32448, 16),
43457 => conv_std_logic_vector(32617, 16),
43458 => conv_std_logic_vector(32786, 16),
43459 => conv_std_logic_vector(32955, 16),
43460 => conv_std_logic_vector(33124, 16),
43461 => conv_std_logic_vector(33293, 16),
43462 => conv_std_logic_vector(33462, 16),
43463 => conv_std_logic_vector(33631, 16),
43464 => conv_std_logic_vector(33800, 16),
43465 => conv_std_logic_vector(33969, 16),
43466 => conv_std_logic_vector(34138, 16),
43467 => conv_std_logic_vector(34307, 16),
43468 => conv_std_logic_vector(34476, 16),
43469 => conv_std_logic_vector(34645, 16),
43470 => conv_std_logic_vector(34814, 16),
43471 => conv_std_logic_vector(34983, 16),
43472 => conv_std_logic_vector(35152, 16),
43473 => conv_std_logic_vector(35321, 16),
43474 => conv_std_logic_vector(35490, 16),
43475 => conv_std_logic_vector(35659, 16),
43476 => conv_std_logic_vector(35828, 16),
43477 => conv_std_logic_vector(35997, 16),
43478 => conv_std_logic_vector(36166, 16),
43479 => conv_std_logic_vector(36335, 16),
43480 => conv_std_logic_vector(36504, 16),
43481 => conv_std_logic_vector(36673, 16),
43482 => conv_std_logic_vector(36842, 16),
43483 => conv_std_logic_vector(37011, 16),
43484 => conv_std_logic_vector(37180, 16),
43485 => conv_std_logic_vector(37349, 16),
43486 => conv_std_logic_vector(37518, 16),
43487 => conv_std_logic_vector(37687, 16),
43488 => conv_std_logic_vector(37856, 16),
43489 => conv_std_logic_vector(38025, 16),
43490 => conv_std_logic_vector(38194, 16),
43491 => conv_std_logic_vector(38363, 16),
43492 => conv_std_logic_vector(38532, 16),
43493 => conv_std_logic_vector(38701, 16),
43494 => conv_std_logic_vector(38870, 16),
43495 => conv_std_logic_vector(39039, 16),
43496 => conv_std_logic_vector(39208, 16),
43497 => conv_std_logic_vector(39377, 16),
43498 => conv_std_logic_vector(39546, 16),
43499 => conv_std_logic_vector(39715, 16),
43500 => conv_std_logic_vector(39884, 16),
43501 => conv_std_logic_vector(40053, 16),
43502 => conv_std_logic_vector(40222, 16),
43503 => conv_std_logic_vector(40391, 16),
43504 => conv_std_logic_vector(40560, 16),
43505 => conv_std_logic_vector(40729, 16),
43506 => conv_std_logic_vector(40898, 16),
43507 => conv_std_logic_vector(41067, 16),
43508 => conv_std_logic_vector(41236, 16),
43509 => conv_std_logic_vector(41405, 16),
43510 => conv_std_logic_vector(41574, 16),
43511 => conv_std_logic_vector(41743, 16),
43512 => conv_std_logic_vector(41912, 16),
43513 => conv_std_logic_vector(42081, 16),
43514 => conv_std_logic_vector(42250, 16),
43515 => conv_std_logic_vector(42419, 16),
43516 => conv_std_logic_vector(42588, 16),
43517 => conv_std_logic_vector(42757, 16),
43518 => conv_std_logic_vector(42926, 16),
43519 => conv_std_logic_vector(43095, 16),
43520 => conv_std_logic_vector(0, 16),
43521 => conv_std_logic_vector(170, 16),
43522 => conv_std_logic_vector(340, 16),
43523 => conv_std_logic_vector(510, 16),
43524 => conv_std_logic_vector(680, 16),
43525 => conv_std_logic_vector(850, 16),
43526 => conv_std_logic_vector(1020, 16),
43527 => conv_std_logic_vector(1190, 16),
43528 => conv_std_logic_vector(1360, 16),
43529 => conv_std_logic_vector(1530, 16),
43530 => conv_std_logic_vector(1700, 16),
43531 => conv_std_logic_vector(1870, 16),
43532 => conv_std_logic_vector(2040, 16),
43533 => conv_std_logic_vector(2210, 16),
43534 => conv_std_logic_vector(2380, 16),
43535 => conv_std_logic_vector(2550, 16),
43536 => conv_std_logic_vector(2720, 16),
43537 => conv_std_logic_vector(2890, 16),
43538 => conv_std_logic_vector(3060, 16),
43539 => conv_std_logic_vector(3230, 16),
43540 => conv_std_logic_vector(3400, 16),
43541 => conv_std_logic_vector(3570, 16),
43542 => conv_std_logic_vector(3740, 16),
43543 => conv_std_logic_vector(3910, 16),
43544 => conv_std_logic_vector(4080, 16),
43545 => conv_std_logic_vector(4250, 16),
43546 => conv_std_logic_vector(4420, 16),
43547 => conv_std_logic_vector(4590, 16),
43548 => conv_std_logic_vector(4760, 16),
43549 => conv_std_logic_vector(4930, 16),
43550 => conv_std_logic_vector(5100, 16),
43551 => conv_std_logic_vector(5270, 16),
43552 => conv_std_logic_vector(5440, 16),
43553 => conv_std_logic_vector(5610, 16),
43554 => conv_std_logic_vector(5780, 16),
43555 => conv_std_logic_vector(5950, 16),
43556 => conv_std_logic_vector(6120, 16),
43557 => conv_std_logic_vector(6290, 16),
43558 => conv_std_logic_vector(6460, 16),
43559 => conv_std_logic_vector(6630, 16),
43560 => conv_std_logic_vector(6800, 16),
43561 => conv_std_logic_vector(6970, 16),
43562 => conv_std_logic_vector(7140, 16),
43563 => conv_std_logic_vector(7310, 16),
43564 => conv_std_logic_vector(7480, 16),
43565 => conv_std_logic_vector(7650, 16),
43566 => conv_std_logic_vector(7820, 16),
43567 => conv_std_logic_vector(7990, 16),
43568 => conv_std_logic_vector(8160, 16),
43569 => conv_std_logic_vector(8330, 16),
43570 => conv_std_logic_vector(8500, 16),
43571 => conv_std_logic_vector(8670, 16),
43572 => conv_std_logic_vector(8840, 16),
43573 => conv_std_logic_vector(9010, 16),
43574 => conv_std_logic_vector(9180, 16),
43575 => conv_std_logic_vector(9350, 16),
43576 => conv_std_logic_vector(9520, 16),
43577 => conv_std_logic_vector(9690, 16),
43578 => conv_std_logic_vector(9860, 16),
43579 => conv_std_logic_vector(10030, 16),
43580 => conv_std_logic_vector(10200, 16),
43581 => conv_std_logic_vector(10370, 16),
43582 => conv_std_logic_vector(10540, 16),
43583 => conv_std_logic_vector(10710, 16),
43584 => conv_std_logic_vector(10880, 16),
43585 => conv_std_logic_vector(11050, 16),
43586 => conv_std_logic_vector(11220, 16),
43587 => conv_std_logic_vector(11390, 16),
43588 => conv_std_logic_vector(11560, 16),
43589 => conv_std_logic_vector(11730, 16),
43590 => conv_std_logic_vector(11900, 16),
43591 => conv_std_logic_vector(12070, 16),
43592 => conv_std_logic_vector(12240, 16),
43593 => conv_std_logic_vector(12410, 16),
43594 => conv_std_logic_vector(12580, 16),
43595 => conv_std_logic_vector(12750, 16),
43596 => conv_std_logic_vector(12920, 16),
43597 => conv_std_logic_vector(13090, 16),
43598 => conv_std_logic_vector(13260, 16),
43599 => conv_std_logic_vector(13430, 16),
43600 => conv_std_logic_vector(13600, 16),
43601 => conv_std_logic_vector(13770, 16),
43602 => conv_std_logic_vector(13940, 16),
43603 => conv_std_logic_vector(14110, 16),
43604 => conv_std_logic_vector(14280, 16),
43605 => conv_std_logic_vector(14450, 16),
43606 => conv_std_logic_vector(14620, 16),
43607 => conv_std_logic_vector(14790, 16),
43608 => conv_std_logic_vector(14960, 16),
43609 => conv_std_logic_vector(15130, 16),
43610 => conv_std_logic_vector(15300, 16),
43611 => conv_std_logic_vector(15470, 16),
43612 => conv_std_logic_vector(15640, 16),
43613 => conv_std_logic_vector(15810, 16),
43614 => conv_std_logic_vector(15980, 16),
43615 => conv_std_logic_vector(16150, 16),
43616 => conv_std_logic_vector(16320, 16),
43617 => conv_std_logic_vector(16490, 16),
43618 => conv_std_logic_vector(16660, 16),
43619 => conv_std_logic_vector(16830, 16),
43620 => conv_std_logic_vector(17000, 16),
43621 => conv_std_logic_vector(17170, 16),
43622 => conv_std_logic_vector(17340, 16),
43623 => conv_std_logic_vector(17510, 16),
43624 => conv_std_logic_vector(17680, 16),
43625 => conv_std_logic_vector(17850, 16),
43626 => conv_std_logic_vector(18020, 16),
43627 => conv_std_logic_vector(18190, 16),
43628 => conv_std_logic_vector(18360, 16),
43629 => conv_std_logic_vector(18530, 16),
43630 => conv_std_logic_vector(18700, 16),
43631 => conv_std_logic_vector(18870, 16),
43632 => conv_std_logic_vector(19040, 16),
43633 => conv_std_logic_vector(19210, 16),
43634 => conv_std_logic_vector(19380, 16),
43635 => conv_std_logic_vector(19550, 16),
43636 => conv_std_logic_vector(19720, 16),
43637 => conv_std_logic_vector(19890, 16),
43638 => conv_std_logic_vector(20060, 16),
43639 => conv_std_logic_vector(20230, 16),
43640 => conv_std_logic_vector(20400, 16),
43641 => conv_std_logic_vector(20570, 16),
43642 => conv_std_logic_vector(20740, 16),
43643 => conv_std_logic_vector(20910, 16),
43644 => conv_std_logic_vector(21080, 16),
43645 => conv_std_logic_vector(21250, 16),
43646 => conv_std_logic_vector(21420, 16),
43647 => conv_std_logic_vector(21590, 16),
43648 => conv_std_logic_vector(21760, 16),
43649 => conv_std_logic_vector(21930, 16),
43650 => conv_std_logic_vector(22100, 16),
43651 => conv_std_logic_vector(22270, 16),
43652 => conv_std_logic_vector(22440, 16),
43653 => conv_std_logic_vector(22610, 16),
43654 => conv_std_logic_vector(22780, 16),
43655 => conv_std_logic_vector(22950, 16),
43656 => conv_std_logic_vector(23120, 16),
43657 => conv_std_logic_vector(23290, 16),
43658 => conv_std_logic_vector(23460, 16),
43659 => conv_std_logic_vector(23630, 16),
43660 => conv_std_logic_vector(23800, 16),
43661 => conv_std_logic_vector(23970, 16),
43662 => conv_std_logic_vector(24140, 16),
43663 => conv_std_logic_vector(24310, 16),
43664 => conv_std_logic_vector(24480, 16),
43665 => conv_std_logic_vector(24650, 16),
43666 => conv_std_logic_vector(24820, 16),
43667 => conv_std_logic_vector(24990, 16),
43668 => conv_std_logic_vector(25160, 16),
43669 => conv_std_logic_vector(25330, 16),
43670 => conv_std_logic_vector(25500, 16),
43671 => conv_std_logic_vector(25670, 16),
43672 => conv_std_logic_vector(25840, 16),
43673 => conv_std_logic_vector(26010, 16),
43674 => conv_std_logic_vector(26180, 16),
43675 => conv_std_logic_vector(26350, 16),
43676 => conv_std_logic_vector(26520, 16),
43677 => conv_std_logic_vector(26690, 16),
43678 => conv_std_logic_vector(26860, 16),
43679 => conv_std_logic_vector(27030, 16),
43680 => conv_std_logic_vector(27200, 16),
43681 => conv_std_logic_vector(27370, 16),
43682 => conv_std_logic_vector(27540, 16),
43683 => conv_std_logic_vector(27710, 16),
43684 => conv_std_logic_vector(27880, 16),
43685 => conv_std_logic_vector(28050, 16),
43686 => conv_std_logic_vector(28220, 16),
43687 => conv_std_logic_vector(28390, 16),
43688 => conv_std_logic_vector(28560, 16),
43689 => conv_std_logic_vector(28730, 16),
43690 => conv_std_logic_vector(28900, 16),
43691 => conv_std_logic_vector(29070, 16),
43692 => conv_std_logic_vector(29240, 16),
43693 => conv_std_logic_vector(29410, 16),
43694 => conv_std_logic_vector(29580, 16),
43695 => conv_std_logic_vector(29750, 16),
43696 => conv_std_logic_vector(29920, 16),
43697 => conv_std_logic_vector(30090, 16),
43698 => conv_std_logic_vector(30260, 16),
43699 => conv_std_logic_vector(30430, 16),
43700 => conv_std_logic_vector(30600, 16),
43701 => conv_std_logic_vector(30770, 16),
43702 => conv_std_logic_vector(30940, 16),
43703 => conv_std_logic_vector(31110, 16),
43704 => conv_std_logic_vector(31280, 16),
43705 => conv_std_logic_vector(31450, 16),
43706 => conv_std_logic_vector(31620, 16),
43707 => conv_std_logic_vector(31790, 16),
43708 => conv_std_logic_vector(31960, 16),
43709 => conv_std_logic_vector(32130, 16),
43710 => conv_std_logic_vector(32300, 16),
43711 => conv_std_logic_vector(32470, 16),
43712 => conv_std_logic_vector(32640, 16),
43713 => conv_std_logic_vector(32810, 16),
43714 => conv_std_logic_vector(32980, 16),
43715 => conv_std_logic_vector(33150, 16),
43716 => conv_std_logic_vector(33320, 16),
43717 => conv_std_logic_vector(33490, 16),
43718 => conv_std_logic_vector(33660, 16),
43719 => conv_std_logic_vector(33830, 16),
43720 => conv_std_logic_vector(34000, 16),
43721 => conv_std_logic_vector(34170, 16),
43722 => conv_std_logic_vector(34340, 16),
43723 => conv_std_logic_vector(34510, 16),
43724 => conv_std_logic_vector(34680, 16),
43725 => conv_std_logic_vector(34850, 16),
43726 => conv_std_logic_vector(35020, 16),
43727 => conv_std_logic_vector(35190, 16),
43728 => conv_std_logic_vector(35360, 16),
43729 => conv_std_logic_vector(35530, 16),
43730 => conv_std_logic_vector(35700, 16),
43731 => conv_std_logic_vector(35870, 16),
43732 => conv_std_logic_vector(36040, 16),
43733 => conv_std_logic_vector(36210, 16),
43734 => conv_std_logic_vector(36380, 16),
43735 => conv_std_logic_vector(36550, 16),
43736 => conv_std_logic_vector(36720, 16),
43737 => conv_std_logic_vector(36890, 16),
43738 => conv_std_logic_vector(37060, 16),
43739 => conv_std_logic_vector(37230, 16),
43740 => conv_std_logic_vector(37400, 16),
43741 => conv_std_logic_vector(37570, 16),
43742 => conv_std_logic_vector(37740, 16),
43743 => conv_std_logic_vector(37910, 16),
43744 => conv_std_logic_vector(38080, 16),
43745 => conv_std_logic_vector(38250, 16),
43746 => conv_std_logic_vector(38420, 16),
43747 => conv_std_logic_vector(38590, 16),
43748 => conv_std_logic_vector(38760, 16),
43749 => conv_std_logic_vector(38930, 16),
43750 => conv_std_logic_vector(39100, 16),
43751 => conv_std_logic_vector(39270, 16),
43752 => conv_std_logic_vector(39440, 16),
43753 => conv_std_logic_vector(39610, 16),
43754 => conv_std_logic_vector(39780, 16),
43755 => conv_std_logic_vector(39950, 16),
43756 => conv_std_logic_vector(40120, 16),
43757 => conv_std_logic_vector(40290, 16),
43758 => conv_std_logic_vector(40460, 16),
43759 => conv_std_logic_vector(40630, 16),
43760 => conv_std_logic_vector(40800, 16),
43761 => conv_std_logic_vector(40970, 16),
43762 => conv_std_logic_vector(41140, 16),
43763 => conv_std_logic_vector(41310, 16),
43764 => conv_std_logic_vector(41480, 16),
43765 => conv_std_logic_vector(41650, 16),
43766 => conv_std_logic_vector(41820, 16),
43767 => conv_std_logic_vector(41990, 16),
43768 => conv_std_logic_vector(42160, 16),
43769 => conv_std_logic_vector(42330, 16),
43770 => conv_std_logic_vector(42500, 16),
43771 => conv_std_logic_vector(42670, 16),
43772 => conv_std_logic_vector(42840, 16),
43773 => conv_std_logic_vector(43010, 16),
43774 => conv_std_logic_vector(43180, 16),
43775 => conv_std_logic_vector(43350, 16),
43776 => conv_std_logic_vector(0, 16),
43777 => conv_std_logic_vector(171, 16),
43778 => conv_std_logic_vector(342, 16),
43779 => conv_std_logic_vector(513, 16),
43780 => conv_std_logic_vector(684, 16),
43781 => conv_std_logic_vector(855, 16),
43782 => conv_std_logic_vector(1026, 16),
43783 => conv_std_logic_vector(1197, 16),
43784 => conv_std_logic_vector(1368, 16),
43785 => conv_std_logic_vector(1539, 16),
43786 => conv_std_logic_vector(1710, 16),
43787 => conv_std_logic_vector(1881, 16),
43788 => conv_std_logic_vector(2052, 16),
43789 => conv_std_logic_vector(2223, 16),
43790 => conv_std_logic_vector(2394, 16),
43791 => conv_std_logic_vector(2565, 16),
43792 => conv_std_logic_vector(2736, 16),
43793 => conv_std_logic_vector(2907, 16),
43794 => conv_std_logic_vector(3078, 16),
43795 => conv_std_logic_vector(3249, 16),
43796 => conv_std_logic_vector(3420, 16),
43797 => conv_std_logic_vector(3591, 16),
43798 => conv_std_logic_vector(3762, 16),
43799 => conv_std_logic_vector(3933, 16),
43800 => conv_std_logic_vector(4104, 16),
43801 => conv_std_logic_vector(4275, 16),
43802 => conv_std_logic_vector(4446, 16),
43803 => conv_std_logic_vector(4617, 16),
43804 => conv_std_logic_vector(4788, 16),
43805 => conv_std_logic_vector(4959, 16),
43806 => conv_std_logic_vector(5130, 16),
43807 => conv_std_logic_vector(5301, 16),
43808 => conv_std_logic_vector(5472, 16),
43809 => conv_std_logic_vector(5643, 16),
43810 => conv_std_logic_vector(5814, 16),
43811 => conv_std_logic_vector(5985, 16),
43812 => conv_std_logic_vector(6156, 16),
43813 => conv_std_logic_vector(6327, 16),
43814 => conv_std_logic_vector(6498, 16),
43815 => conv_std_logic_vector(6669, 16),
43816 => conv_std_logic_vector(6840, 16),
43817 => conv_std_logic_vector(7011, 16),
43818 => conv_std_logic_vector(7182, 16),
43819 => conv_std_logic_vector(7353, 16),
43820 => conv_std_logic_vector(7524, 16),
43821 => conv_std_logic_vector(7695, 16),
43822 => conv_std_logic_vector(7866, 16),
43823 => conv_std_logic_vector(8037, 16),
43824 => conv_std_logic_vector(8208, 16),
43825 => conv_std_logic_vector(8379, 16),
43826 => conv_std_logic_vector(8550, 16),
43827 => conv_std_logic_vector(8721, 16),
43828 => conv_std_logic_vector(8892, 16),
43829 => conv_std_logic_vector(9063, 16),
43830 => conv_std_logic_vector(9234, 16),
43831 => conv_std_logic_vector(9405, 16),
43832 => conv_std_logic_vector(9576, 16),
43833 => conv_std_logic_vector(9747, 16),
43834 => conv_std_logic_vector(9918, 16),
43835 => conv_std_logic_vector(10089, 16),
43836 => conv_std_logic_vector(10260, 16),
43837 => conv_std_logic_vector(10431, 16),
43838 => conv_std_logic_vector(10602, 16),
43839 => conv_std_logic_vector(10773, 16),
43840 => conv_std_logic_vector(10944, 16),
43841 => conv_std_logic_vector(11115, 16),
43842 => conv_std_logic_vector(11286, 16),
43843 => conv_std_logic_vector(11457, 16),
43844 => conv_std_logic_vector(11628, 16),
43845 => conv_std_logic_vector(11799, 16),
43846 => conv_std_logic_vector(11970, 16),
43847 => conv_std_logic_vector(12141, 16),
43848 => conv_std_logic_vector(12312, 16),
43849 => conv_std_logic_vector(12483, 16),
43850 => conv_std_logic_vector(12654, 16),
43851 => conv_std_logic_vector(12825, 16),
43852 => conv_std_logic_vector(12996, 16),
43853 => conv_std_logic_vector(13167, 16),
43854 => conv_std_logic_vector(13338, 16),
43855 => conv_std_logic_vector(13509, 16),
43856 => conv_std_logic_vector(13680, 16),
43857 => conv_std_logic_vector(13851, 16),
43858 => conv_std_logic_vector(14022, 16),
43859 => conv_std_logic_vector(14193, 16),
43860 => conv_std_logic_vector(14364, 16),
43861 => conv_std_logic_vector(14535, 16),
43862 => conv_std_logic_vector(14706, 16),
43863 => conv_std_logic_vector(14877, 16),
43864 => conv_std_logic_vector(15048, 16),
43865 => conv_std_logic_vector(15219, 16),
43866 => conv_std_logic_vector(15390, 16),
43867 => conv_std_logic_vector(15561, 16),
43868 => conv_std_logic_vector(15732, 16),
43869 => conv_std_logic_vector(15903, 16),
43870 => conv_std_logic_vector(16074, 16),
43871 => conv_std_logic_vector(16245, 16),
43872 => conv_std_logic_vector(16416, 16),
43873 => conv_std_logic_vector(16587, 16),
43874 => conv_std_logic_vector(16758, 16),
43875 => conv_std_logic_vector(16929, 16),
43876 => conv_std_logic_vector(17100, 16),
43877 => conv_std_logic_vector(17271, 16),
43878 => conv_std_logic_vector(17442, 16),
43879 => conv_std_logic_vector(17613, 16),
43880 => conv_std_logic_vector(17784, 16),
43881 => conv_std_logic_vector(17955, 16),
43882 => conv_std_logic_vector(18126, 16),
43883 => conv_std_logic_vector(18297, 16),
43884 => conv_std_logic_vector(18468, 16),
43885 => conv_std_logic_vector(18639, 16),
43886 => conv_std_logic_vector(18810, 16),
43887 => conv_std_logic_vector(18981, 16),
43888 => conv_std_logic_vector(19152, 16),
43889 => conv_std_logic_vector(19323, 16),
43890 => conv_std_logic_vector(19494, 16),
43891 => conv_std_logic_vector(19665, 16),
43892 => conv_std_logic_vector(19836, 16),
43893 => conv_std_logic_vector(20007, 16),
43894 => conv_std_logic_vector(20178, 16),
43895 => conv_std_logic_vector(20349, 16),
43896 => conv_std_logic_vector(20520, 16),
43897 => conv_std_logic_vector(20691, 16),
43898 => conv_std_logic_vector(20862, 16),
43899 => conv_std_logic_vector(21033, 16),
43900 => conv_std_logic_vector(21204, 16),
43901 => conv_std_logic_vector(21375, 16),
43902 => conv_std_logic_vector(21546, 16),
43903 => conv_std_logic_vector(21717, 16),
43904 => conv_std_logic_vector(21888, 16),
43905 => conv_std_logic_vector(22059, 16),
43906 => conv_std_logic_vector(22230, 16),
43907 => conv_std_logic_vector(22401, 16),
43908 => conv_std_logic_vector(22572, 16),
43909 => conv_std_logic_vector(22743, 16),
43910 => conv_std_logic_vector(22914, 16),
43911 => conv_std_logic_vector(23085, 16),
43912 => conv_std_logic_vector(23256, 16),
43913 => conv_std_logic_vector(23427, 16),
43914 => conv_std_logic_vector(23598, 16),
43915 => conv_std_logic_vector(23769, 16),
43916 => conv_std_logic_vector(23940, 16),
43917 => conv_std_logic_vector(24111, 16),
43918 => conv_std_logic_vector(24282, 16),
43919 => conv_std_logic_vector(24453, 16),
43920 => conv_std_logic_vector(24624, 16),
43921 => conv_std_logic_vector(24795, 16),
43922 => conv_std_logic_vector(24966, 16),
43923 => conv_std_logic_vector(25137, 16),
43924 => conv_std_logic_vector(25308, 16),
43925 => conv_std_logic_vector(25479, 16),
43926 => conv_std_logic_vector(25650, 16),
43927 => conv_std_logic_vector(25821, 16),
43928 => conv_std_logic_vector(25992, 16),
43929 => conv_std_logic_vector(26163, 16),
43930 => conv_std_logic_vector(26334, 16),
43931 => conv_std_logic_vector(26505, 16),
43932 => conv_std_logic_vector(26676, 16),
43933 => conv_std_logic_vector(26847, 16),
43934 => conv_std_logic_vector(27018, 16),
43935 => conv_std_logic_vector(27189, 16),
43936 => conv_std_logic_vector(27360, 16),
43937 => conv_std_logic_vector(27531, 16),
43938 => conv_std_logic_vector(27702, 16),
43939 => conv_std_logic_vector(27873, 16),
43940 => conv_std_logic_vector(28044, 16),
43941 => conv_std_logic_vector(28215, 16),
43942 => conv_std_logic_vector(28386, 16),
43943 => conv_std_logic_vector(28557, 16),
43944 => conv_std_logic_vector(28728, 16),
43945 => conv_std_logic_vector(28899, 16),
43946 => conv_std_logic_vector(29070, 16),
43947 => conv_std_logic_vector(29241, 16),
43948 => conv_std_logic_vector(29412, 16),
43949 => conv_std_logic_vector(29583, 16),
43950 => conv_std_logic_vector(29754, 16),
43951 => conv_std_logic_vector(29925, 16),
43952 => conv_std_logic_vector(30096, 16),
43953 => conv_std_logic_vector(30267, 16),
43954 => conv_std_logic_vector(30438, 16),
43955 => conv_std_logic_vector(30609, 16),
43956 => conv_std_logic_vector(30780, 16),
43957 => conv_std_logic_vector(30951, 16),
43958 => conv_std_logic_vector(31122, 16),
43959 => conv_std_logic_vector(31293, 16),
43960 => conv_std_logic_vector(31464, 16),
43961 => conv_std_logic_vector(31635, 16),
43962 => conv_std_logic_vector(31806, 16),
43963 => conv_std_logic_vector(31977, 16),
43964 => conv_std_logic_vector(32148, 16),
43965 => conv_std_logic_vector(32319, 16),
43966 => conv_std_logic_vector(32490, 16),
43967 => conv_std_logic_vector(32661, 16),
43968 => conv_std_logic_vector(32832, 16),
43969 => conv_std_logic_vector(33003, 16),
43970 => conv_std_logic_vector(33174, 16),
43971 => conv_std_logic_vector(33345, 16),
43972 => conv_std_logic_vector(33516, 16),
43973 => conv_std_logic_vector(33687, 16),
43974 => conv_std_logic_vector(33858, 16),
43975 => conv_std_logic_vector(34029, 16),
43976 => conv_std_logic_vector(34200, 16),
43977 => conv_std_logic_vector(34371, 16),
43978 => conv_std_logic_vector(34542, 16),
43979 => conv_std_logic_vector(34713, 16),
43980 => conv_std_logic_vector(34884, 16),
43981 => conv_std_logic_vector(35055, 16),
43982 => conv_std_logic_vector(35226, 16),
43983 => conv_std_logic_vector(35397, 16),
43984 => conv_std_logic_vector(35568, 16),
43985 => conv_std_logic_vector(35739, 16),
43986 => conv_std_logic_vector(35910, 16),
43987 => conv_std_logic_vector(36081, 16),
43988 => conv_std_logic_vector(36252, 16),
43989 => conv_std_logic_vector(36423, 16),
43990 => conv_std_logic_vector(36594, 16),
43991 => conv_std_logic_vector(36765, 16),
43992 => conv_std_logic_vector(36936, 16),
43993 => conv_std_logic_vector(37107, 16),
43994 => conv_std_logic_vector(37278, 16),
43995 => conv_std_logic_vector(37449, 16),
43996 => conv_std_logic_vector(37620, 16),
43997 => conv_std_logic_vector(37791, 16),
43998 => conv_std_logic_vector(37962, 16),
43999 => conv_std_logic_vector(38133, 16),
44000 => conv_std_logic_vector(38304, 16),
44001 => conv_std_logic_vector(38475, 16),
44002 => conv_std_logic_vector(38646, 16),
44003 => conv_std_logic_vector(38817, 16),
44004 => conv_std_logic_vector(38988, 16),
44005 => conv_std_logic_vector(39159, 16),
44006 => conv_std_logic_vector(39330, 16),
44007 => conv_std_logic_vector(39501, 16),
44008 => conv_std_logic_vector(39672, 16),
44009 => conv_std_logic_vector(39843, 16),
44010 => conv_std_logic_vector(40014, 16),
44011 => conv_std_logic_vector(40185, 16),
44012 => conv_std_logic_vector(40356, 16),
44013 => conv_std_logic_vector(40527, 16),
44014 => conv_std_logic_vector(40698, 16),
44015 => conv_std_logic_vector(40869, 16),
44016 => conv_std_logic_vector(41040, 16),
44017 => conv_std_logic_vector(41211, 16),
44018 => conv_std_logic_vector(41382, 16),
44019 => conv_std_logic_vector(41553, 16),
44020 => conv_std_logic_vector(41724, 16),
44021 => conv_std_logic_vector(41895, 16),
44022 => conv_std_logic_vector(42066, 16),
44023 => conv_std_logic_vector(42237, 16),
44024 => conv_std_logic_vector(42408, 16),
44025 => conv_std_logic_vector(42579, 16),
44026 => conv_std_logic_vector(42750, 16),
44027 => conv_std_logic_vector(42921, 16),
44028 => conv_std_logic_vector(43092, 16),
44029 => conv_std_logic_vector(43263, 16),
44030 => conv_std_logic_vector(43434, 16),
44031 => conv_std_logic_vector(43605, 16),
44032 => conv_std_logic_vector(0, 16),
44033 => conv_std_logic_vector(172, 16),
44034 => conv_std_logic_vector(344, 16),
44035 => conv_std_logic_vector(516, 16),
44036 => conv_std_logic_vector(688, 16),
44037 => conv_std_logic_vector(860, 16),
44038 => conv_std_logic_vector(1032, 16),
44039 => conv_std_logic_vector(1204, 16),
44040 => conv_std_logic_vector(1376, 16),
44041 => conv_std_logic_vector(1548, 16),
44042 => conv_std_logic_vector(1720, 16),
44043 => conv_std_logic_vector(1892, 16),
44044 => conv_std_logic_vector(2064, 16),
44045 => conv_std_logic_vector(2236, 16),
44046 => conv_std_logic_vector(2408, 16),
44047 => conv_std_logic_vector(2580, 16),
44048 => conv_std_logic_vector(2752, 16),
44049 => conv_std_logic_vector(2924, 16),
44050 => conv_std_logic_vector(3096, 16),
44051 => conv_std_logic_vector(3268, 16),
44052 => conv_std_logic_vector(3440, 16),
44053 => conv_std_logic_vector(3612, 16),
44054 => conv_std_logic_vector(3784, 16),
44055 => conv_std_logic_vector(3956, 16),
44056 => conv_std_logic_vector(4128, 16),
44057 => conv_std_logic_vector(4300, 16),
44058 => conv_std_logic_vector(4472, 16),
44059 => conv_std_logic_vector(4644, 16),
44060 => conv_std_logic_vector(4816, 16),
44061 => conv_std_logic_vector(4988, 16),
44062 => conv_std_logic_vector(5160, 16),
44063 => conv_std_logic_vector(5332, 16),
44064 => conv_std_logic_vector(5504, 16),
44065 => conv_std_logic_vector(5676, 16),
44066 => conv_std_logic_vector(5848, 16),
44067 => conv_std_logic_vector(6020, 16),
44068 => conv_std_logic_vector(6192, 16),
44069 => conv_std_logic_vector(6364, 16),
44070 => conv_std_logic_vector(6536, 16),
44071 => conv_std_logic_vector(6708, 16),
44072 => conv_std_logic_vector(6880, 16),
44073 => conv_std_logic_vector(7052, 16),
44074 => conv_std_logic_vector(7224, 16),
44075 => conv_std_logic_vector(7396, 16),
44076 => conv_std_logic_vector(7568, 16),
44077 => conv_std_logic_vector(7740, 16),
44078 => conv_std_logic_vector(7912, 16),
44079 => conv_std_logic_vector(8084, 16),
44080 => conv_std_logic_vector(8256, 16),
44081 => conv_std_logic_vector(8428, 16),
44082 => conv_std_logic_vector(8600, 16),
44083 => conv_std_logic_vector(8772, 16),
44084 => conv_std_logic_vector(8944, 16),
44085 => conv_std_logic_vector(9116, 16),
44086 => conv_std_logic_vector(9288, 16),
44087 => conv_std_logic_vector(9460, 16),
44088 => conv_std_logic_vector(9632, 16),
44089 => conv_std_logic_vector(9804, 16),
44090 => conv_std_logic_vector(9976, 16),
44091 => conv_std_logic_vector(10148, 16),
44092 => conv_std_logic_vector(10320, 16),
44093 => conv_std_logic_vector(10492, 16),
44094 => conv_std_logic_vector(10664, 16),
44095 => conv_std_logic_vector(10836, 16),
44096 => conv_std_logic_vector(11008, 16),
44097 => conv_std_logic_vector(11180, 16),
44098 => conv_std_logic_vector(11352, 16),
44099 => conv_std_logic_vector(11524, 16),
44100 => conv_std_logic_vector(11696, 16),
44101 => conv_std_logic_vector(11868, 16),
44102 => conv_std_logic_vector(12040, 16),
44103 => conv_std_logic_vector(12212, 16),
44104 => conv_std_logic_vector(12384, 16),
44105 => conv_std_logic_vector(12556, 16),
44106 => conv_std_logic_vector(12728, 16),
44107 => conv_std_logic_vector(12900, 16),
44108 => conv_std_logic_vector(13072, 16),
44109 => conv_std_logic_vector(13244, 16),
44110 => conv_std_logic_vector(13416, 16),
44111 => conv_std_logic_vector(13588, 16),
44112 => conv_std_logic_vector(13760, 16),
44113 => conv_std_logic_vector(13932, 16),
44114 => conv_std_logic_vector(14104, 16),
44115 => conv_std_logic_vector(14276, 16),
44116 => conv_std_logic_vector(14448, 16),
44117 => conv_std_logic_vector(14620, 16),
44118 => conv_std_logic_vector(14792, 16),
44119 => conv_std_logic_vector(14964, 16),
44120 => conv_std_logic_vector(15136, 16),
44121 => conv_std_logic_vector(15308, 16),
44122 => conv_std_logic_vector(15480, 16),
44123 => conv_std_logic_vector(15652, 16),
44124 => conv_std_logic_vector(15824, 16),
44125 => conv_std_logic_vector(15996, 16),
44126 => conv_std_logic_vector(16168, 16),
44127 => conv_std_logic_vector(16340, 16),
44128 => conv_std_logic_vector(16512, 16),
44129 => conv_std_logic_vector(16684, 16),
44130 => conv_std_logic_vector(16856, 16),
44131 => conv_std_logic_vector(17028, 16),
44132 => conv_std_logic_vector(17200, 16),
44133 => conv_std_logic_vector(17372, 16),
44134 => conv_std_logic_vector(17544, 16),
44135 => conv_std_logic_vector(17716, 16),
44136 => conv_std_logic_vector(17888, 16),
44137 => conv_std_logic_vector(18060, 16),
44138 => conv_std_logic_vector(18232, 16),
44139 => conv_std_logic_vector(18404, 16),
44140 => conv_std_logic_vector(18576, 16),
44141 => conv_std_logic_vector(18748, 16),
44142 => conv_std_logic_vector(18920, 16),
44143 => conv_std_logic_vector(19092, 16),
44144 => conv_std_logic_vector(19264, 16),
44145 => conv_std_logic_vector(19436, 16),
44146 => conv_std_logic_vector(19608, 16),
44147 => conv_std_logic_vector(19780, 16),
44148 => conv_std_logic_vector(19952, 16),
44149 => conv_std_logic_vector(20124, 16),
44150 => conv_std_logic_vector(20296, 16),
44151 => conv_std_logic_vector(20468, 16),
44152 => conv_std_logic_vector(20640, 16),
44153 => conv_std_logic_vector(20812, 16),
44154 => conv_std_logic_vector(20984, 16),
44155 => conv_std_logic_vector(21156, 16),
44156 => conv_std_logic_vector(21328, 16),
44157 => conv_std_logic_vector(21500, 16),
44158 => conv_std_logic_vector(21672, 16),
44159 => conv_std_logic_vector(21844, 16),
44160 => conv_std_logic_vector(22016, 16),
44161 => conv_std_logic_vector(22188, 16),
44162 => conv_std_logic_vector(22360, 16),
44163 => conv_std_logic_vector(22532, 16),
44164 => conv_std_logic_vector(22704, 16),
44165 => conv_std_logic_vector(22876, 16),
44166 => conv_std_logic_vector(23048, 16),
44167 => conv_std_logic_vector(23220, 16),
44168 => conv_std_logic_vector(23392, 16),
44169 => conv_std_logic_vector(23564, 16),
44170 => conv_std_logic_vector(23736, 16),
44171 => conv_std_logic_vector(23908, 16),
44172 => conv_std_logic_vector(24080, 16),
44173 => conv_std_logic_vector(24252, 16),
44174 => conv_std_logic_vector(24424, 16),
44175 => conv_std_logic_vector(24596, 16),
44176 => conv_std_logic_vector(24768, 16),
44177 => conv_std_logic_vector(24940, 16),
44178 => conv_std_logic_vector(25112, 16),
44179 => conv_std_logic_vector(25284, 16),
44180 => conv_std_logic_vector(25456, 16),
44181 => conv_std_logic_vector(25628, 16),
44182 => conv_std_logic_vector(25800, 16),
44183 => conv_std_logic_vector(25972, 16),
44184 => conv_std_logic_vector(26144, 16),
44185 => conv_std_logic_vector(26316, 16),
44186 => conv_std_logic_vector(26488, 16),
44187 => conv_std_logic_vector(26660, 16),
44188 => conv_std_logic_vector(26832, 16),
44189 => conv_std_logic_vector(27004, 16),
44190 => conv_std_logic_vector(27176, 16),
44191 => conv_std_logic_vector(27348, 16),
44192 => conv_std_logic_vector(27520, 16),
44193 => conv_std_logic_vector(27692, 16),
44194 => conv_std_logic_vector(27864, 16),
44195 => conv_std_logic_vector(28036, 16),
44196 => conv_std_logic_vector(28208, 16),
44197 => conv_std_logic_vector(28380, 16),
44198 => conv_std_logic_vector(28552, 16),
44199 => conv_std_logic_vector(28724, 16),
44200 => conv_std_logic_vector(28896, 16),
44201 => conv_std_logic_vector(29068, 16),
44202 => conv_std_logic_vector(29240, 16),
44203 => conv_std_logic_vector(29412, 16),
44204 => conv_std_logic_vector(29584, 16),
44205 => conv_std_logic_vector(29756, 16),
44206 => conv_std_logic_vector(29928, 16),
44207 => conv_std_logic_vector(30100, 16),
44208 => conv_std_logic_vector(30272, 16),
44209 => conv_std_logic_vector(30444, 16),
44210 => conv_std_logic_vector(30616, 16),
44211 => conv_std_logic_vector(30788, 16),
44212 => conv_std_logic_vector(30960, 16),
44213 => conv_std_logic_vector(31132, 16),
44214 => conv_std_logic_vector(31304, 16),
44215 => conv_std_logic_vector(31476, 16),
44216 => conv_std_logic_vector(31648, 16),
44217 => conv_std_logic_vector(31820, 16),
44218 => conv_std_logic_vector(31992, 16),
44219 => conv_std_logic_vector(32164, 16),
44220 => conv_std_logic_vector(32336, 16),
44221 => conv_std_logic_vector(32508, 16),
44222 => conv_std_logic_vector(32680, 16),
44223 => conv_std_logic_vector(32852, 16),
44224 => conv_std_logic_vector(33024, 16),
44225 => conv_std_logic_vector(33196, 16),
44226 => conv_std_logic_vector(33368, 16),
44227 => conv_std_logic_vector(33540, 16),
44228 => conv_std_logic_vector(33712, 16),
44229 => conv_std_logic_vector(33884, 16),
44230 => conv_std_logic_vector(34056, 16),
44231 => conv_std_logic_vector(34228, 16),
44232 => conv_std_logic_vector(34400, 16),
44233 => conv_std_logic_vector(34572, 16),
44234 => conv_std_logic_vector(34744, 16),
44235 => conv_std_logic_vector(34916, 16),
44236 => conv_std_logic_vector(35088, 16),
44237 => conv_std_logic_vector(35260, 16),
44238 => conv_std_logic_vector(35432, 16),
44239 => conv_std_logic_vector(35604, 16),
44240 => conv_std_logic_vector(35776, 16),
44241 => conv_std_logic_vector(35948, 16),
44242 => conv_std_logic_vector(36120, 16),
44243 => conv_std_logic_vector(36292, 16),
44244 => conv_std_logic_vector(36464, 16),
44245 => conv_std_logic_vector(36636, 16),
44246 => conv_std_logic_vector(36808, 16),
44247 => conv_std_logic_vector(36980, 16),
44248 => conv_std_logic_vector(37152, 16),
44249 => conv_std_logic_vector(37324, 16),
44250 => conv_std_logic_vector(37496, 16),
44251 => conv_std_logic_vector(37668, 16),
44252 => conv_std_logic_vector(37840, 16),
44253 => conv_std_logic_vector(38012, 16),
44254 => conv_std_logic_vector(38184, 16),
44255 => conv_std_logic_vector(38356, 16),
44256 => conv_std_logic_vector(38528, 16),
44257 => conv_std_logic_vector(38700, 16),
44258 => conv_std_logic_vector(38872, 16),
44259 => conv_std_logic_vector(39044, 16),
44260 => conv_std_logic_vector(39216, 16),
44261 => conv_std_logic_vector(39388, 16),
44262 => conv_std_logic_vector(39560, 16),
44263 => conv_std_logic_vector(39732, 16),
44264 => conv_std_logic_vector(39904, 16),
44265 => conv_std_logic_vector(40076, 16),
44266 => conv_std_logic_vector(40248, 16),
44267 => conv_std_logic_vector(40420, 16),
44268 => conv_std_logic_vector(40592, 16),
44269 => conv_std_logic_vector(40764, 16),
44270 => conv_std_logic_vector(40936, 16),
44271 => conv_std_logic_vector(41108, 16),
44272 => conv_std_logic_vector(41280, 16),
44273 => conv_std_logic_vector(41452, 16),
44274 => conv_std_logic_vector(41624, 16),
44275 => conv_std_logic_vector(41796, 16),
44276 => conv_std_logic_vector(41968, 16),
44277 => conv_std_logic_vector(42140, 16),
44278 => conv_std_logic_vector(42312, 16),
44279 => conv_std_logic_vector(42484, 16),
44280 => conv_std_logic_vector(42656, 16),
44281 => conv_std_logic_vector(42828, 16),
44282 => conv_std_logic_vector(43000, 16),
44283 => conv_std_logic_vector(43172, 16),
44284 => conv_std_logic_vector(43344, 16),
44285 => conv_std_logic_vector(43516, 16),
44286 => conv_std_logic_vector(43688, 16),
44287 => conv_std_logic_vector(43860, 16),
44288 => conv_std_logic_vector(0, 16),
44289 => conv_std_logic_vector(173, 16),
44290 => conv_std_logic_vector(346, 16),
44291 => conv_std_logic_vector(519, 16),
44292 => conv_std_logic_vector(692, 16),
44293 => conv_std_logic_vector(865, 16),
44294 => conv_std_logic_vector(1038, 16),
44295 => conv_std_logic_vector(1211, 16),
44296 => conv_std_logic_vector(1384, 16),
44297 => conv_std_logic_vector(1557, 16),
44298 => conv_std_logic_vector(1730, 16),
44299 => conv_std_logic_vector(1903, 16),
44300 => conv_std_logic_vector(2076, 16),
44301 => conv_std_logic_vector(2249, 16),
44302 => conv_std_logic_vector(2422, 16),
44303 => conv_std_logic_vector(2595, 16),
44304 => conv_std_logic_vector(2768, 16),
44305 => conv_std_logic_vector(2941, 16),
44306 => conv_std_logic_vector(3114, 16),
44307 => conv_std_logic_vector(3287, 16),
44308 => conv_std_logic_vector(3460, 16),
44309 => conv_std_logic_vector(3633, 16),
44310 => conv_std_logic_vector(3806, 16),
44311 => conv_std_logic_vector(3979, 16),
44312 => conv_std_logic_vector(4152, 16),
44313 => conv_std_logic_vector(4325, 16),
44314 => conv_std_logic_vector(4498, 16),
44315 => conv_std_logic_vector(4671, 16),
44316 => conv_std_logic_vector(4844, 16),
44317 => conv_std_logic_vector(5017, 16),
44318 => conv_std_logic_vector(5190, 16),
44319 => conv_std_logic_vector(5363, 16),
44320 => conv_std_logic_vector(5536, 16),
44321 => conv_std_logic_vector(5709, 16),
44322 => conv_std_logic_vector(5882, 16),
44323 => conv_std_logic_vector(6055, 16),
44324 => conv_std_logic_vector(6228, 16),
44325 => conv_std_logic_vector(6401, 16),
44326 => conv_std_logic_vector(6574, 16),
44327 => conv_std_logic_vector(6747, 16),
44328 => conv_std_logic_vector(6920, 16),
44329 => conv_std_logic_vector(7093, 16),
44330 => conv_std_logic_vector(7266, 16),
44331 => conv_std_logic_vector(7439, 16),
44332 => conv_std_logic_vector(7612, 16),
44333 => conv_std_logic_vector(7785, 16),
44334 => conv_std_logic_vector(7958, 16),
44335 => conv_std_logic_vector(8131, 16),
44336 => conv_std_logic_vector(8304, 16),
44337 => conv_std_logic_vector(8477, 16),
44338 => conv_std_logic_vector(8650, 16),
44339 => conv_std_logic_vector(8823, 16),
44340 => conv_std_logic_vector(8996, 16),
44341 => conv_std_logic_vector(9169, 16),
44342 => conv_std_logic_vector(9342, 16),
44343 => conv_std_logic_vector(9515, 16),
44344 => conv_std_logic_vector(9688, 16),
44345 => conv_std_logic_vector(9861, 16),
44346 => conv_std_logic_vector(10034, 16),
44347 => conv_std_logic_vector(10207, 16),
44348 => conv_std_logic_vector(10380, 16),
44349 => conv_std_logic_vector(10553, 16),
44350 => conv_std_logic_vector(10726, 16),
44351 => conv_std_logic_vector(10899, 16),
44352 => conv_std_logic_vector(11072, 16),
44353 => conv_std_logic_vector(11245, 16),
44354 => conv_std_logic_vector(11418, 16),
44355 => conv_std_logic_vector(11591, 16),
44356 => conv_std_logic_vector(11764, 16),
44357 => conv_std_logic_vector(11937, 16),
44358 => conv_std_logic_vector(12110, 16),
44359 => conv_std_logic_vector(12283, 16),
44360 => conv_std_logic_vector(12456, 16),
44361 => conv_std_logic_vector(12629, 16),
44362 => conv_std_logic_vector(12802, 16),
44363 => conv_std_logic_vector(12975, 16),
44364 => conv_std_logic_vector(13148, 16),
44365 => conv_std_logic_vector(13321, 16),
44366 => conv_std_logic_vector(13494, 16),
44367 => conv_std_logic_vector(13667, 16),
44368 => conv_std_logic_vector(13840, 16),
44369 => conv_std_logic_vector(14013, 16),
44370 => conv_std_logic_vector(14186, 16),
44371 => conv_std_logic_vector(14359, 16),
44372 => conv_std_logic_vector(14532, 16),
44373 => conv_std_logic_vector(14705, 16),
44374 => conv_std_logic_vector(14878, 16),
44375 => conv_std_logic_vector(15051, 16),
44376 => conv_std_logic_vector(15224, 16),
44377 => conv_std_logic_vector(15397, 16),
44378 => conv_std_logic_vector(15570, 16),
44379 => conv_std_logic_vector(15743, 16),
44380 => conv_std_logic_vector(15916, 16),
44381 => conv_std_logic_vector(16089, 16),
44382 => conv_std_logic_vector(16262, 16),
44383 => conv_std_logic_vector(16435, 16),
44384 => conv_std_logic_vector(16608, 16),
44385 => conv_std_logic_vector(16781, 16),
44386 => conv_std_logic_vector(16954, 16),
44387 => conv_std_logic_vector(17127, 16),
44388 => conv_std_logic_vector(17300, 16),
44389 => conv_std_logic_vector(17473, 16),
44390 => conv_std_logic_vector(17646, 16),
44391 => conv_std_logic_vector(17819, 16),
44392 => conv_std_logic_vector(17992, 16),
44393 => conv_std_logic_vector(18165, 16),
44394 => conv_std_logic_vector(18338, 16),
44395 => conv_std_logic_vector(18511, 16),
44396 => conv_std_logic_vector(18684, 16),
44397 => conv_std_logic_vector(18857, 16),
44398 => conv_std_logic_vector(19030, 16),
44399 => conv_std_logic_vector(19203, 16),
44400 => conv_std_logic_vector(19376, 16),
44401 => conv_std_logic_vector(19549, 16),
44402 => conv_std_logic_vector(19722, 16),
44403 => conv_std_logic_vector(19895, 16),
44404 => conv_std_logic_vector(20068, 16),
44405 => conv_std_logic_vector(20241, 16),
44406 => conv_std_logic_vector(20414, 16),
44407 => conv_std_logic_vector(20587, 16),
44408 => conv_std_logic_vector(20760, 16),
44409 => conv_std_logic_vector(20933, 16),
44410 => conv_std_logic_vector(21106, 16),
44411 => conv_std_logic_vector(21279, 16),
44412 => conv_std_logic_vector(21452, 16),
44413 => conv_std_logic_vector(21625, 16),
44414 => conv_std_logic_vector(21798, 16),
44415 => conv_std_logic_vector(21971, 16),
44416 => conv_std_logic_vector(22144, 16),
44417 => conv_std_logic_vector(22317, 16),
44418 => conv_std_logic_vector(22490, 16),
44419 => conv_std_logic_vector(22663, 16),
44420 => conv_std_logic_vector(22836, 16),
44421 => conv_std_logic_vector(23009, 16),
44422 => conv_std_logic_vector(23182, 16),
44423 => conv_std_logic_vector(23355, 16),
44424 => conv_std_logic_vector(23528, 16),
44425 => conv_std_logic_vector(23701, 16),
44426 => conv_std_logic_vector(23874, 16),
44427 => conv_std_logic_vector(24047, 16),
44428 => conv_std_logic_vector(24220, 16),
44429 => conv_std_logic_vector(24393, 16),
44430 => conv_std_logic_vector(24566, 16),
44431 => conv_std_logic_vector(24739, 16),
44432 => conv_std_logic_vector(24912, 16),
44433 => conv_std_logic_vector(25085, 16),
44434 => conv_std_logic_vector(25258, 16),
44435 => conv_std_logic_vector(25431, 16),
44436 => conv_std_logic_vector(25604, 16),
44437 => conv_std_logic_vector(25777, 16),
44438 => conv_std_logic_vector(25950, 16),
44439 => conv_std_logic_vector(26123, 16),
44440 => conv_std_logic_vector(26296, 16),
44441 => conv_std_logic_vector(26469, 16),
44442 => conv_std_logic_vector(26642, 16),
44443 => conv_std_logic_vector(26815, 16),
44444 => conv_std_logic_vector(26988, 16),
44445 => conv_std_logic_vector(27161, 16),
44446 => conv_std_logic_vector(27334, 16),
44447 => conv_std_logic_vector(27507, 16),
44448 => conv_std_logic_vector(27680, 16),
44449 => conv_std_logic_vector(27853, 16),
44450 => conv_std_logic_vector(28026, 16),
44451 => conv_std_logic_vector(28199, 16),
44452 => conv_std_logic_vector(28372, 16),
44453 => conv_std_logic_vector(28545, 16),
44454 => conv_std_logic_vector(28718, 16),
44455 => conv_std_logic_vector(28891, 16),
44456 => conv_std_logic_vector(29064, 16),
44457 => conv_std_logic_vector(29237, 16),
44458 => conv_std_logic_vector(29410, 16),
44459 => conv_std_logic_vector(29583, 16),
44460 => conv_std_logic_vector(29756, 16),
44461 => conv_std_logic_vector(29929, 16),
44462 => conv_std_logic_vector(30102, 16),
44463 => conv_std_logic_vector(30275, 16),
44464 => conv_std_logic_vector(30448, 16),
44465 => conv_std_logic_vector(30621, 16),
44466 => conv_std_logic_vector(30794, 16),
44467 => conv_std_logic_vector(30967, 16),
44468 => conv_std_logic_vector(31140, 16),
44469 => conv_std_logic_vector(31313, 16),
44470 => conv_std_logic_vector(31486, 16),
44471 => conv_std_logic_vector(31659, 16),
44472 => conv_std_logic_vector(31832, 16),
44473 => conv_std_logic_vector(32005, 16),
44474 => conv_std_logic_vector(32178, 16),
44475 => conv_std_logic_vector(32351, 16),
44476 => conv_std_logic_vector(32524, 16),
44477 => conv_std_logic_vector(32697, 16),
44478 => conv_std_logic_vector(32870, 16),
44479 => conv_std_logic_vector(33043, 16),
44480 => conv_std_logic_vector(33216, 16),
44481 => conv_std_logic_vector(33389, 16),
44482 => conv_std_logic_vector(33562, 16),
44483 => conv_std_logic_vector(33735, 16),
44484 => conv_std_logic_vector(33908, 16),
44485 => conv_std_logic_vector(34081, 16),
44486 => conv_std_logic_vector(34254, 16),
44487 => conv_std_logic_vector(34427, 16),
44488 => conv_std_logic_vector(34600, 16),
44489 => conv_std_logic_vector(34773, 16),
44490 => conv_std_logic_vector(34946, 16),
44491 => conv_std_logic_vector(35119, 16),
44492 => conv_std_logic_vector(35292, 16),
44493 => conv_std_logic_vector(35465, 16),
44494 => conv_std_logic_vector(35638, 16),
44495 => conv_std_logic_vector(35811, 16),
44496 => conv_std_logic_vector(35984, 16),
44497 => conv_std_logic_vector(36157, 16),
44498 => conv_std_logic_vector(36330, 16),
44499 => conv_std_logic_vector(36503, 16),
44500 => conv_std_logic_vector(36676, 16),
44501 => conv_std_logic_vector(36849, 16),
44502 => conv_std_logic_vector(37022, 16),
44503 => conv_std_logic_vector(37195, 16),
44504 => conv_std_logic_vector(37368, 16),
44505 => conv_std_logic_vector(37541, 16),
44506 => conv_std_logic_vector(37714, 16),
44507 => conv_std_logic_vector(37887, 16),
44508 => conv_std_logic_vector(38060, 16),
44509 => conv_std_logic_vector(38233, 16),
44510 => conv_std_logic_vector(38406, 16),
44511 => conv_std_logic_vector(38579, 16),
44512 => conv_std_logic_vector(38752, 16),
44513 => conv_std_logic_vector(38925, 16),
44514 => conv_std_logic_vector(39098, 16),
44515 => conv_std_logic_vector(39271, 16),
44516 => conv_std_logic_vector(39444, 16),
44517 => conv_std_logic_vector(39617, 16),
44518 => conv_std_logic_vector(39790, 16),
44519 => conv_std_logic_vector(39963, 16),
44520 => conv_std_logic_vector(40136, 16),
44521 => conv_std_logic_vector(40309, 16),
44522 => conv_std_logic_vector(40482, 16),
44523 => conv_std_logic_vector(40655, 16),
44524 => conv_std_logic_vector(40828, 16),
44525 => conv_std_logic_vector(41001, 16),
44526 => conv_std_logic_vector(41174, 16),
44527 => conv_std_logic_vector(41347, 16),
44528 => conv_std_logic_vector(41520, 16),
44529 => conv_std_logic_vector(41693, 16),
44530 => conv_std_logic_vector(41866, 16),
44531 => conv_std_logic_vector(42039, 16),
44532 => conv_std_logic_vector(42212, 16),
44533 => conv_std_logic_vector(42385, 16),
44534 => conv_std_logic_vector(42558, 16),
44535 => conv_std_logic_vector(42731, 16),
44536 => conv_std_logic_vector(42904, 16),
44537 => conv_std_logic_vector(43077, 16),
44538 => conv_std_logic_vector(43250, 16),
44539 => conv_std_logic_vector(43423, 16),
44540 => conv_std_logic_vector(43596, 16),
44541 => conv_std_logic_vector(43769, 16),
44542 => conv_std_logic_vector(43942, 16),
44543 => conv_std_logic_vector(44115, 16),
44544 => conv_std_logic_vector(0, 16),
44545 => conv_std_logic_vector(174, 16),
44546 => conv_std_logic_vector(348, 16),
44547 => conv_std_logic_vector(522, 16),
44548 => conv_std_logic_vector(696, 16),
44549 => conv_std_logic_vector(870, 16),
44550 => conv_std_logic_vector(1044, 16),
44551 => conv_std_logic_vector(1218, 16),
44552 => conv_std_logic_vector(1392, 16),
44553 => conv_std_logic_vector(1566, 16),
44554 => conv_std_logic_vector(1740, 16),
44555 => conv_std_logic_vector(1914, 16),
44556 => conv_std_logic_vector(2088, 16),
44557 => conv_std_logic_vector(2262, 16),
44558 => conv_std_logic_vector(2436, 16),
44559 => conv_std_logic_vector(2610, 16),
44560 => conv_std_logic_vector(2784, 16),
44561 => conv_std_logic_vector(2958, 16),
44562 => conv_std_logic_vector(3132, 16),
44563 => conv_std_logic_vector(3306, 16),
44564 => conv_std_logic_vector(3480, 16),
44565 => conv_std_logic_vector(3654, 16),
44566 => conv_std_logic_vector(3828, 16),
44567 => conv_std_logic_vector(4002, 16),
44568 => conv_std_logic_vector(4176, 16),
44569 => conv_std_logic_vector(4350, 16),
44570 => conv_std_logic_vector(4524, 16),
44571 => conv_std_logic_vector(4698, 16),
44572 => conv_std_logic_vector(4872, 16),
44573 => conv_std_logic_vector(5046, 16),
44574 => conv_std_logic_vector(5220, 16),
44575 => conv_std_logic_vector(5394, 16),
44576 => conv_std_logic_vector(5568, 16),
44577 => conv_std_logic_vector(5742, 16),
44578 => conv_std_logic_vector(5916, 16),
44579 => conv_std_logic_vector(6090, 16),
44580 => conv_std_logic_vector(6264, 16),
44581 => conv_std_logic_vector(6438, 16),
44582 => conv_std_logic_vector(6612, 16),
44583 => conv_std_logic_vector(6786, 16),
44584 => conv_std_logic_vector(6960, 16),
44585 => conv_std_logic_vector(7134, 16),
44586 => conv_std_logic_vector(7308, 16),
44587 => conv_std_logic_vector(7482, 16),
44588 => conv_std_logic_vector(7656, 16),
44589 => conv_std_logic_vector(7830, 16),
44590 => conv_std_logic_vector(8004, 16),
44591 => conv_std_logic_vector(8178, 16),
44592 => conv_std_logic_vector(8352, 16),
44593 => conv_std_logic_vector(8526, 16),
44594 => conv_std_logic_vector(8700, 16),
44595 => conv_std_logic_vector(8874, 16),
44596 => conv_std_logic_vector(9048, 16),
44597 => conv_std_logic_vector(9222, 16),
44598 => conv_std_logic_vector(9396, 16),
44599 => conv_std_logic_vector(9570, 16),
44600 => conv_std_logic_vector(9744, 16),
44601 => conv_std_logic_vector(9918, 16),
44602 => conv_std_logic_vector(10092, 16),
44603 => conv_std_logic_vector(10266, 16),
44604 => conv_std_logic_vector(10440, 16),
44605 => conv_std_logic_vector(10614, 16),
44606 => conv_std_logic_vector(10788, 16),
44607 => conv_std_logic_vector(10962, 16),
44608 => conv_std_logic_vector(11136, 16),
44609 => conv_std_logic_vector(11310, 16),
44610 => conv_std_logic_vector(11484, 16),
44611 => conv_std_logic_vector(11658, 16),
44612 => conv_std_logic_vector(11832, 16),
44613 => conv_std_logic_vector(12006, 16),
44614 => conv_std_logic_vector(12180, 16),
44615 => conv_std_logic_vector(12354, 16),
44616 => conv_std_logic_vector(12528, 16),
44617 => conv_std_logic_vector(12702, 16),
44618 => conv_std_logic_vector(12876, 16),
44619 => conv_std_logic_vector(13050, 16),
44620 => conv_std_logic_vector(13224, 16),
44621 => conv_std_logic_vector(13398, 16),
44622 => conv_std_logic_vector(13572, 16),
44623 => conv_std_logic_vector(13746, 16),
44624 => conv_std_logic_vector(13920, 16),
44625 => conv_std_logic_vector(14094, 16),
44626 => conv_std_logic_vector(14268, 16),
44627 => conv_std_logic_vector(14442, 16),
44628 => conv_std_logic_vector(14616, 16),
44629 => conv_std_logic_vector(14790, 16),
44630 => conv_std_logic_vector(14964, 16),
44631 => conv_std_logic_vector(15138, 16),
44632 => conv_std_logic_vector(15312, 16),
44633 => conv_std_logic_vector(15486, 16),
44634 => conv_std_logic_vector(15660, 16),
44635 => conv_std_logic_vector(15834, 16),
44636 => conv_std_logic_vector(16008, 16),
44637 => conv_std_logic_vector(16182, 16),
44638 => conv_std_logic_vector(16356, 16),
44639 => conv_std_logic_vector(16530, 16),
44640 => conv_std_logic_vector(16704, 16),
44641 => conv_std_logic_vector(16878, 16),
44642 => conv_std_logic_vector(17052, 16),
44643 => conv_std_logic_vector(17226, 16),
44644 => conv_std_logic_vector(17400, 16),
44645 => conv_std_logic_vector(17574, 16),
44646 => conv_std_logic_vector(17748, 16),
44647 => conv_std_logic_vector(17922, 16),
44648 => conv_std_logic_vector(18096, 16),
44649 => conv_std_logic_vector(18270, 16),
44650 => conv_std_logic_vector(18444, 16),
44651 => conv_std_logic_vector(18618, 16),
44652 => conv_std_logic_vector(18792, 16),
44653 => conv_std_logic_vector(18966, 16),
44654 => conv_std_logic_vector(19140, 16),
44655 => conv_std_logic_vector(19314, 16),
44656 => conv_std_logic_vector(19488, 16),
44657 => conv_std_logic_vector(19662, 16),
44658 => conv_std_logic_vector(19836, 16),
44659 => conv_std_logic_vector(20010, 16),
44660 => conv_std_logic_vector(20184, 16),
44661 => conv_std_logic_vector(20358, 16),
44662 => conv_std_logic_vector(20532, 16),
44663 => conv_std_logic_vector(20706, 16),
44664 => conv_std_logic_vector(20880, 16),
44665 => conv_std_logic_vector(21054, 16),
44666 => conv_std_logic_vector(21228, 16),
44667 => conv_std_logic_vector(21402, 16),
44668 => conv_std_logic_vector(21576, 16),
44669 => conv_std_logic_vector(21750, 16),
44670 => conv_std_logic_vector(21924, 16),
44671 => conv_std_logic_vector(22098, 16),
44672 => conv_std_logic_vector(22272, 16),
44673 => conv_std_logic_vector(22446, 16),
44674 => conv_std_logic_vector(22620, 16),
44675 => conv_std_logic_vector(22794, 16),
44676 => conv_std_logic_vector(22968, 16),
44677 => conv_std_logic_vector(23142, 16),
44678 => conv_std_logic_vector(23316, 16),
44679 => conv_std_logic_vector(23490, 16),
44680 => conv_std_logic_vector(23664, 16),
44681 => conv_std_logic_vector(23838, 16),
44682 => conv_std_logic_vector(24012, 16),
44683 => conv_std_logic_vector(24186, 16),
44684 => conv_std_logic_vector(24360, 16),
44685 => conv_std_logic_vector(24534, 16),
44686 => conv_std_logic_vector(24708, 16),
44687 => conv_std_logic_vector(24882, 16),
44688 => conv_std_logic_vector(25056, 16),
44689 => conv_std_logic_vector(25230, 16),
44690 => conv_std_logic_vector(25404, 16),
44691 => conv_std_logic_vector(25578, 16),
44692 => conv_std_logic_vector(25752, 16),
44693 => conv_std_logic_vector(25926, 16),
44694 => conv_std_logic_vector(26100, 16),
44695 => conv_std_logic_vector(26274, 16),
44696 => conv_std_logic_vector(26448, 16),
44697 => conv_std_logic_vector(26622, 16),
44698 => conv_std_logic_vector(26796, 16),
44699 => conv_std_logic_vector(26970, 16),
44700 => conv_std_logic_vector(27144, 16),
44701 => conv_std_logic_vector(27318, 16),
44702 => conv_std_logic_vector(27492, 16),
44703 => conv_std_logic_vector(27666, 16),
44704 => conv_std_logic_vector(27840, 16),
44705 => conv_std_logic_vector(28014, 16),
44706 => conv_std_logic_vector(28188, 16),
44707 => conv_std_logic_vector(28362, 16),
44708 => conv_std_logic_vector(28536, 16),
44709 => conv_std_logic_vector(28710, 16),
44710 => conv_std_logic_vector(28884, 16),
44711 => conv_std_logic_vector(29058, 16),
44712 => conv_std_logic_vector(29232, 16),
44713 => conv_std_logic_vector(29406, 16),
44714 => conv_std_logic_vector(29580, 16),
44715 => conv_std_logic_vector(29754, 16),
44716 => conv_std_logic_vector(29928, 16),
44717 => conv_std_logic_vector(30102, 16),
44718 => conv_std_logic_vector(30276, 16),
44719 => conv_std_logic_vector(30450, 16),
44720 => conv_std_logic_vector(30624, 16),
44721 => conv_std_logic_vector(30798, 16),
44722 => conv_std_logic_vector(30972, 16),
44723 => conv_std_logic_vector(31146, 16),
44724 => conv_std_logic_vector(31320, 16),
44725 => conv_std_logic_vector(31494, 16),
44726 => conv_std_logic_vector(31668, 16),
44727 => conv_std_logic_vector(31842, 16),
44728 => conv_std_logic_vector(32016, 16),
44729 => conv_std_logic_vector(32190, 16),
44730 => conv_std_logic_vector(32364, 16),
44731 => conv_std_logic_vector(32538, 16),
44732 => conv_std_logic_vector(32712, 16),
44733 => conv_std_logic_vector(32886, 16),
44734 => conv_std_logic_vector(33060, 16),
44735 => conv_std_logic_vector(33234, 16),
44736 => conv_std_logic_vector(33408, 16),
44737 => conv_std_logic_vector(33582, 16),
44738 => conv_std_logic_vector(33756, 16),
44739 => conv_std_logic_vector(33930, 16),
44740 => conv_std_logic_vector(34104, 16),
44741 => conv_std_logic_vector(34278, 16),
44742 => conv_std_logic_vector(34452, 16),
44743 => conv_std_logic_vector(34626, 16),
44744 => conv_std_logic_vector(34800, 16),
44745 => conv_std_logic_vector(34974, 16),
44746 => conv_std_logic_vector(35148, 16),
44747 => conv_std_logic_vector(35322, 16),
44748 => conv_std_logic_vector(35496, 16),
44749 => conv_std_logic_vector(35670, 16),
44750 => conv_std_logic_vector(35844, 16),
44751 => conv_std_logic_vector(36018, 16),
44752 => conv_std_logic_vector(36192, 16),
44753 => conv_std_logic_vector(36366, 16),
44754 => conv_std_logic_vector(36540, 16),
44755 => conv_std_logic_vector(36714, 16),
44756 => conv_std_logic_vector(36888, 16),
44757 => conv_std_logic_vector(37062, 16),
44758 => conv_std_logic_vector(37236, 16),
44759 => conv_std_logic_vector(37410, 16),
44760 => conv_std_logic_vector(37584, 16),
44761 => conv_std_logic_vector(37758, 16),
44762 => conv_std_logic_vector(37932, 16),
44763 => conv_std_logic_vector(38106, 16),
44764 => conv_std_logic_vector(38280, 16),
44765 => conv_std_logic_vector(38454, 16),
44766 => conv_std_logic_vector(38628, 16),
44767 => conv_std_logic_vector(38802, 16),
44768 => conv_std_logic_vector(38976, 16),
44769 => conv_std_logic_vector(39150, 16),
44770 => conv_std_logic_vector(39324, 16),
44771 => conv_std_logic_vector(39498, 16),
44772 => conv_std_logic_vector(39672, 16),
44773 => conv_std_logic_vector(39846, 16),
44774 => conv_std_logic_vector(40020, 16),
44775 => conv_std_logic_vector(40194, 16),
44776 => conv_std_logic_vector(40368, 16),
44777 => conv_std_logic_vector(40542, 16),
44778 => conv_std_logic_vector(40716, 16),
44779 => conv_std_logic_vector(40890, 16),
44780 => conv_std_logic_vector(41064, 16),
44781 => conv_std_logic_vector(41238, 16),
44782 => conv_std_logic_vector(41412, 16),
44783 => conv_std_logic_vector(41586, 16),
44784 => conv_std_logic_vector(41760, 16),
44785 => conv_std_logic_vector(41934, 16),
44786 => conv_std_logic_vector(42108, 16),
44787 => conv_std_logic_vector(42282, 16),
44788 => conv_std_logic_vector(42456, 16),
44789 => conv_std_logic_vector(42630, 16),
44790 => conv_std_logic_vector(42804, 16),
44791 => conv_std_logic_vector(42978, 16),
44792 => conv_std_logic_vector(43152, 16),
44793 => conv_std_logic_vector(43326, 16),
44794 => conv_std_logic_vector(43500, 16),
44795 => conv_std_logic_vector(43674, 16),
44796 => conv_std_logic_vector(43848, 16),
44797 => conv_std_logic_vector(44022, 16),
44798 => conv_std_logic_vector(44196, 16),
44799 => conv_std_logic_vector(44370, 16),
44800 => conv_std_logic_vector(0, 16),
44801 => conv_std_logic_vector(175, 16),
44802 => conv_std_logic_vector(350, 16),
44803 => conv_std_logic_vector(525, 16),
44804 => conv_std_logic_vector(700, 16),
44805 => conv_std_logic_vector(875, 16),
44806 => conv_std_logic_vector(1050, 16),
44807 => conv_std_logic_vector(1225, 16),
44808 => conv_std_logic_vector(1400, 16),
44809 => conv_std_logic_vector(1575, 16),
44810 => conv_std_logic_vector(1750, 16),
44811 => conv_std_logic_vector(1925, 16),
44812 => conv_std_logic_vector(2100, 16),
44813 => conv_std_logic_vector(2275, 16),
44814 => conv_std_logic_vector(2450, 16),
44815 => conv_std_logic_vector(2625, 16),
44816 => conv_std_logic_vector(2800, 16),
44817 => conv_std_logic_vector(2975, 16),
44818 => conv_std_logic_vector(3150, 16),
44819 => conv_std_logic_vector(3325, 16),
44820 => conv_std_logic_vector(3500, 16),
44821 => conv_std_logic_vector(3675, 16),
44822 => conv_std_logic_vector(3850, 16),
44823 => conv_std_logic_vector(4025, 16),
44824 => conv_std_logic_vector(4200, 16),
44825 => conv_std_logic_vector(4375, 16),
44826 => conv_std_logic_vector(4550, 16),
44827 => conv_std_logic_vector(4725, 16),
44828 => conv_std_logic_vector(4900, 16),
44829 => conv_std_logic_vector(5075, 16),
44830 => conv_std_logic_vector(5250, 16),
44831 => conv_std_logic_vector(5425, 16),
44832 => conv_std_logic_vector(5600, 16),
44833 => conv_std_logic_vector(5775, 16),
44834 => conv_std_logic_vector(5950, 16),
44835 => conv_std_logic_vector(6125, 16),
44836 => conv_std_logic_vector(6300, 16),
44837 => conv_std_logic_vector(6475, 16),
44838 => conv_std_logic_vector(6650, 16),
44839 => conv_std_logic_vector(6825, 16),
44840 => conv_std_logic_vector(7000, 16),
44841 => conv_std_logic_vector(7175, 16),
44842 => conv_std_logic_vector(7350, 16),
44843 => conv_std_logic_vector(7525, 16),
44844 => conv_std_logic_vector(7700, 16),
44845 => conv_std_logic_vector(7875, 16),
44846 => conv_std_logic_vector(8050, 16),
44847 => conv_std_logic_vector(8225, 16),
44848 => conv_std_logic_vector(8400, 16),
44849 => conv_std_logic_vector(8575, 16),
44850 => conv_std_logic_vector(8750, 16),
44851 => conv_std_logic_vector(8925, 16),
44852 => conv_std_logic_vector(9100, 16),
44853 => conv_std_logic_vector(9275, 16),
44854 => conv_std_logic_vector(9450, 16),
44855 => conv_std_logic_vector(9625, 16),
44856 => conv_std_logic_vector(9800, 16),
44857 => conv_std_logic_vector(9975, 16),
44858 => conv_std_logic_vector(10150, 16),
44859 => conv_std_logic_vector(10325, 16),
44860 => conv_std_logic_vector(10500, 16),
44861 => conv_std_logic_vector(10675, 16),
44862 => conv_std_logic_vector(10850, 16),
44863 => conv_std_logic_vector(11025, 16),
44864 => conv_std_logic_vector(11200, 16),
44865 => conv_std_logic_vector(11375, 16),
44866 => conv_std_logic_vector(11550, 16),
44867 => conv_std_logic_vector(11725, 16),
44868 => conv_std_logic_vector(11900, 16),
44869 => conv_std_logic_vector(12075, 16),
44870 => conv_std_logic_vector(12250, 16),
44871 => conv_std_logic_vector(12425, 16),
44872 => conv_std_logic_vector(12600, 16),
44873 => conv_std_logic_vector(12775, 16),
44874 => conv_std_logic_vector(12950, 16),
44875 => conv_std_logic_vector(13125, 16),
44876 => conv_std_logic_vector(13300, 16),
44877 => conv_std_logic_vector(13475, 16),
44878 => conv_std_logic_vector(13650, 16),
44879 => conv_std_logic_vector(13825, 16),
44880 => conv_std_logic_vector(14000, 16),
44881 => conv_std_logic_vector(14175, 16),
44882 => conv_std_logic_vector(14350, 16),
44883 => conv_std_logic_vector(14525, 16),
44884 => conv_std_logic_vector(14700, 16),
44885 => conv_std_logic_vector(14875, 16),
44886 => conv_std_logic_vector(15050, 16),
44887 => conv_std_logic_vector(15225, 16),
44888 => conv_std_logic_vector(15400, 16),
44889 => conv_std_logic_vector(15575, 16),
44890 => conv_std_logic_vector(15750, 16),
44891 => conv_std_logic_vector(15925, 16),
44892 => conv_std_logic_vector(16100, 16),
44893 => conv_std_logic_vector(16275, 16),
44894 => conv_std_logic_vector(16450, 16),
44895 => conv_std_logic_vector(16625, 16),
44896 => conv_std_logic_vector(16800, 16),
44897 => conv_std_logic_vector(16975, 16),
44898 => conv_std_logic_vector(17150, 16),
44899 => conv_std_logic_vector(17325, 16),
44900 => conv_std_logic_vector(17500, 16),
44901 => conv_std_logic_vector(17675, 16),
44902 => conv_std_logic_vector(17850, 16),
44903 => conv_std_logic_vector(18025, 16),
44904 => conv_std_logic_vector(18200, 16),
44905 => conv_std_logic_vector(18375, 16),
44906 => conv_std_logic_vector(18550, 16),
44907 => conv_std_logic_vector(18725, 16),
44908 => conv_std_logic_vector(18900, 16),
44909 => conv_std_logic_vector(19075, 16),
44910 => conv_std_logic_vector(19250, 16),
44911 => conv_std_logic_vector(19425, 16),
44912 => conv_std_logic_vector(19600, 16),
44913 => conv_std_logic_vector(19775, 16),
44914 => conv_std_logic_vector(19950, 16),
44915 => conv_std_logic_vector(20125, 16),
44916 => conv_std_logic_vector(20300, 16),
44917 => conv_std_logic_vector(20475, 16),
44918 => conv_std_logic_vector(20650, 16),
44919 => conv_std_logic_vector(20825, 16),
44920 => conv_std_logic_vector(21000, 16),
44921 => conv_std_logic_vector(21175, 16),
44922 => conv_std_logic_vector(21350, 16),
44923 => conv_std_logic_vector(21525, 16),
44924 => conv_std_logic_vector(21700, 16),
44925 => conv_std_logic_vector(21875, 16),
44926 => conv_std_logic_vector(22050, 16),
44927 => conv_std_logic_vector(22225, 16),
44928 => conv_std_logic_vector(22400, 16),
44929 => conv_std_logic_vector(22575, 16),
44930 => conv_std_logic_vector(22750, 16),
44931 => conv_std_logic_vector(22925, 16),
44932 => conv_std_logic_vector(23100, 16),
44933 => conv_std_logic_vector(23275, 16),
44934 => conv_std_logic_vector(23450, 16),
44935 => conv_std_logic_vector(23625, 16),
44936 => conv_std_logic_vector(23800, 16),
44937 => conv_std_logic_vector(23975, 16),
44938 => conv_std_logic_vector(24150, 16),
44939 => conv_std_logic_vector(24325, 16),
44940 => conv_std_logic_vector(24500, 16),
44941 => conv_std_logic_vector(24675, 16),
44942 => conv_std_logic_vector(24850, 16),
44943 => conv_std_logic_vector(25025, 16),
44944 => conv_std_logic_vector(25200, 16),
44945 => conv_std_logic_vector(25375, 16),
44946 => conv_std_logic_vector(25550, 16),
44947 => conv_std_logic_vector(25725, 16),
44948 => conv_std_logic_vector(25900, 16),
44949 => conv_std_logic_vector(26075, 16),
44950 => conv_std_logic_vector(26250, 16),
44951 => conv_std_logic_vector(26425, 16),
44952 => conv_std_logic_vector(26600, 16),
44953 => conv_std_logic_vector(26775, 16),
44954 => conv_std_logic_vector(26950, 16),
44955 => conv_std_logic_vector(27125, 16),
44956 => conv_std_logic_vector(27300, 16),
44957 => conv_std_logic_vector(27475, 16),
44958 => conv_std_logic_vector(27650, 16),
44959 => conv_std_logic_vector(27825, 16),
44960 => conv_std_logic_vector(28000, 16),
44961 => conv_std_logic_vector(28175, 16),
44962 => conv_std_logic_vector(28350, 16),
44963 => conv_std_logic_vector(28525, 16),
44964 => conv_std_logic_vector(28700, 16),
44965 => conv_std_logic_vector(28875, 16),
44966 => conv_std_logic_vector(29050, 16),
44967 => conv_std_logic_vector(29225, 16),
44968 => conv_std_logic_vector(29400, 16),
44969 => conv_std_logic_vector(29575, 16),
44970 => conv_std_logic_vector(29750, 16),
44971 => conv_std_logic_vector(29925, 16),
44972 => conv_std_logic_vector(30100, 16),
44973 => conv_std_logic_vector(30275, 16),
44974 => conv_std_logic_vector(30450, 16),
44975 => conv_std_logic_vector(30625, 16),
44976 => conv_std_logic_vector(30800, 16),
44977 => conv_std_logic_vector(30975, 16),
44978 => conv_std_logic_vector(31150, 16),
44979 => conv_std_logic_vector(31325, 16),
44980 => conv_std_logic_vector(31500, 16),
44981 => conv_std_logic_vector(31675, 16),
44982 => conv_std_logic_vector(31850, 16),
44983 => conv_std_logic_vector(32025, 16),
44984 => conv_std_logic_vector(32200, 16),
44985 => conv_std_logic_vector(32375, 16),
44986 => conv_std_logic_vector(32550, 16),
44987 => conv_std_logic_vector(32725, 16),
44988 => conv_std_logic_vector(32900, 16),
44989 => conv_std_logic_vector(33075, 16),
44990 => conv_std_logic_vector(33250, 16),
44991 => conv_std_logic_vector(33425, 16),
44992 => conv_std_logic_vector(33600, 16),
44993 => conv_std_logic_vector(33775, 16),
44994 => conv_std_logic_vector(33950, 16),
44995 => conv_std_logic_vector(34125, 16),
44996 => conv_std_logic_vector(34300, 16),
44997 => conv_std_logic_vector(34475, 16),
44998 => conv_std_logic_vector(34650, 16),
44999 => conv_std_logic_vector(34825, 16),
45000 => conv_std_logic_vector(35000, 16),
45001 => conv_std_logic_vector(35175, 16),
45002 => conv_std_logic_vector(35350, 16),
45003 => conv_std_logic_vector(35525, 16),
45004 => conv_std_logic_vector(35700, 16),
45005 => conv_std_logic_vector(35875, 16),
45006 => conv_std_logic_vector(36050, 16),
45007 => conv_std_logic_vector(36225, 16),
45008 => conv_std_logic_vector(36400, 16),
45009 => conv_std_logic_vector(36575, 16),
45010 => conv_std_logic_vector(36750, 16),
45011 => conv_std_logic_vector(36925, 16),
45012 => conv_std_logic_vector(37100, 16),
45013 => conv_std_logic_vector(37275, 16),
45014 => conv_std_logic_vector(37450, 16),
45015 => conv_std_logic_vector(37625, 16),
45016 => conv_std_logic_vector(37800, 16),
45017 => conv_std_logic_vector(37975, 16),
45018 => conv_std_logic_vector(38150, 16),
45019 => conv_std_logic_vector(38325, 16),
45020 => conv_std_logic_vector(38500, 16),
45021 => conv_std_logic_vector(38675, 16),
45022 => conv_std_logic_vector(38850, 16),
45023 => conv_std_logic_vector(39025, 16),
45024 => conv_std_logic_vector(39200, 16),
45025 => conv_std_logic_vector(39375, 16),
45026 => conv_std_logic_vector(39550, 16),
45027 => conv_std_logic_vector(39725, 16),
45028 => conv_std_logic_vector(39900, 16),
45029 => conv_std_logic_vector(40075, 16),
45030 => conv_std_logic_vector(40250, 16),
45031 => conv_std_logic_vector(40425, 16),
45032 => conv_std_logic_vector(40600, 16),
45033 => conv_std_logic_vector(40775, 16),
45034 => conv_std_logic_vector(40950, 16),
45035 => conv_std_logic_vector(41125, 16),
45036 => conv_std_logic_vector(41300, 16),
45037 => conv_std_logic_vector(41475, 16),
45038 => conv_std_logic_vector(41650, 16),
45039 => conv_std_logic_vector(41825, 16),
45040 => conv_std_logic_vector(42000, 16),
45041 => conv_std_logic_vector(42175, 16),
45042 => conv_std_logic_vector(42350, 16),
45043 => conv_std_logic_vector(42525, 16),
45044 => conv_std_logic_vector(42700, 16),
45045 => conv_std_logic_vector(42875, 16),
45046 => conv_std_logic_vector(43050, 16),
45047 => conv_std_logic_vector(43225, 16),
45048 => conv_std_logic_vector(43400, 16),
45049 => conv_std_logic_vector(43575, 16),
45050 => conv_std_logic_vector(43750, 16),
45051 => conv_std_logic_vector(43925, 16),
45052 => conv_std_logic_vector(44100, 16),
45053 => conv_std_logic_vector(44275, 16),
45054 => conv_std_logic_vector(44450, 16),
45055 => conv_std_logic_vector(44625, 16),
45056 => conv_std_logic_vector(0, 16),
45057 => conv_std_logic_vector(176, 16),
45058 => conv_std_logic_vector(352, 16),
45059 => conv_std_logic_vector(528, 16),
45060 => conv_std_logic_vector(704, 16),
45061 => conv_std_logic_vector(880, 16),
45062 => conv_std_logic_vector(1056, 16),
45063 => conv_std_logic_vector(1232, 16),
45064 => conv_std_logic_vector(1408, 16),
45065 => conv_std_logic_vector(1584, 16),
45066 => conv_std_logic_vector(1760, 16),
45067 => conv_std_logic_vector(1936, 16),
45068 => conv_std_logic_vector(2112, 16),
45069 => conv_std_logic_vector(2288, 16),
45070 => conv_std_logic_vector(2464, 16),
45071 => conv_std_logic_vector(2640, 16),
45072 => conv_std_logic_vector(2816, 16),
45073 => conv_std_logic_vector(2992, 16),
45074 => conv_std_logic_vector(3168, 16),
45075 => conv_std_logic_vector(3344, 16),
45076 => conv_std_logic_vector(3520, 16),
45077 => conv_std_logic_vector(3696, 16),
45078 => conv_std_logic_vector(3872, 16),
45079 => conv_std_logic_vector(4048, 16),
45080 => conv_std_logic_vector(4224, 16),
45081 => conv_std_logic_vector(4400, 16),
45082 => conv_std_logic_vector(4576, 16),
45083 => conv_std_logic_vector(4752, 16),
45084 => conv_std_logic_vector(4928, 16),
45085 => conv_std_logic_vector(5104, 16),
45086 => conv_std_logic_vector(5280, 16),
45087 => conv_std_logic_vector(5456, 16),
45088 => conv_std_logic_vector(5632, 16),
45089 => conv_std_logic_vector(5808, 16),
45090 => conv_std_logic_vector(5984, 16),
45091 => conv_std_logic_vector(6160, 16),
45092 => conv_std_logic_vector(6336, 16),
45093 => conv_std_logic_vector(6512, 16),
45094 => conv_std_logic_vector(6688, 16),
45095 => conv_std_logic_vector(6864, 16),
45096 => conv_std_logic_vector(7040, 16),
45097 => conv_std_logic_vector(7216, 16),
45098 => conv_std_logic_vector(7392, 16),
45099 => conv_std_logic_vector(7568, 16),
45100 => conv_std_logic_vector(7744, 16),
45101 => conv_std_logic_vector(7920, 16),
45102 => conv_std_logic_vector(8096, 16),
45103 => conv_std_logic_vector(8272, 16),
45104 => conv_std_logic_vector(8448, 16),
45105 => conv_std_logic_vector(8624, 16),
45106 => conv_std_logic_vector(8800, 16),
45107 => conv_std_logic_vector(8976, 16),
45108 => conv_std_logic_vector(9152, 16),
45109 => conv_std_logic_vector(9328, 16),
45110 => conv_std_logic_vector(9504, 16),
45111 => conv_std_logic_vector(9680, 16),
45112 => conv_std_logic_vector(9856, 16),
45113 => conv_std_logic_vector(10032, 16),
45114 => conv_std_logic_vector(10208, 16),
45115 => conv_std_logic_vector(10384, 16),
45116 => conv_std_logic_vector(10560, 16),
45117 => conv_std_logic_vector(10736, 16),
45118 => conv_std_logic_vector(10912, 16),
45119 => conv_std_logic_vector(11088, 16),
45120 => conv_std_logic_vector(11264, 16),
45121 => conv_std_logic_vector(11440, 16),
45122 => conv_std_logic_vector(11616, 16),
45123 => conv_std_logic_vector(11792, 16),
45124 => conv_std_logic_vector(11968, 16),
45125 => conv_std_logic_vector(12144, 16),
45126 => conv_std_logic_vector(12320, 16),
45127 => conv_std_logic_vector(12496, 16),
45128 => conv_std_logic_vector(12672, 16),
45129 => conv_std_logic_vector(12848, 16),
45130 => conv_std_logic_vector(13024, 16),
45131 => conv_std_logic_vector(13200, 16),
45132 => conv_std_logic_vector(13376, 16),
45133 => conv_std_logic_vector(13552, 16),
45134 => conv_std_logic_vector(13728, 16),
45135 => conv_std_logic_vector(13904, 16),
45136 => conv_std_logic_vector(14080, 16),
45137 => conv_std_logic_vector(14256, 16),
45138 => conv_std_logic_vector(14432, 16),
45139 => conv_std_logic_vector(14608, 16),
45140 => conv_std_logic_vector(14784, 16),
45141 => conv_std_logic_vector(14960, 16),
45142 => conv_std_logic_vector(15136, 16),
45143 => conv_std_logic_vector(15312, 16),
45144 => conv_std_logic_vector(15488, 16),
45145 => conv_std_logic_vector(15664, 16),
45146 => conv_std_logic_vector(15840, 16),
45147 => conv_std_logic_vector(16016, 16),
45148 => conv_std_logic_vector(16192, 16),
45149 => conv_std_logic_vector(16368, 16),
45150 => conv_std_logic_vector(16544, 16),
45151 => conv_std_logic_vector(16720, 16),
45152 => conv_std_logic_vector(16896, 16),
45153 => conv_std_logic_vector(17072, 16),
45154 => conv_std_logic_vector(17248, 16),
45155 => conv_std_logic_vector(17424, 16),
45156 => conv_std_logic_vector(17600, 16),
45157 => conv_std_logic_vector(17776, 16),
45158 => conv_std_logic_vector(17952, 16),
45159 => conv_std_logic_vector(18128, 16),
45160 => conv_std_logic_vector(18304, 16),
45161 => conv_std_logic_vector(18480, 16),
45162 => conv_std_logic_vector(18656, 16),
45163 => conv_std_logic_vector(18832, 16),
45164 => conv_std_logic_vector(19008, 16),
45165 => conv_std_logic_vector(19184, 16),
45166 => conv_std_logic_vector(19360, 16),
45167 => conv_std_logic_vector(19536, 16),
45168 => conv_std_logic_vector(19712, 16),
45169 => conv_std_logic_vector(19888, 16),
45170 => conv_std_logic_vector(20064, 16),
45171 => conv_std_logic_vector(20240, 16),
45172 => conv_std_logic_vector(20416, 16),
45173 => conv_std_logic_vector(20592, 16),
45174 => conv_std_logic_vector(20768, 16),
45175 => conv_std_logic_vector(20944, 16),
45176 => conv_std_logic_vector(21120, 16),
45177 => conv_std_logic_vector(21296, 16),
45178 => conv_std_logic_vector(21472, 16),
45179 => conv_std_logic_vector(21648, 16),
45180 => conv_std_logic_vector(21824, 16),
45181 => conv_std_logic_vector(22000, 16),
45182 => conv_std_logic_vector(22176, 16),
45183 => conv_std_logic_vector(22352, 16),
45184 => conv_std_logic_vector(22528, 16),
45185 => conv_std_logic_vector(22704, 16),
45186 => conv_std_logic_vector(22880, 16),
45187 => conv_std_logic_vector(23056, 16),
45188 => conv_std_logic_vector(23232, 16),
45189 => conv_std_logic_vector(23408, 16),
45190 => conv_std_logic_vector(23584, 16),
45191 => conv_std_logic_vector(23760, 16),
45192 => conv_std_logic_vector(23936, 16),
45193 => conv_std_logic_vector(24112, 16),
45194 => conv_std_logic_vector(24288, 16),
45195 => conv_std_logic_vector(24464, 16),
45196 => conv_std_logic_vector(24640, 16),
45197 => conv_std_logic_vector(24816, 16),
45198 => conv_std_logic_vector(24992, 16),
45199 => conv_std_logic_vector(25168, 16),
45200 => conv_std_logic_vector(25344, 16),
45201 => conv_std_logic_vector(25520, 16),
45202 => conv_std_logic_vector(25696, 16),
45203 => conv_std_logic_vector(25872, 16),
45204 => conv_std_logic_vector(26048, 16),
45205 => conv_std_logic_vector(26224, 16),
45206 => conv_std_logic_vector(26400, 16),
45207 => conv_std_logic_vector(26576, 16),
45208 => conv_std_logic_vector(26752, 16),
45209 => conv_std_logic_vector(26928, 16),
45210 => conv_std_logic_vector(27104, 16),
45211 => conv_std_logic_vector(27280, 16),
45212 => conv_std_logic_vector(27456, 16),
45213 => conv_std_logic_vector(27632, 16),
45214 => conv_std_logic_vector(27808, 16),
45215 => conv_std_logic_vector(27984, 16),
45216 => conv_std_logic_vector(28160, 16),
45217 => conv_std_logic_vector(28336, 16),
45218 => conv_std_logic_vector(28512, 16),
45219 => conv_std_logic_vector(28688, 16),
45220 => conv_std_logic_vector(28864, 16),
45221 => conv_std_logic_vector(29040, 16),
45222 => conv_std_logic_vector(29216, 16),
45223 => conv_std_logic_vector(29392, 16),
45224 => conv_std_logic_vector(29568, 16),
45225 => conv_std_logic_vector(29744, 16),
45226 => conv_std_logic_vector(29920, 16),
45227 => conv_std_logic_vector(30096, 16),
45228 => conv_std_logic_vector(30272, 16),
45229 => conv_std_logic_vector(30448, 16),
45230 => conv_std_logic_vector(30624, 16),
45231 => conv_std_logic_vector(30800, 16),
45232 => conv_std_logic_vector(30976, 16),
45233 => conv_std_logic_vector(31152, 16),
45234 => conv_std_logic_vector(31328, 16),
45235 => conv_std_logic_vector(31504, 16),
45236 => conv_std_logic_vector(31680, 16),
45237 => conv_std_logic_vector(31856, 16),
45238 => conv_std_logic_vector(32032, 16),
45239 => conv_std_logic_vector(32208, 16),
45240 => conv_std_logic_vector(32384, 16),
45241 => conv_std_logic_vector(32560, 16),
45242 => conv_std_logic_vector(32736, 16),
45243 => conv_std_logic_vector(32912, 16),
45244 => conv_std_logic_vector(33088, 16),
45245 => conv_std_logic_vector(33264, 16),
45246 => conv_std_logic_vector(33440, 16),
45247 => conv_std_logic_vector(33616, 16),
45248 => conv_std_logic_vector(33792, 16),
45249 => conv_std_logic_vector(33968, 16),
45250 => conv_std_logic_vector(34144, 16),
45251 => conv_std_logic_vector(34320, 16),
45252 => conv_std_logic_vector(34496, 16),
45253 => conv_std_logic_vector(34672, 16),
45254 => conv_std_logic_vector(34848, 16),
45255 => conv_std_logic_vector(35024, 16),
45256 => conv_std_logic_vector(35200, 16),
45257 => conv_std_logic_vector(35376, 16),
45258 => conv_std_logic_vector(35552, 16),
45259 => conv_std_logic_vector(35728, 16),
45260 => conv_std_logic_vector(35904, 16),
45261 => conv_std_logic_vector(36080, 16),
45262 => conv_std_logic_vector(36256, 16),
45263 => conv_std_logic_vector(36432, 16),
45264 => conv_std_logic_vector(36608, 16),
45265 => conv_std_logic_vector(36784, 16),
45266 => conv_std_logic_vector(36960, 16),
45267 => conv_std_logic_vector(37136, 16),
45268 => conv_std_logic_vector(37312, 16),
45269 => conv_std_logic_vector(37488, 16),
45270 => conv_std_logic_vector(37664, 16),
45271 => conv_std_logic_vector(37840, 16),
45272 => conv_std_logic_vector(38016, 16),
45273 => conv_std_logic_vector(38192, 16),
45274 => conv_std_logic_vector(38368, 16),
45275 => conv_std_logic_vector(38544, 16),
45276 => conv_std_logic_vector(38720, 16),
45277 => conv_std_logic_vector(38896, 16),
45278 => conv_std_logic_vector(39072, 16),
45279 => conv_std_logic_vector(39248, 16),
45280 => conv_std_logic_vector(39424, 16),
45281 => conv_std_logic_vector(39600, 16),
45282 => conv_std_logic_vector(39776, 16),
45283 => conv_std_logic_vector(39952, 16),
45284 => conv_std_logic_vector(40128, 16),
45285 => conv_std_logic_vector(40304, 16),
45286 => conv_std_logic_vector(40480, 16),
45287 => conv_std_logic_vector(40656, 16),
45288 => conv_std_logic_vector(40832, 16),
45289 => conv_std_logic_vector(41008, 16),
45290 => conv_std_logic_vector(41184, 16),
45291 => conv_std_logic_vector(41360, 16),
45292 => conv_std_logic_vector(41536, 16),
45293 => conv_std_logic_vector(41712, 16),
45294 => conv_std_logic_vector(41888, 16),
45295 => conv_std_logic_vector(42064, 16),
45296 => conv_std_logic_vector(42240, 16),
45297 => conv_std_logic_vector(42416, 16),
45298 => conv_std_logic_vector(42592, 16),
45299 => conv_std_logic_vector(42768, 16),
45300 => conv_std_logic_vector(42944, 16),
45301 => conv_std_logic_vector(43120, 16),
45302 => conv_std_logic_vector(43296, 16),
45303 => conv_std_logic_vector(43472, 16),
45304 => conv_std_logic_vector(43648, 16),
45305 => conv_std_logic_vector(43824, 16),
45306 => conv_std_logic_vector(44000, 16),
45307 => conv_std_logic_vector(44176, 16),
45308 => conv_std_logic_vector(44352, 16),
45309 => conv_std_logic_vector(44528, 16),
45310 => conv_std_logic_vector(44704, 16),
45311 => conv_std_logic_vector(44880, 16),
45312 => conv_std_logic_vector(0, 16),
45313 => conv_std_logic_vector(177, 16),
45314 => conv_std_logic_vector(354, 16),
45315 => conv_std_logic_vector(531, 16),
45316 => conv_std_logic_vector(708, 16),
45317 => conv_std_logic_vector(885, 16),
45318 => conv_std_logic_vector(1062, 16),
45319 => conv_std_logic_vector(1239, 16),
45320 => conv_std_logic_vector(1416, 16),
45321 => conv_std_logic_vector(1593, 16),
45322 => conv_std_logic_vector(1770, 16),
45323 => conv_std_logic_vector(1947, 16),
45324 => conv_std_logic_vector(2124, 16),
45325 => conv_std_logic_vector(2301, 16),
45326 => conv_std_logic_vector(2478, 16),
45327 => conv_std_logic_vector(2655, 16),
45328 => conv_std_logic_vector(2832, 16),
45329 => conv_std_logic_vector(3009, 16),
45330 => conv_std_logic_vector(3186, 16),
45331 => conv_std_logic_vector(3363, 16),
45332 => conv_std_logic_vector(3540, 16),
45333 => conv_std_logic_vector(3717, 16),
45334 => conv_std_logic_vector(3894, 16),
45335 => conv_std_logic_vector(4071, 16),
45336 => conv_std_logic_vector(4248, 16),
45337 => conv_std_logic_vector(4425, 16),
45338 => conv_std_logic_vector(4602, 16),
45339 => conv_std_logic_vector(4779, 16),
45340 => conv_std_logic_vector(4956, 16),
45341 => conv_std_logic_vector(5133, 16),
45342 => conv_std_logic_vector(5310, 16),
45343 => conv_std_logic_vector(5487, 16),
45344 => conv_std_logic_vector(5664, 16),
45345 => conv_std_logic_vector(5841, 16),
45346 => conv_std_logic_vector(6018, 16),
45347 => conv_std_logic_vector(6195, 16),
45348 => conv_std_logic_vector(6372, 16),
45349 => conv_std_logic_vector(6549, 16),
45350 => conv_std_logic_vector(6726, 16),
45351 => conv_std_logic_vector(6903, 16),
45352 => conv_std_logic_vector(7080, 16),
45353 => conv_std_logic_vector(7257, 16),
45354 => conv_std_logic_vector(7434, 16),
45355 => conv_std_logic_vector(7611, 16),
45356 => conv_std_logic_vector(7788, 16),
45357 => conv_std_logic_vector(7965, 16),
45358 => conv_std_logic_vector(8142, 16),
45359 => conv_std_logic_vector(8319, 16),
45360 => conv_std_logic_vector(8496, 16),
45361 => conv_std_logic_vector(8673, 16),
45362 => conv_std_logic_vector(8850, 16),
45363 => conv_std_logic_vector(9027, 16),
45364 => conv_std_logic_vector(9204, 16),
45365 => conv_std_logic_vector(9381, 16),
45366 => conv_std_logic_vector(9558, 16),
45367 => conv_std_logic_vector(9735, 16),
45368 => conv_std_logic_vector(9912, 16),
45369 => conv_std_logic_vector(10089, 16),
45370 => conv_std_logic_vector(10266, 16),
45371 => conv_std_logic_vector(10443, 16),
45372 => conv_std_logic_vector(10620, 16),
45373 => conv_std_logic_vector(10797, 16),
45374 => conv_std_logic_vector(10974, 16),
45375 => conv_std_logic_vector(11151, 16),
45376 => conv_std_logic_vector(11328, 16),
45377 => conv_std_logic_vector(11505, 16),
45378 => conv_std_logic_vector(11682, 16),
45379 => conv_std_logic_vector(11859, 16),
45380 => conv_std_logic_vector(12036, 16),
45381 => conv_std_logic_vector(12213, 16),
45382 => conv_std_logic_vector(12390, 16),
45383 => conv_std_logic_vector(12567, 16),
45384 => conv_std_logic_vector(12744, 16),
45385 => conv_std_logic_vector(12921, 16),
45386 => conv_std_logic_vector(13098, 16),
45387 => conv_std_logic_vector(13275, 16),
45388 => conv_std_logic_vector(13452, 16),
45389 => conv_std_logic_vector(13629, 16),
45390 => conv_std_logic_vector(13806, 16),
45391 => conv_std_logic_vector(13983, 16),
45392 => conv_std_logic_vector(14160, 16),
45393 => conv_std_logic_vector(14337, 16),
45394 => conv_std_logic_vector(14514, 16),
45395 => conv_std_logic_vector(14691, 16),
45396 => conv_std_logic_vector(14868, 16),
45397 => conv_std_logic_vector(15045, 16),
45398 => conv_std_logic_vector(15222, 16),
45399 => conv_std_logic_vector(15399, 16),
45400 => conv_std_logic_vector(15576, 16),
45401 => conv_std_logic_vector(15753, 16),
45402 => conv_std_logic_vector(15930, 16),
45403 => conv_std_logic_vector(16107, 16),
45404 => conv_std_logic_vector(16284, 16),
45405 => conv_std_logic_vector(16461, 16),
45406 => conv_std_logic_vector(16638, 16),
45407 => conv_std_logic_vector(16815, 16),
45408 => conv_std_logic_vector(16992, 16),
45409 => conv_std_logic_vector(17169, 16),
45410 => conv_std_logic_vector(17346, 16),
45411 => conv_std_logic_vector(17523, 16),
45412 => conv_std_logic_vector(17700, 16),
45413 => conv_std_logic_vector(17877, 16),
45414 => conv_std_logic_vector(18054, 16),
45415 => conv_std_logic_vector(18231, 16),
45416 => conv_std_logic_vector(18408, 16),
45417 => conv_std_logic_vector(18585, 16),
45418 => conv_std_logic_vector(18762, 16),
45419 => conv_std_logic_vector(18939, 16),
45420 => conv_std_logic_vector(19116, 16),
45421 => conv_std_logic_vector(19293, 16),
45422 => conv_std_logic_vector(19470, 16),
45423 => conv_std_logic_vector(19647, 16),
45424 => conv_std_logic_vector(19824, 16),
45425 => conv_std_logic_vector(20001, 16),
45426 => conv_std_logic_vector(20178, 16),
45427 => conv_std_logic_vector(20355, 16),
45428 => conv_std_logic_vector(20532, 16),
45429 => conv_std_logic_vector(20709, 16),
45430 => conv_std_logic_vector(20886, 16),
45431 => conv_std_logic_vector(21063, 16),
45432 => conv_std_logic_vector(21240, 16),
45433 => conv_std_logic_vector(21417, 16),
45434 => conv_std_logic_vector(21594, 16),
45435 => conv_std_logic_vector(21771, 16),
45436 => conv_std_logic_vector(21948, 16),
45437 => conv_std_logic_vector(22125, 16),
45438 => conv_std_logic_vector(22302, 16),
45439 => conv_std_logic_vector(22479, 16),
45440 => conv_std_logic_vector(22656, 16),
45441 => conv_std_logic_vector(22833, 16),
45442 => conv_std_logic_vector(23010, 16),
45443 => conv_std_logic_vector(23187, 16),
45444 => conv_std_logic_vector(23364, 16),
45445 => conv_std_logic_vector(23541, 16),
45446 => conv_std_logic_vector(23718, 16),
45447 => conv_std_logic_vector(23895, 16),
45448 => conv_std_logic_vector(24072, 16),
45449 => conv_std_logic_vector(24249, 16),
45450 => conv_std_logic_vector(24426, 16),
45451 => conv_std_logic_vector(24603, 16),
45452 => conv_std_logic_vector(24780, 16),
45453 => conv_std_logic_vector(24957, 16),
45454 => conv_std_logic_vector(25134, 16),
45455 => conv_std_logic_vector(25311, 16),
45456 => conv_std_logic_vector(25488, 16),
45457 => conv_std_logic_vector(25665, 16),
45458 => conv_std_logic_vector(25842, 16),
45459 => conv_std_logic_vector(26019, 16),
45460 => conv_std_logic_vector(26196, 16),
45461 => conv_std_logic_vector(26373, 16),
45462 => conv_std_logic_vector(26550, 16),
45463 => conv_std_logic_vector(26727, 16),
45464 => conv_std_logic_vector(26904, 16),
45465 => conv_std_logic_vector(27081, 16),
45466 => conv_std_logic_vector(27258, 16),
45467 => conv_std_logic_vector(27435, 16),
45468 => conv_std_logic_vector(27612, 16),
45469 => conv_std_logic_vector(27789, 16),
45470 => conv_std_logic_vector(27966, 16),
45471 => conv_std_logic_vector(28143, 16),
45472 => conv_std_logic_vector(28320, 16),
45473 => conv_std_logic_vector(28497, 16),
45474 => conv_std_logic_vector(28674, 16),
45475 => conv_std_logic_vector(28851, 16),
45476 => conv_std_logic_vector(29028, 16),
45477 => conv_std_logic_vector(29205, 16),
45478 => conv_std_logic_vector(29382, 16),
45479 => conv_std_logic_vector(29559, 16),
45480 => conv_std_logic_vector(29736, 16),
45481 => conv_std_logic_vector(29913, 16),
45482 => conv_std_logic_vector(30090, 16),
45483 => conv_std_logic_vector(30267, 16),
45484 => conv_std_logic_vector(30444, 16),
45485 => conv_std_logic_vector(30621, 16),
45486 => conv_std_logic_vector(30798, 16),
45487 => conv_std_logic_vector(30975, 16),
45488 => conv_std_logic_vector(31152, 16),
45489 => conv_std_logic_vector(31329, 16),
45490 => conv_std_logic_vector(31506, 16),
45491 => conv_std_logic_vector(31683, 16),
45492 => conv_std_logic_vector(31860, 16),
45493 => conv_std_logic_vector(32037, 16),
45494 => conv_std_logic_vector(32214, 16),
45495 => conv_std_logic_vector(32391, 16),
45496 => conv_std_logic_vector(32568, 16),
45497 => conv_std_logic_vector(32745, 16),
45498 => conv_std_logic_vector(32922, 16),
45499 => conv_std_logic_vector(33099, 16),
45500 => conv_std_logic_vector(33276, 16),
45501 => conv_std_logic_vector(33453, 16),
45502 => conv_std_logic_vector(33630, 16),
45503 => conv_std_logic_vector(33807, 16),
45504 => conv_std_logic_vector(33984, 16),
45505 => conv_std_logic_vector(34161, 16),
45506 => conv_std_logic_vector(34338, 16),
45507 => conv_std_logic_vector(34515, 16),
45508 => conv_std_logic_vector(34692, 16),
45509 => conv_std_logic_vector(34869, 16),
45510 => conv_std_logic_vector(35046, 16),
45511 => conv_std_logic_vector(35223, 16),
45512 => conv_std_logic_vector(35400, 16),
45513 => conv_std_logic_vector(35577, 16),
45514 => conv_std_logic_vector(35754, 16),
45515 => conv_std_logic_vector(35931, 16),
45516 => conv_std_logic_vector(36108, 16),
45517 => conv_std_logic_vector(36285, 16),
45518 => conv_std_logic_vector(36462, 16),
45519 => conv_std_logic_vector(36639, 16),
45520 => conv_std_logic_vector(36816, 16),
45521 => conv_std_logic_vector(36993, 16),
45522 => conv_std_logic_vector(37170, 16),
45523 => conv_std_logic_vector(37347, 16),
45524 => conv_std_logic_vector(37524, 16),
45525 => conv_std_logic_vector(37701, 16),
45526 => conv_std_logic_vector(37878, 16),
45527 => conv_std_logic_vector(38055, 16),
45528 => conv_std_logic_vector(38232, 16),
45529 => conv_std_logic_vector(38409, 16),
45530 => conv_std_logic_vector(38586, 16),
45531 => conv_std_logic_vector(38763, 16),
45532 => conv_std_logic_vector(38940, 16),
45533 => conv_std_logic_vector(39117, 16),
45534 => conv_std_logic_vector(39294, 16),
45535 => conv_std_logic_vector(39471, 16),
45536 => conv_std_logic_vector(39648, 16),
45537 => conv_std_logic_vector(39825, 16),
45538 => conv_std_logic_vector(40002, 16),
45539 => conv_std_logic_vector(40179, 16),
45540 => conv_std_logic_vector(40356, 16),
45541 => conv_std_logic_vector(40533, 16),
45542 => conv_std_logic_vector(40710, 16),
45543 => conv_std_logic_vector(40887, 16),
45544 => conv_std_logic_vector(41064, 16),
45545 => conv_std_logic_vector(41241, 16),
45546 => conv_std_logic_vector(41418, 16),
45547 => conv_std_logic_vector(41595, 16),
45548 => conv_std_logic_vector(41772, 16),
45549 => conv_std_logic_vector(41949, 16),
45550 => conv_std_logic_vector(42126, 16),
45551 => conv_std_logic_vector(42303, 16),
45552 => conv_std_logic_vector(42480, 16),
45553 => conv_std_logic_vector(42657, 16),
45554 => conv_std_logic_vector(42834, 16),
45555 => conv_std_logic_vector(43011, 16),
45556 => conv_std_logic_vector(43188, 16),
45557 => conv_std_logic_vector(43365, 16),
45558 => conv_std_logic_vector(43542, 16),
45559 => conv_std_logic_vector(43719, 16),
45560 => conv_std_logic_vector(43896, 16),
45561 => conv_std_logic_vector(44073, 16),
45562 => conv_std_logic_vector(44250, 16),
45563 => conv_std_logic_vector(44427, 16),
45564 => conv_std_logic_vector(44604, 16),
45565 => conv_std_logic_vector(44781, 16),
45566 => conv_std_logic_vector(44958, 16),
45567 => conv_std_logic_vector(45135, 16),
45568 => conv_std_logic_vector(0, 16),
45569 => conv_std_logic_vector(178, 16),
45570 => conv_std_logic_vector(356, 16),
45571 => conv_std_logic_vector(534, 16),
45572 => conv_std_logic_vector(712, 16),
45573 => conv_std_logic_vector(890, 16),
45574 => conv_std_logic_vector(1068, 16),
45575 => conv_std_logic_vector(1246, 16),
45576 => conv_std_logic_vector(1424, 16),
45577 => conv_std_logic_vector(1602, 16),
45578 => conv_std_logic_vector(1780, 16),
45579 => conv_std_logic_vector(1958, 16),
45580 => conv_std_logic_vector(2136, 16),
45581 => conv_std_logic_vector(2314, 16),
45582 => conv_std_logic_vector(2492, 16),
45583 => conv_std_logic_vector(2670, 16),
45584 => conv_std_logic_vector(2848, 16),
45585 => conv_std_logic_vector(3026, 16),
45586 => conv_std_logic_vector(3204, 16),
45587 => conv_std_logic_vector(3382, 16),
45588 => conv_std_logic_vector(3560, 16),
45589 => conv_std_logic_vector(3738, 16),
45590 => conv_std_logic_vector(3916, 16),
45591 => conv_std_logic_vector(4094, 16),
45592 => conv_std_logic_vector(4272, 16),
45593 => conv_std_logic_vector(4450, 16),
45594 => conv_std_logic_vector(4628, 16),
45595 => conv_std_logic_vector(4806, 16),
45596 => conv_std_logic_vector(4984, 16),
45597 => conv_std_logic_vector(5162, 16),
45598 => conv_std_logic_vector(5340, 16),
45599 => conv_std_logic_vector(5518, 16),
45600 => conv_std_logic_vector(5696, 16),
45601 => conv_std_logic_vector(5874, 16),
45602 => conv_std_logic_vector(6052, 16),
45603 => conv_std_logic_vector(6230, 16),
45604 => conv_std_logic_vector(6408, 16),
45605 => conv_std_logic_vector(6586, 16),
45606 => conv_std_logic_vector(6764, 16),
45607 => conv_std_logic_vector(6942, 16),
45608 => conv_std_logic_vector(7120, 16),
45609 => conv_std_logic_vector(7298, 16),
45610 => conv_std_logic_vector(7476, 16),
45611 => conv_std_logic_vector(7654, 16),
45612 => conv_std_logic_vector(7832, 16),
45613 => conv_std_logic_vector(8010, 16),
45614 => conv_std_logic_vector(8188, 16),
45615 => conv_std_logic_vector(8366, 16),
45616 => conv_std_logic_vector(8544, 16),
45617 => conv_std_logic_vector(8722, 16),
45618 => conv_std_logic_vector(8900, 16),
45619 => conv_std_logic_vector(9078, 16),
45620 => conv_std_logic_vector(9256, 16),
45621 => conv_std_logic_vector(9434, 16),
45622 => conv_std_logic_vector(9612, 16),
45623 => conv_std_logic_vector(9790, 16),
45624 => conv_std_logic_vector(9968, 16),
45625 => conv_std_logic_vector(10146, 16),
45626 => conv_std_logic_vector(10324, 16),
45627 => conv_std_logic_vector(10502, 16),
45628 => conv_std_logic_vector(10680, 16),
45629 => conv_std_logic_vector(10858, 16),
45630 => conv_std_logic_vector(11036, 16),
45631 => conv_std_logic_vector(11214, 16),
45632 => conv_std_logic_vector(11392, 16),
45633 => conv_std_logic_vector(11570, 16),
45634 => conv_std_logic_vector(11748, 16),
45635 => conv_std_logic_vector(11926, 16),
45636 => conv_std_logic_vector(12104, 16),
45637 => conv_std_logic_vector(12282, 16),
45638 => conv_std_logic_vector(12460, 16),
45639 => conv_std_logic_vector(12638, 16),
45640 => conv_std_logic_vector(12816, 16),
45641 => conv_std_logic_vector(12994, 16),
45642 => conv_std_logic_vector(13172, 16),
45643 => conv_std_logic_vector(13350, 16),
45644 => conv_std_logic_vector(13528, 16),
45645 => conv_std_logic_vector(13706, 16),
45646 => conv_std_logic_vector(13884, 16),
45647 => conv_std_logic_vector(14062, 16),
45648 => conv_std_logic_vector(14240, 16),
45649 => conv_std_logic_vector(14418, 16),
45650 => conv_std_logic_vector(14596, 16),
45651 => conv_std_logic_vector(14774, 16),
45652 => conv_std_logic_vector(14952, 16),
45653 => conv_std_logic_vector(15130, 16),
45654 => conv_std_logic_vector(15308, 16),
45655 => conv_std_logic_vector(15486, 16),
45656 => conv_std_logic_vector(15664, 16),
45657 => conv_std_logic_vector(15842, 16),
45658 => conv_std_logic_vector(16020, 16),
45659 => conv_std_logic_vector(16198, 16),
45660 => conv_std_logic_vector(16376, 16),
45661 => conv_std_logic_vector(16554, 16),
45662 => conv_std_logic_vector(16732, 16),
45663 => conv_std_logic_vector(16910, 16),
45664 => conv_std_logic_vector(17088, 16),
45665 => conv_std_logic_vector(17266, 16),
45666 => conv_std_logic_vector(17444, 16),
45667 => conv_std_logic_vector(17622, 16),
45668 => conv_std_logic_vector(17800, 16),
45669 => conv_std_logic_vector(17978, 16),
45670 => conv_std_logic_vector(18156, 16),
45671 => conv_std_logic_vector(18334, 16),
45672 => conv_std_logic_vector(18512, 16),
45673 => conv_std_logic_vector(18690, 16),
45674 => conv_std_logic_vector(18868, 16),
45675 => conv_std_logic_vector(19046, 16),
45676 => conv_std_logic_vector(19224, 16),
45677 => conv_std_logic_vector(19402, 16),
45678 => conv_std_logic_vector(19580, 16),
45679 => conv_std_logic_vector(19758, 16),
45680 => conv_std_logic_vector(19936, 16),
45681 => conv_std_logic_vector(20114, 16),
45682 => conv_std_logic_vector(20292, 16),
45683 => conv_std_logic_vector(20470, 16),
45684 => conv_std_logic_vector(20648, 16),
45685 => conv_std_logic_vector(20826, 16),
45686 => conv_std_logic_vector(21004, 16),
45687 => conv_std_logic_vector(21182, 16),
45688 => conv_std_logic_vector(21360, 16),
45689 => conv_std_logic_vector(21538, 16),
45690 => conv_std_logic_vector(21716, 16),
45691 => conv_std_logic_vector(21894, 16),
45692 => conv_std_logic_vector(22072, 16),
45693 => conv_std_logic_vector(22250, 16),
45694 => conv_std_logic_vector(22428, 16),
45695 => conv_std_logic_vector(22606, 16),
45696 => conv_std_logic_vector(22784, 16),
45697 => conv_std_logic_vector(22962, 16),
45698 => conv_std_logic_vector(23140, 16),
45699 => conv_std_logic_vector(23318, 16),
45700 => conv_std_logic_vector(23496, 16),
45701 => conv_std_logic_vector(23674, 16),
45702 => conv_std_logic_vector(23852, 16),
45703 => conv_std_logic_vector(24030, 16),
45704 => conv_std_logic_vector(24208, 16),
45705 => conv_std_logic_vector(24386, 16),
45706 => conv_std_logic_vector(24564, 16),
45707 => conv_std_logic_vector(24742, 16),
45708 => conv_std_logic_vector(24920, 16),
45709 => conv_std_logic_vector(25098, 16),
45710 => conv_std_logic_vector(25276, 16),
45711 => conv_std_logic_vector(25454, 16),
45712 => conv_std_logic_vector(25632, 16),
45713 => conv_std_logic_vector(25810, 16),
45714 => conv_std_logic_vector(25988, 16),
45715 => conv_std_logic_vector(26166, 16),
45716 => conv_std_logic_vector(26344, 16),
45717 => conv_std_logic_vector(26522, 16),
45718 => conv_std_logic_vector(26700, 16),
45719 => conv_std_logic_vector(26878, 16),
45720 => conv_std_logic_vector(27056, 16),
45721 => conv_std_logic_vector(27234, 16),
45722 => conv_std_logic_vector(27412, 16),
45723 => conv_std_logic_vector(27590, 16),
45724 => conv_std_logic_vector(27768, 16),
45725 => conv_std_logic_vector(27946, 16),
45726 => conv_std_logic_vector(28124, 16),
45727 => conv_std_logic_vector(28302, 16),
45728 => conv_std_logic_vector(28480, 16),
45729 => conv_std_logic_vector(28658, 16),
45730 => conv_std_logic_vector(28836, 16),
45731 => conv_std_logic_vector(29014, 16),
45732 => conv_std_logic_vector(29192, 16),
45733 => conv_std_logic_vector(29370, 16),
45734 => conv_std_logic_vector(29548, 16),
45735 => conv_std_logic_vector(29726, 16),
45736 => conv_std_logic_vector(29904, 16),
45737 => conv_std_logic_vector(30082, 16),
45738 => conv_std_logic_vector(30260, 16),
45739 => conv_std_logic_vector(30438, 16),
45740 => conv_std_logic_vector(30616, 16),
45741 => conv_std_logic_vector(30794, 16),
45742 => conv_std_logic_vector(30972, 16),
45743 => conv_std_logic_vector(31150, 16),
45744 => conv_std_logic_vector(31328, 16),
45745 => conv_std_logic_vector(31506, 16),
45746 => conv_std_logic_vector(31684, 16),
45747 => conv_std_logic_vector(31862, 16),
45748 => conv_std_logic_vector(32040, 16),
45749 => conv_std_logic_vector(32218, 16),
45750 => conv_std_logic_vector(32396, 16),
45751 => conv_std_logic_vector(32574, 16),
45752 => conv_std_logic_vector(32752, 16),
45753 => conv_std_logic_vector(32930, 16),
45754 => conv_std_logic_vector(33108, 16),
45755 => conv_std_logic_vector(33286, 16),
45756 => conv_std_logic_vector(33464, 16),
45757 => conv_std_logic_vector(33642, 16),
45758 => conv_std_logic_vector(33820, 16),
45759 => conv_std_logic_vector(33998, 16),
45760 => conv_std_logic_vector(34176, 16),
45761 => conv_std_logic_vector(34354, 16),
45762 => conv_std_logic_vector(34532, 16),
45763 => conv_std_logic_vector(34710, 16),
45764 => conv_std_logic_vector(34888, 16),
45765 => conv_std_logic_vector(35066, 16),
45766 => conv_std_logic_vector(35244, 16),
45767 => conv_std_logic_vector(35422, 16),
45768 => conv_std_logic_vector(35600, 16),
45769 => conv_std_logic_vector(35778, 16),
45770 => conv_std_logic_vector(35956, 16),
45771 => conv_std_logic_vector(36134, 16),
45772 => conv_std_logic_vector(36312, 16),
45773 => conv_std_logic_vector(36490, 16),
45774 => conv_std_logic_vector(36668, 16),
45775 => conv_std_logic_vector(36846, 16),
45776 => conv_std_logic_vector(37024, 16),
45777 => conv_std_logic_vector(37202, 16),
45778 => conv_std_logic_vector(37380, 16),
45779 => conv_std_logic_vector(37558, 16),
45780 => conv_std_logic_vector(37736, 16),
45781 => conv_std_logic_vector(37914, 16),
45782 => conv_std_logic_vector(38092, 16),
45783 => conv_std_logic_vector(38270, 16),
45784 => conv_std_logic_vector(38448, 16),
45785 => conv_std_logic_vector(38626, 16),
45786 => conv_std_logic_vector(38804, 16),
45787 => conv_std_logic_vector(38982, 16),
45788 => conv_std_logic_vector(39160, 16),
45789 => conv_std_logic_vector(39338, 16),
45790 => conv_std_logic_vector(39516, 16),
45791 => conv_std_logic_vector(39694, 16),
45792 => conv_std_logic_vector(39872, 16),
45793 => conv_std_logic_vector(40050, 16),
45794 => conv_std_logic_vector(40228, 16),
45795 => conv_std_logic_vector(40406, 16),
45796 => conv_std_logic_vector(40584, 16),
45797 => conv_std_logic_vector(40762, 16),
45798 => conv_std_logic_vector(40940, 16),
45799 => conv_std_logic_vector(41118, 16),
45800 => conv_std_logic_vector(41296, 16),
45801 => conv_std_logic_vector(41474, 16),
45802 => conv_std_logic_vector(41652, 16),
45803 => conv_std_logic_vector(41830, 16),
45804 => conv_std_logic_vector(42008, 16),
45805 => conv_std_logic_vector(42186, 16),
45806 => conv_std_logic_vector(42364, 16),
45807 => conv_std_logic_vector(42542, 16),
45808 => conv_std_logic_vector(42720, 16),
45809 => conv_std_logic_vector(42898, 16),
45810 => conv_std_logic_vector(43076, 16),
45811 => conv_std_logic_vector(43254, 16),
45812 => conv_std_logic_vector(43432, 16),
45813 => conv_std_logic_vector(43610, 16),
45814 => conv_std_logic_vector(43788, 16),
45815 => conv_std_logic_vector(43966, 16),
45816 => conv_std_logic_vector(44144, 16),
45817 => conv_std_logic_vector(44322, 16),
45818 => conv_std_logic_vector(44500, 16),
45819 => conv_std_logic_vector(44678, 16),
45820 => conv_std_logic_vector(44856, 16),
45821 => conv_std_logic_vector(45034, 16),
45822 => conv_std_logic_vector(45212, 16),
45823 => conv_std_logic_vector(45390, 16),
45824 => conv_std_logic_vector(0, 16),
45825 => conv_std_logic_vector(179, 16),
45826 => conv_std_logic_vector(358, 16),
45827 => conv_std_logic_vector(537, 16),
45828 => conv_std_logic_vector(716, 16),
45829 => conv_std_logic_vector(895, 16),
45830 => conv_std_logic_vector(1074, 16),
45831 => conv_std_logic_vector(1253, 16),
45832 => conv_std_logic_vector(1432, 16),
45833 => conv_std_logic_vector(1611, 16),
45834 => conv_std_logic_vector(1790, 16),
45835 => conv_std_logic_vector(1969, 16),
45836 => conv_std_logic_vector(2148, 16),
45837 => conv_std_logic_vector(2327, 16),
45838 => conv_std_logic_vector(2506, 16),
45839 => conv_std_logic_vector(2685, 16),
45840 => conv_std_logic_vector(2864, 16),
45841 => conv_std_logic_vector(3043, 16),
45842 => conv_std_logic_vector(3222, 16),
45843 => conv_std_logic_vector(3401, 16),
45844 => conv_std_logic_vector(3580, 16),
45845 => conv_std_logic_vector(3759, 16),
45846 => conv_std_logic_vector(3938, 16),
45847 => conv_std_logic_vector(4117, 16),
45848 => conv_std_logic_vector(4296, 16),
45849 => conv_std_logic_vector(4475, 16),
45850 => conv_std_logic_vector(4654, 16),
45851 => conv_std_logic_vector(4833, 16),
45852 => conv_std_logic_vector(5012, 16),
45853 => conv_std_logic_vector(5191, 16),
45854 => conv_std_logic_vector(5370, 16),
45855 => conv_std_logic_vector(5549, 16),
45856 => conv_std_logic_vector(5728, 16),
45857 => conv_std_logic_vector(5907, 16),
45858 => conv_std_logic_vector(6086, 16),
45859 => conv_std_logic_vector(6265, 16),
45860 => conv_std_logic_vector(6444, 16),
45861 => conv_std_logic_vector(6623, 16),
45862 => conv_std_logic_vector(6802, 16),
45863 => conv_std_logic_vector(6981, 16),
45864 => conv_std_logic_vector(7160, 16),
45865 => conv_std_logic_vector(7339, 16),
45866 => conv_std_logic_vector(7518, 16),
45867 => conv_std_logic_vector(7697, 16),
45868 => conv_std_logic_vector(7876, 16),
45869 => conv_std_logic_vector(8055, 16),
45870 => conv_std_logic_vector(8234, 16),
45871 => conv_std_logic_vector(8413, 16),
45872 => conv_std_logic_vector(8592, 16),
45873 => conv_std_logic_vector(8771, 16),
45874 => conv_std_logic_vector(8950, 16),
45875 => conv_std_logic_vector(9129, 16),
45876 => conv_std_logic_vector(9308, 16),
45877 => conv_std_logic_vector(9487, 16),
45878 => conv_std_logic_vector(9666, 16),
45879 => conv_std_logic_vector(9845, 16),
45880 => conv_std_logic_vector(10024, 16),
45881 => conv_std_logic_vector(10203, 16),
45882 => conv_std_logic_vector(10382, 16),
45883 => conv_std_logic_vector(10561, 16),
45884 => conv_std_logic_vector(10740, 16),
45885 => conv_std_logic_vector(10919, 16),
45886 => conv_std_logic_vector(11098, 16),
45887 => conv_std_logic_vector(11277, 16),
45888 => conv_std_logic_vector(11456, 16),
45889 => conv_std_logic_vector(11635, 16),
45890 => conv_std_logic_vector(11814, 16),
45891 => conv_std_logic_vector(11993, 16),
45892 => conv_std_logic_vector(12172, 16),
45893 => conv_std_logic_vector(12351, 16),
45894 => conv_std_logic_vector(12530, 16),
45895 => conv_std_logic_vector(12709, 16),
45896 => conv_std_logic_vector(12888, 16),
45897 => conv_std_logic_vector(13067, 16),
45898 => conv_std_logic_vector(13246, 16),
45899 => conv_std_logic_vector(13425, 16),
45900 => conv_std_logic_vector(13604, 16),
45901 => conv_std_logic_vector(13783, 16),
45902 => conv_std_logic_vector(13962, 16),
45903 => conv_std_logic_vector(14141, 16),
45904 => conv_std_logic_vector(14320, 16),
45905 => conv_std_logic_vector(14499, 16),
45906 => conv_std_logic_vector(14678, 16),
45907 => conv_std_logic_vector(14857, 16),
45908 => conv_std_logic_vector(15036, 16),
45909 => conv_std_logic_vector(15215, 16),
45910 => conv_std_logic_vector(15394, 16),
45911 => conv_std_logic_vector(15573, 16),
45912 => conv_std_logic_vector(15752, 16),
45913 => conv_std_logic_vector(15931, 16),
45914 => conv_std_logic_vector(16110, 16),
45915 => conv_std_logic_vector(16289, 16),
45916 => conv_std_logic_vector(16468, 16),
45917 => conv_std_logic_vector(16647, 16),
45918 => conv_std_logic_vector(16826, 16),
45919 => conv_std_logic_vector(17005, 16),
45920 => conv_std_logic_vector(17184, 16),
45921 => conv_std_logic_vector(17363, 16),
45922 => conv_std_logic_vector(17542, 16),
45923 => conv_std_logic_vector(17721, 16),
45924 => conv_std_logic_vector(17900, 16),
45925 => conv_std_logic_vector(18079, 16),
45926 => conv_std_logic_vector(18258, 16),
45927 => conv_std_logic_vector(18437, 16),
45928 => conv_std_logic_vector(18616, 16),
45929 => conv_std_logic_vector(18795, 16),
45930 => conv_std_logic_vector(18974, 16),
45931 => conv_std_logic_vector(19153, 16),
45932 => conv_std_logic_vector(19332, 16),
45933 => conv_std_logic_vector(19511, 16),
45934 => conv_std_logic_vector(19690, 16),
45935 => conv_std_logic_vector(19869, 16),
45936 => conv_std_logic_vector(20048, 16),
45937 => conv_std_logic_vector(20227, 16),
45938 => conv_std_logic_vector(20406, 16),
45939 => conv_std_logic_vector(20585, 16),
45940 => conv_std_logic_vector(20764, 16),
45941 => conv_std_logic_vector(20943, 16),
45942 => conv_std_logic_vector(21122, 16),
45943 => conv_std_logic_vector(21301, 16),
45944 => conv_std_logic_vector(21480, 16),
45945 => conv_std_logic_vector(21659, 16),
45946 => conv_std_logic_vector(21838, 16),
45947 => conv_std_logic_vector(22017, 16),
45948 => conv_std_logic_vector(22196, 16),
45949 => conv_std_logic_vector(22375, 16),
45950 => conv_std_logic_vector(22554, 16),
45951 => conv_std_logic_vector(22733, 16),
45952 => conv_std_logic_vector(22912, 16),
45953 => conv_std_logic_vector(23091, 16),
45954 => conv_std_logic_vector(23270, 16),
45955 => conv_std_logic_vector(23449, 16),
45956 => conv_std_logic_vector(23628, 16),
45957 => conv_std_logic_vector(23807, 16),
45958 => conv_std_logic_vector(23986, 16),
45959 => conv_std_logic_vector(24165, 16),
45960 => conv_std_logic_vector(24344, 16),
45961 => conv_std_logic_vector(24523, 16),
45962 => conv_std_logic_vector(24702, 16),
45963 => conv_std_logic_vector(24881, 16),
45964 => conv_std_logic_vector(25060, 16),
45965 => conv_std_logic_vector(25239, 16),
45966 => conv_std_logic_vector(25418, 16),
45967 => conv_std_logic_vector(25597, 16),
45968 => conv_std_logic_vector(25776, 16),
45969 => conv_std_logic_vector(25955, 16),
45970 => conv_std_logic_vector(26134, 16),
45971 => conv_std_logic_vector(26313, 16),
45972 => conv_std_logic_vector(26492, 16),
45973 => conv_std_logic_vector(26671, 16),
45974 => conv_std_logic_vector(26850, 16),
45975 => conv_std_logic_vector(27029, 16),
45976 => conv_std_logic_vector(27208, 16),
45977 => conv_std_logic_vector(27387, 16),
45978 => conv_std_logic_vector(27566, 16),
45979 => conv_std_logic_vector(27745, 16),
45980 => conv_std_logic_vector(27924, 16),
45981 => conv_std_logic_vector(28103, 16),
45982 => conv_std_logic_vector(28282, 16),
45983 => conv_std_logic_vector(28461, 16),
45984 => conv_std_logic_vector(28640, 16),
45985 => conv_std_logic_vector(28819, 16),
45986 => conv_std_logic_vector(28998, 16),
45987 => conv_std_logic_vector(29177, 16),
45988 => conv_std_logic_vector(29356, 16),
45989 => conv_std_logic_vector(29535, 16),
45990 => conv_std_logic_vector(29714, 16),
45991 => conv_std_logic_vector(29893, 16),
45992 => conv_std_logic_vector(30072, 16),
45993 => conv_std_logic_vector(30251, 16),
45994 => conv_std_logic_vector(30430, 16),
45995 => conv_std_logic_vector(30609, 16),
45996 => conv_std_logic_vector(30788, 16),
45997 => conv_std_logic_vector(30967, 16),
45998 => conv_std_logic_vector(31146, 16),
45999 => conv_std_logic_vector(31325, 16),
46000 => conv_std_logic_vector(31504, 16),
46001 => conv_std_logic_vector(31683, 16),
46002 => conv_std_logic_vector(31862, 16),
46003 => conv_std_logic_vector(32041, 16),
46004 => conv_std_logic_vector(32220, 16),
46005 => conv_std_logic_vector(32399, 16),
46006 => conv_std_logic_vector(32578, 16),
46007 => conv_std_logic_vector(32757, 16),
46008 => conv_std_logic_vector(32936, 16),
46009 => conv_std_logic_vector(33115, 16),
46010 => conv_std_logic_vector(33294, 16),
46011 => conv_std_logic_vector(33473, 16),
46012 => conv_std_logic_vector(33652, 16),
46013 => conv_std_logic_vector(33831, 16),
46014 => conv_std_logic_vector(34010, 16),
46015 => conv_std_logic_vector(34189, 16),
46016 => conv_std_logic_vector(34368, 16),
46017 => conv_std_logic_vector(34547, 16),
46018 => conv_std_logic_vector(34726, 16),
46019 => conv_std_logic_vector(34905, 16),
46020 => conv_std_logic_vector(35084, 16),
46021 => conv_std_logic_vector(35263, 16),
46022 => conv_std_logic_vector(35442, 16),
46023 => conv_std_logic_vector(35621, 16),
46024 => conv_std_logic_vector(35800, 16),
46025 => conv_std_logic_vector(35979, 16),
46026 => conv_std_logic_vector(36158, 16),
46027 => conv_std_logic_vector(36337, 16),
46028 => conv_std_logic_vector(36516, 16),
46029 => conv_std_logic_vector(36695, 16),
46030 => conv_std_logic_vector(36874, 16),
46031 => conv_std_logic_vector(37053, 16),
46032 => conv_std_logic_vector(37232, 16),
46033 => conv_std_logic_vector(37411, 16),
46034 => conv_std_logic_vector(37590, 16),
46035 => conv_std_logic_vector(37769, 16),
46036 => conv_std_logic_vector(37948, 16),
46037 => conv_std_logic_vector(38127, 16),
46038 => conv_std_logic_vector(38306, 16),
46039 => conv_std_logic_vector(38485, 16),
46040 => conv_std_logic_vector(38664, 16),
46041 => conv_std_logic_vector(38843, 16),
46042 => conv_std_logic_vector(39022, 16),
46043 => conv_std_logic_vector(39201, 16),
46044 => conv_std_logic_vector(39380, 16),
46045 => conv_std_logic_vector(39559, 16),
46046 => conv_std_logic_vector(39738, 16),
46047 => conv_std_logic_vector(39917, 16),
46048 => conv_std_logic_vector(40096, 16),
46049 => conv_std_logic_vector(40275, 16),
46050 => conv_std_logic_vector(40454, 16),
46051 => conv_std_logic_vector(40633, 16),
46052 => conv_std_logic_vector(40812, 16),
46053 => conv_std_logic_vector(40991, 16),
46054 => conv_std_logic_vector(41170, 16),
46055 => conv_std_logic_vector(41349, 16),
46056 => conv_std_logic_vector(41528, 16),
46057 => conv_std_logic_vector(41707, 16),
46058 => conv_std_logic_vector(41886, 16),
46059 => conv_std_logic_vector(42065, 16),
46060 => conv_std_logic_vector(42244, 16),
46061 => conv_std_logic_vector(42423, 16),
46062 => conv_std_logic_vector(42602, 16),
46063 => conv_std_logic_vector(42781, 16),
46064 => conv_std_logic_vector(42960, 16),
46065 => conv_std_logic_vector(43139, 16),
46066 => conv_std_logic_vector(43318, 16),
46067 => conv_std_logic_vector(43497, 16),
46068 => conv_std_logic_vector(43676, 16),
46069 => conv_std_logic_vector(43855, 16),
46070 => conv_std_logic_vector(44034, 16),
46071 => conv_std_logic_vector(44213, 16),
46072 => conv_std_logic_vector(44392, 16),
46073 => conv_std_logic_vector(44571, 16),
46074 => conv_std_logic_vector(44750, 16),
46075 => conv_std_logic_vector(44929, 16),
46076 => conv_std_logic_vector(45108, 16),
46077 => conv_std_logic_vector(45287, 16),
46078 => conv_std_logic_vector(45466, 16),
46079 => conv_std_logic_vector(45645, 16),
46080 => conv_std_logic_vector(0, 16),
46081 => conv_std_logic_vector(180, 16),
46082 => conv_std_logic_vector(360, 16),
46083 => conv_std_logic_vector(540, 16),
46084 => conv_std_logic_vector(720, 16),
46085 => conv_std_logic_vector(900, 16),
46086 => conv_std_logic_vector(1080, 16),
46087 => conv_std_logic_vector(1260, 16),
46088 => conv_std_logic_vector(1440, 16),
46089 => conv_std_logic_vector(1620, 16),
46090 => conv_std_logic_vector(1800, 16),
46091 => conv_std_logic_vector(1980, 16),
46092 => conv_std_logic_vector(2160, 16),
46093 => conv_std_logic_vector(2340, 16),
46094 => conv_std_logic_vector(2520, 16),
46095 => conv_std_logic_vector(2700, 16),
46096 => conv_std_logic_vector(2880, 16),
46097 => conv_std_logic_vector(3060, 16),
46098 => conv_std_logic_vector(3240, 16),
46099 => conv_std_logic_vector(3420, 16),
46100 => conv_std_logic_vector(3600, 16),
46101 => conv_std_logic_vector(3780, 16),
46102 => conv_std_logic_vector(3960, 16),
46103 => conv_std_logic_vector(4140, 16),
46104 => conv_std_logic_vector(4320, 16),
46105 => conv_std_logic_vector(4500, 16),
46106 => conv_std_logic_vector(4680, 16),
46107 => conv_std_logic_vector(4860, 16),
46108 => conv_std_logic_vector(5040, 16),
46109 => conv_std_logic_vector(5220, 16),
46110 => conv_std_logic_vector(5400, 16),
46111 => conv_std_logic_vector(5580, 16),
46112 => conv_std_logic_vector(5760, 16),
46113 => conv_std_logic_vector(5940, 16),
46114 => conv_std_logic_vector(6120, 16),
46115 => conv_std_logic_vector(6300, 16),
46116 => conv_std_logic_vector(6480, 16),
46117 => conv_std_logic_vector(6660, 16),
46118 => conv_std_logic_vector(6840, 16),
46119 => conv_std_logic_vector(7020, 16),
46120 => conv_std_logic_vector(7200, 16),
46121 => conv_std_logic_vector(7380, 16),
46122 => conv_std_logic_vector(7560, 16),
46123 => conv_std_logic_vector(7740, 16),
46124 => conv_std_logic_vector(7920, 16),
46125 => conv_std_logic_vector(8100, 16),
46126 => conv_std_logic_vector(8280, 16),
46127 => conv_std_logic_vector(8460, 16),
46128 => conv_std_logic_vector(8640, 16),
46129 => conv_std_logic_vector(8820, 16),
46130 => conv_std_logic_vector(9000, 16),
46131 => conv_std_logic_vector(9180, 16),
46132 => conv_std_logic_vector(9360, 16),
46133 => conv_std_logic_vector(9540, 16),
46134 => conv_std_logic_vector(9720, 16),
46135 => conv_std_logic_vector(9900, 16),
46136 => conv_std_logic_vector(10080, 16),
46137 => conv_std_logic_vector(10260, 16),
46138 => conv_std_logic_vector(10440, 16),
46139 => conv_std_logic_vector(10620, 16),
46140 => conv_std_logic_vector(10800, 16),
46141 => conv_std_logic_vector(10980, 16),
46142 => conv_std_logic_vector(11160, 16),
46143 => conv_std_logic_vector(11340, 16),
46144 => conv_std_logic_vector(11520, 16),
46145 => conv_std_logic_vector(11700, 16),
46146 => conv_std_logic_vector(11880, 16),
46147 => conv_std_logic_vector(12060, 16),
46148 => conv_std_logic_vector(12240, 16),
46149 => conv_std_logic_vector(12420, 16),
46150 => conv_std_logic_vector(12600, 16),
46151 => conv_std_logic_vector(12780, 16),
46152 => conv_std_logic_vector(12960, 16),
46153 => conv_std_logic_vector(13140, 16),
46154 => conv_std_logic_vector(13320, 16),
46155 => conv_std_logic_vector(13500, 16),
46156 => conv_std_logic_vector(13680, 16),
46157 => conv_std_logic_vector(13860, 16),
46158 => conv_std_logic_vector(14040, 16),
46159 => conv_std_logic_vector(14220, 16),
46160 => conv_std_logic_vector(14400, 16),
46161 => conv_std_logic_vector(14580, 16),
46162 => conv_std_logic_vector(14760, 16),
46163 => conv_std_logic_vector(14940, 16),
46164 => conv_std_logic_vector(15120, 16),
46165 => conv_std_logic_vector(15300, 16),
46166 => conv_std_logic_vector(15480, 16),
46167 => conv_std_logic_vector(15660, 16),
46168 => conv_std_logic_vector(15840, 16),
46169 => conv_std_logic_vector(16020, 16),
46170 => conv_std_logic_vector(16200, 16),
46171 => conv_std_logic_vector(16380, 16),
46172 => conv_std_logic_vector(16560, 16),
46173 => conv_std_logic_vector(16740, 16),
46174 => conv_std_logic_vector(16920, 16),
46175 => conv_std_logic_vector(17100, 16),
46176 => conv_std_logic_vector(17280, 16),
46177 => conv_std_logic_vector(17460, 16),
46178 => conv_std_logic_vector(17640, 16),
46179 => conv_std_logic_vector(17820, 16),
46180 => conv_std_logic_vector(18000, 16),
46181 => conv_std_logic_vector(18180, 16),
46182 => conv_std_logic_vector(18360, 16),
46183 => conv_std_logic_vector(18540, 16),
46184 => conv_std_logic_vector(18720, 16),
46185 => conv_std_logic_vector(18900, 16),
46186 => conv_std_logic_vector(19080, 16),
46187 => conv_std_logic_vector(19260, 16),
46188 => conv_std_logic_vector(19440, 16),
46189 => conv_std_logic_vector(19620, 16),
46190 => conv_std_logic_vector(19800, 16),
46191 => conv_std_logic_vector(19980, 16),
46192 => conv_std_logic_vector(20160, 16),
46193 => conv_std_logic_vector(20340, 16),
46194 => conv_std_logic_vector(20520, 16),
46195 => conv_std_logic_vector(20700, 16),
46196 => conv_std_logic_vector(20880, 16),
46197 => conv_std_logic_vector(21060, 16),
46198 => conv_std_logic_vector(21240, 16),
46199 => conv_std_logic_vector(21420, 16),
46200 => conv_std_logic_vector(21600, 16),
46201 => conv_std_logic_vector(21780, 16),
46202 => conv_std_logic_vector(21960, 16),
46203 => conv_std_logic_vector(22140, 16),
46204 => conv_std_logic_vector(22320, 16),
46205 => conv_std_logic_vector(22500, 16),
46206 => conv_std_logic_vector(22680, 16),
46207 => conv_std_logic_vector(22860, 16),
46208 => conv_std_logic_vector(23040, 16),
46209 => conv_std_logic_vector(23220, 16),
46210 => conv_std_logic_vector(23400, 16),
46211 => conv_std_logic_vector(23580, 16),
46212 => conv_std_logic_vector(23760, 16),
46213 => conv_std_logic_vector(23940, 16),
46214 => conv_std_logic_vector(24120, 16),
46215 => conv_std_logic_vector(24300, 16),
46216 => conv_std_logic_vector(24480, 16),
46217 => conv_std_logic_vector(24660, 16),
46218 => conv_std_logic_vector(24840, 16),
46219 => conv_std_logic_vector(25020, 16),
46220 => conv_std_logic_vector(25200, 16),
46221 => conv_std_logic_vector(25380, 16),
46222 => conv_std_logic_vector(25560, 16),
46223 => conv_std_logic_vector(25740, 16),
46224 => conv_std_logic_vector(25920, 16),
46225 => conv_std_logic_vector(26100, 16),
46226 => conv_std_logic_vector(26280, 16),
46227 => conv_std_logic_vector(26460, 16),
46228 => conv_std_logic_vector(26640, 16),
46229 => conv_std_logic_vector(26820, 16),
46230 => conv_std_logic_vector(27000, 16),
46231 => conv_std_logic_vector(27180, 16),
46232 => conv_std_logic_vector(27360, 16),
46233 => conv_std_logic_vector(27540, 16),
46234 => conv_std_logic_vector(27720, 16),
46235 => conv_std_logic_vector(27900, 16),
46236 => conv_std_logic_vector(28080, 16),
46237 => conv_std_logic_vector(28260, 16),
46238 => conv_std_logic_vector(28440, 16),
46239 => conv_std_logic_vector(28620, 16),
46240 => conv_std_logic_vector(28800, 16),
46241 => conv_std_logic_vector(28980, 16),
46242 => conv_std_logic_vector(29160, 16),
46243 => conv_std_logic_vector(29340, 16),
46244 => conv_std_logic_vector(29520, 16),
46245 => conv_std_logic_vector(29700, 16),
46246 => conv_std_logic_vector(29880, 16),
46247 => conv_std_logic_vector(30060, 16),
46248 => conv_std_logic_vector(30240, 16),
46249 => conv_std_logic_vector(30420, 16),
46250 => conv_std_logic_vector(30600, 16),
46251 => conv_std_logic_vector(30780, 16),
46252 => conv_std_logic_vector(30960, 16),
46253 => conv_std_logic_vector(31140, 16),
46254 => conv_std_logic_vector(31320, 16),
46255 => conv_std_logic_vector(31500, 16),
46256 => conv_std_logic_vector(31680, 16),
46257 => conv_std_logic_vector(31860, 16),
46258 => conv_std_logic_vector(32040, 16),
46259 => conv_std_logic_vector(32220, 16),
46260 => conv_std_logic_vector(32400, 16),
46261 => conv_std_logic_vector(32580, 16),
46262 => conv_std_logic_vector(32760, 16),
46263 => conv_std_logic_vector(32940, 16),
46264 => conv_std_logic_vector(33120, 16),
46265 => conv_std_logic_vector(33300, 16),
46266 => conv_std_logic_vector(33480, 16),
46267 => conv_std_logic_vector(33660, 16),
46268 => conv_std_logic_vector(33840, 16),
46269 => conv_std_logic_vector(34020, 16),
46270 => conv_std_logic_vector(34200, 16),
46271 => conv_std_logic_vector(34380, 16),
46272 => conv_std_logic_vector(34560, 16),
46273 => conv_std_logic_vector(34740, 16),
46274 => conv_std_logic_vector(34920, 16),
46275 => conv_std_logic_vector(35100, 16),
46276 => conv_std_logic_vector(35280, 16),
46277 => conv_std_logic_vector(35460, 16),
46278 => conv_std_logic_vector(35640, 16),
46279 => conv_std_logic_vector(35820, 16),
46280 => conv_std_logic_vector(36000, 16),
46281 => conv_std_logic_vector(36180, 16),
46282 => conv_std_logic_vector(36360, 16),
46283 => conv_std_logic_vector(36540, 16),
46284 => conv_std_logic_vector(36720, 16),
46285 => conv_std_logic_vector(36900, 16),
46286 => conv_std_logic_vector(37080, 16),
46287 => conv_std_logic_vector(37260, 16),
46288 => conv_std_logic_vector(37440, 16),
46289 => conv_std_logic_vector(37620, 16),
46290 => conv_std_logic_vector(37800, 16),
46291 => conv_std_logic_vector(37980, 16),
46292 => conv_std_logic_vector(38160, 16),
46293 => conv_std_logic_vector(38340, 16),
46294 => conv_std_logic_vector(38520, 16),
46295 => conv_std_logic_vector(38700, 16),
46296 => conv_std_logic_vector(38880, 16),
46297 => conv_std_logic_vector(39060, 16),
46298 => conv_std_logic_vector(39240, 16),
46299 => conv_std_logic_vector(39420, 16),
46300 => conv_std_logic_vector(39600, 16),
46301 => conv_std_logic_vector(39780, 16),
46302 => conv_std_logic_vector(39960, 16),
46303 => conv_std_logic_vector(40140, 16),
46304 => conv_std_logic_vector(40320, 16),
46305 => conv_std_logic_vector(40500, 16),
46306 => conv_std_logic_vector(40680, 16),
46307 => conv_std_logic_vector(40860, 16),
46308 => conv_std_logic_vector(41040, 16),
46309 => conv_std_logic_vector(41220, 16),
46310 => conv_std_logic_vector(41400, 16),
46311 => conv_std_logic_vector(41580, 16),
46312 => conv_std_logic_vector(41760, 16),
46313 => conv_std_logic_vector(41940, 16),
46314 => conv_std_logic_vector(42120, 16),
46315 => conv_std_logic_vector(42300, 16),
46316 => conv_std_logic_vector(42480, 16),
46317 => conv_std_logic_vector(42660, 16),
46318 => conv_std_logic_vector(42840, 16),
46319 => conv_std_logic_vector(43020, 16),
46320 => conv_std_logic_vector(43200, 16),
46321 => conv_std_logic_vector(43380, 16),
46322 => conv_std_logic_vector(43560, 16),
46323 => conv_std_logic_vector(43740, 16),
46324 => conv_std_logic_vector(43920, 16),
46325 => conv_std_logic_vector(44100, 16),
46326 => conv_std_logic_vector(44280, 16),
46327 => conv_std_logic_vector(44460, 16),
46328 => conv_std_logic_vector(44640, 16),
46329 => conv_std_logic_vector(44820, 16),
46330 => conv_std_logic_vector(45000, 16),
46331 => conv_std_logic_vector(45180, 16),
46332 => conv_std_logic_vector(45360, 16),
46333 => conv_std_logic_vector(45540, 16),
46334 => conv_std_logic_vector(45720, 16),
46335 => conv_std_logic_vector(45900, 16),
46336 => conv_std_logic_vector(0, 16),
46337 => conv_std_logic_vector(181, 16),
46338 => conv_std_logic_vector(362, 16),
46339 => conv_std_logic_vector(543, 16),
46340 => conv_std_logic_vector(724, 16),
46341 => conv_std_logic_vector(905, 16),
46342 => conv_std_logic_vector(1086, 16),
46343 => conv_std_logic_vector(1267, 16),
46344 => conv_std_logic_vector(1448, 16),
46345 => conv_std_logic_vector(1629, 16),
46346 => conv_std_logic_vector(1810, 16),
46347 => conv_std_logic_vector(1991, 16),
46348 => conv_std_logic_vector(2172, 16),
46349 => conv_std_logic_vector(2353, 16),
46350 => conv_std_logic_vector(2534, 16),
46351 => conv_std_logic_vector(2715, 16),
46352 => conv_std_logic_vector(2896, 16),
46353 => conv_std_logic_vector(3077, 16),
46354 => conv_std_logic_vector(3258, 16),
46355 => conv_std_logic_vector(3439, 16),
46356 => conv_std_logic_vector(3620, 16),
46357 => conv_std_logic_vector(3801, 16),
46358 => conv_std_logic_vector(3982, 16),
46359 => conv_std_logic_vector(4163, 16),
46360 => conv_std_logic_vector(4344, 16),
46361 => conv_std_logic_vector(4525, 16),
46362 => conv_std_logic_vector(4706, 16),
46363 => conv_std_logic_vector(4887, 16),
46364 => conv_std_logic_vector(5068, 16),
46365 => conv_std_logic_vector(5249, 16),
46366 => conv_std_logic_vector(5430, 16),
46367 => conv_std_logic_vector(5611, 16),
46368 => conv_std_logic_vector(5792, 16),
46369 => conv_std_logic_vector(5973, 16),
46370 => conv_std_logic_vector(6154, 16),
46371 => conv_std_logic_vector(6335, 16),
46372 => conv_std_logic_vector(6516, 16),
46373 => conv_std_logic_vector(6697, 16),
46374 => conv_std_logic_vector(6878, 16),
46375 => conv_std_logic_vector(7059, 16),
46376 => conv_std_logic_vector(7240, 16),
46377 => conv_std_logic_vector(7421, 16),
46378 => conv_std_logic_vector(7602, 16),
46379 => conv_std_logic_vector(7783, 16),
46380 => conv_std_logic_vector(7964, 16),
46381 => conv_std_logic_vector(8145, 16),
46382 => conv_std_logic_vector(8326, 16),
46383 => conv_std_logic_vector(8507, 16),
46384 => conv_std_logic_vector(8688, 16),
46385 => conv_std_logic_vector(8869, 16),
46386 => conv_std_logic_vector(9050, 16),
46387 => conv_std_logic_vector(9231, 16),
46388 => conv_std_logic_vector(9412, 16),
46389 => conv_std_logic_vector(9593, 16),
46390 => conv_std_logic_vector(9774, 16),
46391 => conv_std_logic_vector(9955, 16),
46392 => conv_std_logic_vector(10136, 16),
46393 => conv_std_logic_vector(10317, 16),
46394 => conv_std_logic_vector(10498, 16),
46395 => conv_std_logic_vector(10679, 16),
46396 => conv_std_logic_vector(10860, 16),
46397 => conv_std_logic_vector(11041, 16),
46398 => conv_std_logic_vector(11222, 16),
46399 => conv_std_logic_vector(11403, 16),
46400 => conv_std_logic_vector(11584, 16),
46401 => conv_std_logic_vector(11765, 16),
46402 => conv_std_logic_vector(11946, 16),
46403 => conv_std_logic_vector(12127, 16),
46404 => conv_std_logic_vector(12308, 16),
46405 => conv_std_logic_vector(12489, 16),
46406 => conv_std_logic_vector(12670, 16),
46407 => conv_std_logic_vector(12851, 16),
46408 => conv_std_logic_vector(13032, 16),
46409 => conv_std_logic_vector(13213, 16),
46410 => conv_std_logic_vector(13394, 16),
46411 => conv_std_logic_vector(13575, 16),
46412 => conv_std_logic_vector(13756, 16),
46413 => conv_std_logic_vector(13937, 16),
46414 => conv_std_logic_vector(14118, 16),
46415 => conv_std_logic_vector(14299, 16),
46416 => conv_std_logic_vector(14480, 16),
46417 => conv_std_logic_vector(14661, 16),
46418 => conv_std_logic_vector(14842, 16),
46419 => conv_std_logic_vector(15023, 16),
46420 => conv_std_logic_vector(15204, 16),
46421 => conv_std_logic_vector(15385, 16),
46422 => conv_std_logic_vector(15566, 16),
46423 => conv_std_logic_vector(15747, 16),
46424 => conv_std_logic_vector(15928, 16),
46425 => conv_std_logic_vector(16109, 16),
46426 => conv_std_logic_vector(16290, 16),
46427 => conv_std_logic_vector(16471, 16),
46428 => conv_std_logic_vector(16652, 16),
46429 => conv_std_logic_vector(16833, 16),
46430 => conv_std_logic_vector(17014, 16),
46431 => conv_std_logic_vector(17195, 16),
46432 => conv_std_logic_vector(17376, 16),
46433 => conv_std_logic_vector(17557, 16),
46434 => conv_std_logic_vector(17738, 16),
46435 => conv_std_logic_vector(17919, 16),
46436 => conv_std_logic_vector(18100, 16),
46437 => conv_std_logic_vector(18281, 16),
46438 => conv_std_logic_vector(18462, 16),
46439 => conv_std_logic_vector(18643, 16),
46440 => conv_std_logic_vector(18824, 16),
46441 => conv_std_logic_vector(19005, 16),
46442 => conv_std_logic_vector(19186, 16),
46443 => conv_std_logic_vector(19367, 16),
46444 => conv_std_logic_vector(19548, 16),
46445 => conv_std_logic_vector(19729, 16),
46446 => conv_std_logic_vector(19910, 16),
46447 => conv_std_logic_vector(20091, 16),
46448 => conv_std_logic_vector(20272, 16),
46449 => conv_std_logic_vector(20453, 16),
46450 => conv_std_logic_vector(20634, 16),
46451 => conv_std_logic_vector(20815, 16),
46452 => conv_std_logic_vector(20996, 16),
46453 => conv_std_logic_vector(21177, 16),
46454 => conv_std_logic_vector(21358, 16),
46455 => conv_std_logic_vector(21539, 16),
46456 => conv_std_logic_vector(21720, 16),
46457 => conv_std_logic_vector(21901, 16),
46458 => conv_std_logic_vector(22082, 16),
46459 => conv_std_logic_vector(22263, 16),
46460 => conv_std_logic_vector(22444, 16),
46461 => conv_std_logic_vector(22625, 16),
46462 => conv_std_logic_vector(22806, 16),
46463 => conv_std_logic_vector(22987, 16),
46464 => conv_std_logic_vector(23168, 16),
46465 => conv_std_logic_vector(23349, 16),
46466 => conv_std_logic_vector(23530, 16),
46467 => conv_std_logic_vector(23711, 16),
46468 => conv_std_logic_vector(23892, 16),
46469 => conv_std_logic_vector(24073, 16),
46470 => conv_std_logic_vector(24254, 16),
46471 => conv_std_logic_vector(24435, 16),
46472 => conv_std_logic_vector(24616, 16),
46473 => conv_std_logic_vector(24797, 16),
46474 => conv_std_logic_vector(24978, 16),
46475 => conv_std_logic_vector(25159, 16),
46476 => conv_std_logic_vector(25340, 16),
46477 => conv_std_logic_vector(25521, 16),
46478 => conv_std_logic_vector(25702, 16),
46479 => conv_std_logic_vector(25883, 16),
46480 => conv_std_logic_vector(26064, 16),
46481 => conv_std_logic_vector(26245, 16),
46482 => conv_std_logic_vector(26426, 16),
46483 => conv_std_logic_vector(26607, 16),
46484 => conv_std_logic_vector(26788, 16),
46485 => conv_std_logic_vector(26969, 16),
46486 => conv_std_logic_vector(27150, 16),
46487 => conv_std_logic_vector(27331, 16),
46488 => conv_std_logic_vector(27512, 16),
46489 => conv_std_logic_vector(27693, 16),
46490 => conv_std_logic_vector(27874, 16),
46491 => conv_std_logic_vector(28055, 16),
46492 => conv_std_logic_vector(28236, 16),
46493 => conv_std_logic_vector(28417, 16),
46494 => conv_std_logic_vector(28598, 16),
46495 => conv_std_logic_vector(28779, 16),
46496 => conv_std_logic_vector(28960, 16),
46497 => conv_std_logic_vector(29141, 16),
46498 => conv_std_logic_vector(29322, 16),
46499 => conv_std_logic_vector(29503, 16),
46500 => conv_std_logic_vector(29684, 16),
46501 => conv_std_logic_vector(29865, 16),
46502 => conv_std_logic_vector(30046, 16),
46503 => conv_std_logic_vector(30227, 16),
46504 => conv_std_logic_vector(30408, 16),
46505 => conv_std_logic_vector(30589, 16),
46506 => conv_std_logic_vector(30770, 16),
46507 => conv_std_logic_vector(30951, 16),
46508 => conv_std_logic_vector(31132, 16),
46509 => conv_std_logic_vector(31313, 16),
46510 => conv_std_logic_vector(31494, 16),
46511 => conv_std_logic_vector(31675, 16),
46512 => conv_std_logic_vector(31856, 16),
46513 => conv_std_logic_vector(32037, 16),
46514 => conv_std_logic_vector(32218, 16),
46515 => conv_std_logic_vector(32399, 16),
46516 => conv_std_logic_vector(32580, 16),
46517 => conv_std_logic_vector(32761, 16),
46518 => conv_std_logic_vector(32942, 16),
46519 => conv_std_logic_vector(33123, 16),
46520 => conv_std_logic_vector(33304, 16),
46521 => conv_std_logic_vector(33485, 16),
46522 => conv_std_logic_vector(33666, 16),
46523 => conv_std_logic_vector(33847, 16),
46524 => conv_std_logic_vector(34028, 16),
46525 => conv_std_logic_vector(34209, 16),
46526 => conv_std_logic_vector(34390, 16),
46527 => conv_std_logic_vector(34571, 16),
46528 => conv_std_logic_vector(34752, 16),
46529 => conv_std_logic_vector(34933, 16),
46530 => conv_std_logic_vector(35114, 16),
46531 => conv_std_logic_vector(35295, 16),
46532 => conv_std_logic_vector(35476, 16),
46533 => conv_std_logic_vector(35657, 16),
46534 => conv_std_logic_vector(35838, 16),
46535 => conv_std_logic_vector(36019, 16),
46536 => conv_std_logic_vector(36200, 16),
46537 => conv_std_logic_vector(36381, 16),
46538 => conv_std_logic_vector(36562, 16),
46539 => conv_std_logic_vector(36743, 16),
46540 => conv_std_logic_vector(36924, 16),
46541 => conv_std_logic_vector(37105, 16),
46542 => conv_std_logic_vector(37286, 16),
46543 => conv_std_logic_vector(37467, 16),
46544 => conv_std_logic_vector(37648, 16),
46545 => conv_std_logic_vector(37829, 16),
46546 => conv_std_logic_vector(38010, 16),
46547 => conv_std_logic_vector(38191, 16),
46548 => conv_std_logic_vector(38372, 16),
46549 => conv_std_logic_vector(38553, 16),
46550 => conv_std_logic_vector(38734, 16),
46551 => conv_std_logic_vector(38915, 16),
46552 => conv_std_logic_vector(39096, 16),
46553 => conv_std_logic_vector(39277, 16),
46554 => conv_std_logic_vector(39458, 16),
46555 => conv_std_logic_vector(39639, 16),
46556 => conv_std_logic_vector(39820, 16),
46557 => conv_std_logic_vector(40001, 16),
46558 => conv_std_logic_vector(40182, 16),
46559 => conv_std_logic_vector(40363, 16),
46560 => conv_std_logic_vector(40544, 16),
46561 => conv_std_logic_vector(40725, 16),
46562 => conv_std_logic_vector(40906, 16),
46563 => conv_std_logic_vector(41087, 16),
46564 => conv_std_logic_vector(41268, 16),
46565 => conv_std_logic_vector(41449, 16),
46566 => conv_std_logic_vector(41630, 16),
46567 => conv_std_logic_vector(41811, 16),
46568 => conv_std_logic_vector(41992, 16),
46569 => conv_std_logic_vector(42173, 16),
46570 => conv_std_logic_vector(42354, 16),
46571 => conv_std_logic_vector(42535, 16),
46572 => conv_std_logic_vector(42716, 16),
46573 => conv_std_logic_vector(42897, 16),
46574 => conv_std_logic_vector(43078, 16),
46575 => conv_std_logic_vector(43259, 16),
46576 => conv_std_logic_vector(43440, 16),
46577 => conv_std_logic_vector(43621, 16),
46578 => conv_std_logic_vector(43802, 16),
46579 => conv_std_logic_vector(43983, 16),
46580 => conv_std_logic_vector(44164, 16),
46581 => conv_std_logic_vector(44345, 16),
46582 => conv_std_logic_vector(44526, 16),
46583 => conv_std_logic_vector(44707, 16),
46584 => conv_std_logic_vector(44888, 16),
46585 => conv_std_logic_vector(45069, 16),
46586 => conv_std_logic_vector(45250, 16),
46587 => conv_std_logic_vector(45431, 16),
46588 => conv_std_logic_vector(45612, 16),
46589 => conv_std_logic_vector(45793, 16),
46590 => conv_std_logic_vector(45974, 16),
46591 => conv_std_logic_vector(46155, 16),
46592 => conv_std_logic_vector(0, 16),
46593 => conv_std_logic_vector(182, 16),
46594 => conv_std_logic_vector(364, 16),
46595 => conv_std_logic_vector(546, 16),
46596 => conv_std_logic_vector(728, 16),
46597 => conv_std_logic_vector(910, 16),
46598 => conv_std_logic_vector(1092, 16),
46599 => conv_std_logic_vector(1274, 16),
46600 => conv_std_logic_vector(1456, 16),
46601 => conv_std_logic_vector(1638, 16),
46602 => conv_std_logic_vector(1820, 16),
46603 => conv_std_logic_vector(2002, 16),
46604 => conv_std_logic_vector(2184, 16),
46605 => conv_std_logic_vector(2366, 16),
46606 => conv_std_logic_vector(2548, 16),
46607 => conv_std_logic_vector(2730, 16),
46608 => conv_std_logic_vector(2912, 16),
46609 => conv_std_logic_vector(3094, 16),
46610 => conv_std_logic_vector(3276, 16),
46611 => conv_std_logic_vector(3458, 16),
46612 => conv_std_logic_vector(3640, 16),
46613 => conv_std_logic_vector(3822, 16),
46614 => conv_std_logic_vector(4004, 16),
46615 => conv_std_logic_vector(4186, 16),
46616 => conv_std_logic_vector(4368, 16),
46617 => conv_std_logic_vector(4550, 16),
46618 => conv_std_logic_vector(4732, 16),
46619 => conv_std_logic_vector(4914, 16),
46620 => conv_std_logic_vector(5096, 16),
46621 => conv_std_logic_vector(5278, 16),
46622 => conv_std_logic_vector(5460, 16),
46623 => conv_std_logic_vector(5642, 16),
46624 => conv_std_logic_vector(5824, 16),
46625 => conv_std_logic_vector(6006, 16),
46626 => conv_std_logic_vector(6188, 16),
46627 => conv_std_logic_vector(6370, 16),
46628 => conv_std_logic_vector(6552, 16),
46629 => conv_std_logic_vector(6734, 16),
46630 => conv_std_logic_vector(6916, 16),
46631 => conv_std_logic_vector(7098, 16),
46632 => conv_std_logic_vector(7280, 16),
46633 => conv_std_logic_vector(7462, 16),
46634 => conv_std_logic_vector(7644, 16),
46635 => conv_std_logic_vector(7826, 16),
46636 => conv_std_logic_vector(8008, 16),
46637 => conv_std_logic_vector(8190, 16),
46638 => conv_std_logic_vector(8372, 16),
46639 => conv_std_logic_vector(8554, 16),
46640 => conv_std_logic_vector(8736, 16),
46641 => conv_std_logic_vector(8918, 16),
46642 => conv_std_logic_vector(9100, 16),
46643 => conv_std_logic_vector(9282, 16),
46644 => conv_std_logic_vector(9464, 16),
46645 => conv_std_logic_vector(9646, 16),
46646 => conv_std_logic_vector(9828, 16),
46647 => conv_std_logic_vector(10010, 16),
46648 => conv_std_logic_vector(10192, 16),
46649 => conv_std_logic_vector(10374, 16),
46650 => conv_std_logic_vector(10556, 16),
46651 => conv_std_logic_vector(10738, 16),
46652 => conv_std_logic_vector(10920, 16),
46653 => conv_std_logic_vector(11102, 16),
46654 => conv_std_logic_vector(11284, 16),
46655 => conv_std_logic_vector(11466, 16),
46656 => conv_std_logic_vector(11648, 16),
46657 => conv_std_logic_vector(11830, 16),
46658 => conv_std_logic_vector(12012, 16),
46659 => conv_std_logic_vector(12194, 16),
46660 => conv_std_logic_vector(12376, 16),
46661 => conv_std_logic_vector(12558, 16),
46662 => conv_std_logic_vector(12740, 16),
46663 => conv_std_logic_vector(12922, 16),
46664 => conv_std_logic_vector(13104, 16),
46665 => conv_std_logic_vector(13286, 16),
46666 => conv_std_logic_vector(13468, 16),
46667 => conv_std_logic_vector(13650, 16),
46668 => conv_std_logic_vector(13832, 16),
46669 => conv_std_logic_vector(14014, 16),
46670 => conv_std_logic_vector(14196, 16),
46671 => conv_std_logic_vector(14378, 16),
46672 => conv_std_logic_vector(14560, 16),
46673 => conv_std_logic_vector(14742, 16),
46674 => conv_std_logic_vector(14924, 16),
46675 => conv_std_logic_vector(15106, 16),
46676 => conv_std_logic_vector(15288, 16),
46677 => conv_std_logic_vector(15470, 16),
46678 => conv_std_logic_vector(15652, 16),
46679 => conv_std_logic_vector(15834, 16),
46680 => conv_std_logic_vector(16016, 16),
46681 => conv_std_logic_vector(16198, 16),
46682 => conv_std_logic_vector(16380, 16),
46683 => conv_std_logic_vector(16562, 16),
46684 => conv_std_logic_vector(16744, 16),
46685 => conv_std_logic_vector(16926, 16),
46686 => conv_std_logic_vector(17108, 16),
46687 => conv_std_logic_vector(17290, 16),
46688 => conv_std_logic_vector(17472, 16),
46689 => conv_std_logic_vector(17654, 16),
46690 => conv_std_logic_vector(17836, 16),
46691 => conv_std_logic_vector(18018, 16),
46692 => conv_std_logic_vector(18200, 16),
46693 => conv_std_logic_vector(18382, 16),
46694 => conv_std_logic_vector(18564, 16),
46695 => conv_std_logic_vector(18746, 16),
46696 => conv_std_logic_vector(18928, 16),
46697 => conv_std_logic_vector(19110, 16),
46698 => conv_std_logic_vector(19292, 16),
46699 => conv_std_logic_vector(19474, 16),
46700 => conv_std_logic_vector(19656, 16),
46701 => conv_std_logic_vector(19838, 16),
46702 => conv_std_logic_vector(20020, 16),
46703 => conv_std_logic_vector(20202, 16),
46704 => conv_std_logic_vector(20384, 16),
46705 => conv_std_logic_vector(20566, 16),
46706 => conv_std_logic_vector(20748, 16),
46707 => conv_std_logic_vector(20930, 16),
46708 => conv_std_logic_vector(21112, 16),
46709 => conv_std_logic_vector(21294, 16),
46710 => conv_std_logic_vector(21476, 16),
46711 => conv_std_logic_vector(21658, 16),
46712 => conv_std_logic_vector(21840, 16),
46713 => conv_std_logic_vector(22022, 16),
46714 => conv_std_logic_vector(22204, 16),
46715 => conv_std_logic_vector(22386, 16),
46716 => conv_std_logic_vector(22568, 16),
46717 => conv_std_logic_vector(22750, 16),
46718 => conv_std_logic_vector(22932, 16),
46719 => conv_std_logic_vector(23114, 16),
46720 => conv_std_logic_vector(23296, 16),
46721 => conv_std_logic_vector(23478, 16),
46722 => conv_std_logic_vector(23660, 16),
46723 => conv_std_logic_vector(23842, 16),
46724 => conv_std_logic_vector(24024, 16),
46725 => conv_std_logic_vector(24206, 16),
46726 => conv_std_logic_vector(24388, 16),
46727 => conv_std_logic_vector(24570, 16),
46728 => conv_std_logic_vector(24752, 16),
46729 => conv_std_logic_vector(24934, 16),
46730 => conv_std_logic_vector(25116, 16),
46731 => conv_std_logic_vector(25298, 16),
46732 => conv_std_logic_vector(25480, 16),
46733 => conv_std_logic_vector(25662, 16),
46734 => conv_std_logic_vector(25844, 16),
46735 => conv_std_logic_vector(26026, 16),
46736 => conv_std_logic_vector(26208, 16),
46737 => conv_std_logic_vector(26390, 16),
46738 => conv_std_logic_vector(26572, 16),
46739 => conv_std_logic_vector(26754, 16),
46740 => conv_std_logic_vector(26936, 16),
46741 => conv_std_logic_vector(27118, 16),
46742 => conv_std_logic_vector(27300, 16),
46743 => conv_std_logic_vector(27482, 16),
46744 => conv_std_logic_vector(27664, 16),
46745 => conv_std_logic_vector(27846, 16),
46746 => conv_std_logic_vector(28028, 16),
46747 => conv_std_logic_vector(28210, 16),
46748 => conv_std_logic_vector(28392, 16),
46749 => conv_std_logic_vector(28574, 16),
46750 => conv_std_logic_vector(28756, 16),
46751 => conv_std_logic_vector(28938, 16),
46752 => conv_std_logic_vector(29120, 16),
46753 => conv_std_logic_vector(29302, 16),
46754 => conv_std_logic_vector(29484, 16),
46755 => conv_std_logic_vector(29666, 16),
46756 => conv_std_logic_vector(29848, 16),
46757 => conv_std_logic_vector(30030, 16),
46758 => conv_std_logic_vector(30212, 16),
46759 => conv_std_logic_vector(30394, 16),
46760 => conv_std_logic_vector(30576, 16),
46761 => conv_std_logic_vector(30758, 16),
46762 => conv_std_logic_vector(30940, 16),
46763 => conv_std_logic_vector(31122, 16),
46764 => conv_std_logic_vector(31304, 16),
46765 => conv_std_logic_vector(31486, 16),
46766 => conv_std_logic_vector(31668, 16),
46767 => conv_std_logic_vector(31850, 16),
46768 => conv_std_logic_vector(32032, 16),
46769 => conv_std_logic_vector(32214, 16),
46770 => conv_std_logic_vector(32396, 16),
46771 => conv_std_logic_vector(32578, 16),
46772 => conv_std_logic_vector(32760, 16),
46773 => conv_std_logic_vector(32942, 16),
46774 => conv_std_logic_vector(33124, 16),
46775 => conv_std_logic_vector(33306, 16),
46776 => conv_std_logic_vector(33488, 16),
46777 => conv_std_logic_vector(33670, 16),
46778 => conv_std_logic_vector(33852, 16),
46779 => conv_std_logic_vector(34034, 16),
46780 => conv_std_logic_vector(34216, 16),
46781 => conv_std_logic_vector(34398, 16),
46782 => conv_std_logic_vector(34580, 16),
46783 => conv_std_logic_vector(34762, 16),
46784 => conv_std_logic_vector(34944, 16),
46785 => conv_std_logic_vector(35126, 16),
46786 => conv_std_logic_vector(35308, 16),
46787 => conv_std_logic_vector(35490, 16),
46788 => conv_std_logic_vector(35672, 16),
46789 => conv_std_logic_vector(35854, 16),
46790 => conv_std_logic_vector(36036, 16),
46791 => conv_std_logic_vector(36218, 16),
46792 => conv_std_logic_vector(36400, 16),
46793 => conv_std_logic_vector(36582, 16),
46794 => conv_std_logic_vector(36764, 16),
46795 => conv_std_logic_vector(36946, 16),
46796 => conv_std_logic_vector(37128, 16),
46797 => conv_std_logic_vector(37310, 16),
46798 => conv_std_logic_vector(37492, 16),
46799 => conv_std_logic_vector(37674, 16),
46800 => conv_std_logic_vector(37856, 16),
46801 => conv_std_logic_vector(38038, 16),
46802 => conv_std_logic_vector(38220, 16),
46803 => conv_std_logic_vector(38402, 16),
46804 => conv_std_logic_vector(38584, 16),
46805 => conv_std_logic_vector(38766, 16),
46806 => conv_std_logic_vector(38948, 16),
46807 => conv_std_logic_vector(39130, 16),
46808 => conv_std_logic_vector(39312, 16),
46809 => conv_std_logic_vector(39494, 16),
46810 => conv_std_logic_vector(39676, 16),
46811 => conv_std_logic_vector(39858, 16),
46812 => conv_std_logic_vector(40040, 16),
46813 => conv_std_logic_vector(40222, 16),
46814 => conv_std_logic_vector(40404, 16),
46815 => conv_std_logic_vector(40586, 16),
46816 => conv_std_logic_vector(40768, 16),
46817 => conv_std_logic_vector(40950, 16),
46818 => conv_std_logic_vector(41132, 16),
46819 => conv_std_logic_vector(41314, 16),
46820 => conv_std_logic_vector(41496, 16),
46821 => conv_std_logic_vector(41678, 16),
46822 => conv_std_logic_vector(41860, 16),
46823 => conv_std_logic_vector(42042, 16),
46824 => conv_std_logic_vector(42224, 16),
46825 => conv_std_logic_vector(42406, 16),
46826 => conv_std_logic_vector(42588, 16),
46827 => conv_std_logic_vector(42770, 16),
46828 => conv_std_logic_vector(42952, 16),
46829 => conv_std_logic_vector(43134, 16),
46830 => conv_std_logic_vector(43316, 16),
46831 => conv_std_logic_vector(43498, 16),
46832 => conv_std_logic_vector(43680, 16),
46833 => conv_std_logic_vector(43862, 16),
46834 => conv_std_logic_vector(44044, 16),
46835 => conv_std_logic_vector(44226, 16),
46836 => conv_std_logic_vector(44408, 16),
46837 => conv_std_logic_vector(44590, 16),
46838 => conv_std_logic_vector(44772, 16),
46839 => conv_std_logic_vector(44954, 16),
46840 => conv_std_logic_vector(45136, 16),
46841 => conv_std_logic_vector(45318, 16),
46842 => conv_std_logic_vector(45500, 16),
46843 => conv_std_logic_vector(45682, 16),
46844 => conv_std_logic_vector(45864, 16),
46845 => conv_std_logic_vector(46046, 16),
46846 => conv_std_logic_vector(46228, 16),
46847 => conv_std_logic_vector(46410, 16),
46848 => conv_std_logic_vector(0, 16),
46849 => conv_std_logic_vector(183, 16),
46850 => conv_std_logic_vector(366, 16),
46851 => conv_std_logic_vector(549, 16),
46852 => conv_std_logic_vector(732, 16),
46853 => conv_std_logic_vector(915, 16),
46854 => conv_std_logic_vector(1098, 16),
46855 => conv_std_logic_vector(1281, 16),
46856 => conv_std_logic_vector(1464, 16),
46857 => conv_std_logic_vector(1647, 16),
46858 => conv_std_logic_vector(1830, 16),
46859 => conv_std_logic_vector(2013, 16),
46860 => conv_std_logic_vector(2196, 16),
46861 => conv_std_logic_vector(2379, 16),
46862 => conv_std_logic_vector(2562, 16),
46863 => conv_std_logic_vector(2745, 16),
46864 => conv_std_logic_vector(2928, 16),
46865 => conv_std_logic_vector(3111, 16),
46866 => conv_std_logic_vector(3294, 16),
46867 => conv_std_logic_vector(3477, 16),
46868 => conv_std_logic_vector(3660, 16),
46869 => conv_std_logic_vector(3843, 16),
46870 => conv_std_logic_vector(4026, 16),
46871 => conv_std_logic_vector(4209, 16),
46872 => conv_std_logic_vector(4392, 16),
46873 => conv_std_logic_vector(4575, 16),
46874 => conv_std_logic_vector(4758, 16),
46875 => conv_std_logic_vector(4941, 16),
46876 => conv_std_logic_vector(5124, 16),
46877 => conv_std_logic_vector(5307, 16),
46878 => conv_std_logic_vector(5490, 16),
46879 => conv_std_logic_vector(5673, 16),
46880 => conv_std_logic_vector(5856, 16),
46881 => conv_std_logic_vector(6039, 16),
46882 => conv_std_logic_vector(6222, 16),
46883 => conv_std_logic_vector(6405, 16),
46884 => conv_std_logic_vector(6588, 16),
46885 => conv_std_logic_vector(6771, 16),
46886 => conv_std_logic_vector(6954, 16),
46887 => conv_std_logic_vector(7137, 16),
46888 => conv_std_logic_vector(7320, 16),
46889 => conv_std_logic_vector(7503, 16),
46890 => conv_std_logic_vector(7686, 16),
46891 => conv_std_logic_vector(7869, 16),
46892 => conv_std_logic_vector(8052, 16),
46893 => conv_std_logic_vector(8235, 16),
46894 => conv_std_logic_vector(8418, 16),
46895 => conv_std_logic_vector(8601, 16),
46896 => conv_std_logic_vector(8784, 16),
46897 => conv_std_logic_vector(8967, 16),
46898 => conv_std_logic_vector(9150, 16),
46899 => conv_std_logic_vector(9333, 16),
46900 => conv_std_logic_vector(9516, 16),
46901 => conv_std_logic_vector(9699, 16),
46902 => conv_std_logic_vector(9882, 16),
46903 => conv_std_logic_vector(10065, 16),
46904 => conv_std_logic_vector(10248, 16),
46905 => conv_std_logic_vector(10431, 16),
46906 => conv_std_logic_vector(10614, 16),
46907 => conv_std_logic_vector(10797, 16),
46908 => conv_std_logic_vector(10980, 16),
46909 => conv_std_logic_vector(11163, 16),
46910 => conv_std_logic_vector(11346, 16),
46911 => conv_std_logic_vector(11529, 16),
46912 => conv_std_logic_vector(11712, 16),
46913 => conv_std_logic_vector(11895, 16),
46914 => conv_std_logic_vector(12078, 16),
46915 => conv_std_logic_vector(12261, 16),
46916 => conv_std_logic_vector(12444, 16),
46917 => conv_std_logic_vector(12627, 16),
46918 => conv_std_logic_vector(12810, 16),
46919 => conv_std_logic_vector(12993, 16),
46920 => conv_std_logic_vector(13176, 16),
46921 => conv_std_logic_vector(13359, 16),
46922 => conv_std_logic_vector(13542, 16),
46923 => conv_std_logic_vector(13725, 16),
46924 => conv_std_logic_vector(13908, 16),
46925 => conv_std_logic_vector(14091, 16),
46926 => conv_std_logic_vector(14274, 16),
46927 => conv_std_logic_vector(14457, 16),
46928 => conv_std_logic_vector(14640, 16),
46929 => conv_std_logic_vector(14823, 16),
46930 => conv_std_logic_vector(15006, 16),
46931 => conv_std_logic_vector(15189, 16),
46932 => conv_std_logic_vector(15372, 16),
46933 => conv_std_logic_vector(15555, 16),
46934 => conv_std_logic_vector(15738, 16),
46935 => conv_std_logic_vector(15921, 16),
46936 => conv_std_logic_vector(16104, 16),
46937 => conv_std_logic_vector(16287, 16),
46938 => conv_std_logic_vector(16470, 16),
46939 => conv_std_logic_vector(16653, 16),
46940 => conv_std_logic_vector(16836, 16),
46941 => conv_std_logic_vector(17019, 16),
46942 => conv_std_logic_vector(17202, 16),
46943 => conv_std_logic_vector(17385, 16),
46944 => conv_std_logic_vector(17568, 16),
46945 => conv_std_logic_vector(17751, 16),
46946 => conv_std_logic_vector(17934, 16),
46947 => conv_std_logic_vector(18117, 16),
46948 => conv_std_logic_vector(18300, 16),
46949 => conv_std_logic_vector(18483, 16),
46950 => conv_std_logic_vector(18666, 16),
46951 => conv_std_logic_vector(18849, 16),
46952 => conv_std_logic_vector(19032, 16),
46953 => conv_std_logic_vector(19215, 16),
46954 => conv_std_logic_vector(19398, 16),
46955 => conv_std_logic_vector(19581, 16),
46956 => conv_std_logic_vector(19764, 16),
46957 => conv_std_logic_vector(19947, 16),
46958 => conv_std_logic_vector(20130, 16),
46959 => conv_std_logic_vector(20313, 16),
46960 => conv_std_logic_vector(20496, 16),
46961 => conv_std_logic_vector(20679, 16),
46962 => conv_std_logic_vector(20862, 16),
46963 => conv_std_logic_vector(21045, 16),
46964 => conv_std_logic_vector(21228, 16),
46965 => conv_std_logic_vector(21411, 16),
46966 => conv_std_logic_vector(21594, 16),
46967 => conv_std_logic_vector(21777, 16),
46968 => conv_std_logic_vector(21960, 16),
46969 => conv_std_logic_vector(22143, 16),
46970 => conv_std_logic_vector(22326, 16),
46971 => conv_std_logic_vector(22509, 16),
46972 => conv_std_logic_vector(22692, 16),
46973 => conv_std_logic_vector(22875, 16),
46974 => conv_std_logic_vector(23058, 16),
46975 => conv_std_logic_vector(23241, 16),
46976 => conv_std_logic_vector(23424, 16),
46977 => conv_std_logic_vector(23607, 16),
46978 => conv_std_logic_vector(23790, 16),
46979 => conv_std_logic_vector(23973, 16),
46980 => conv_std_logic_vector(24156, 16),
46981 => conv_std_logic_vector(24339, 16),
46982 => conv_std_logic_vector(24522, 16),
46983 => conv_std_logic_vector(24705, 16),
46984 => conv_std_logic_vector(24888, 16),
46985 => conv_std_logic_vector(25071, 16),
46986 => conv_std_logic_vector(25254, 16),
46987 => conv_std_logic_vector(25437, 16),
46988 => conv_std_logic_vector(25620, 16),
46989 => conv_std_logic_vector(25803, 16),
46990 => conv_std_logic_vector(25986, 16),
46991 => conv_std_logic_vector(26169, 16),
46992 => conv_std_logic_vector(26352, 16),
46993 => conv_std_logic_vector(26535, 16),
46994 => conv_std_logic_vector(26718, 16),
46995 => conv_std_logic_vector(26901, 16),
46996 => conv_std_logic_vector(27084, 16),
46997 => conv_std_logic_vector(27267, 16),
46998 => conv_std_logic_vector(27450, 16),
46999 => conv_std_logic_vector(27633, 16),
47000 => conv_std_logic_vector(27816, 16),
47001 => conv_std_logic_vector(27999, 16),
47002 => conv_std_logic_vector(28182, 16),
47003 => conv_std_logic_vector(28365, 16),
47004 => conv_std_logic_vector(28548, 16),
47005 => conv_std_logic_vector(28731, 16),
47006 => conv_std_logic_vector(28914, 16),
47007 => conv_std_logic_vector(29097, 16),
47008 => conv_std_logic_vector(29280, 16),
47009 => conv_std_logic_vector(29463, 16),
47010 => conv_std_logic_vector(29646, 16),
47011 => conv_std_logic_vector(29829, 16),
47012 => conv_std_logic_vector(30012, 16),
47013 => conv_std_logic_vector(30195, 16),
47014 => conv_std_logic_vector(30378, 16),
47015 => conv_std_logic_vector(30561, 16),
47016 => conv_std_logic_vector(30744, 16),
47017 => conv_std_logic_vector(30927, 16),
47018 => conv_std_logic_vector(31110, 16),
47019 => conv_std_logic_vector(31293, 16),
47020 => conv_std_logic_vector(31476, 16),
47021 => conv_std_logic_vector(31659, 16),
47022 => conv_std_logic_vector(31842, 16),
47023 => conv_std_logic_vector(32025, 16),
47024 => conv_std_logic_vector(32208, 16),
47025 => conv_std_logic_vector(32391, 16),
47026 => conv_std_logic_vector(32574, 16),
47027 => conv_std_logic_vector(32757, 16),
47028 => conv_std_logic_vector(32940, 16),
47029 => conv_std_logic_vector(33123, 16),
47030 => conv_std_logic_vector(33306, 16),
47031 => conv_std_logic_vector(33489, 16),
47032 => conv_std_logic_vector(33672, 16),
47033 => conv_std_logic_vector(33855, 16),
47034 => conv_std_logic_vector(34038, 16),
47035 => conv_std_logic_vector(34221, 16),
47036 => conv_std_logic_vector(34404, 16),
47037 => conv_std_logic_vector(34587, 16),
47038 => conv_std_logic_vector(34770, 16),
47039 => conv_std_logic_vector(34953, 16),
47040 => conv_std_logic_vector(35136, 16),
47041 => conv_std_logic_vector(35319, 16),
47042 => conv_std_logic_vector(35502, 16),
47043 => conv_std_logic_vector(35685, 16),
47044 => conv_std_logic_vector(35868, 16),
47045 => conv_std_logic_vector(36051, 16),
47046 => conv_std_logic_vector(36234, 16),
47047 => conv_std_logic_vector(36417, 16),
47048 => conv_std_logic_vector(36600, 16),
47049 => conv_std_logic_vector(36783, 16),
47050 => conv_std_logic_vector(36966, 16),
47051 => conv_std_logic_vector(37149, 16),
47052 => conv_std_logic_vector(37332, 16),
47053 => conv_std_logic_vector(37515, 16),
47054 => conv_std_logic_vector(37698, 16),
47055 => conv_std_logic_vector(37881, 16),
47056 => conv_std_logic_vector(38064, 16),
47057 => conv_std_logic_vector(38247, 16),
47058 => conv_std_logic_vector(38430, 16),
47059 => conv_std_logic_vector(38613, 16),
47060 => conv_std_logic_vector(38796, 16),
47061 => conv_std_logic_vector(38979, 16),
47062 => conv_std_logic_vector(39162, 16),
47063 => conv_std_logic_vector(39345, 16),
47064 => conv_std_logic_vector(39528, 16),
47065 => conv_std_logic_vector(39711, 16),
47066 => conv_std_logic_vector(39894, 16),
47067 => conv_std_logic_vector(40077, 16),
47068 => conv_std_logic_vector(40260, 16),
47069 => conv_std_logic_vector(40443, 16),
47070 => conv_std_logic_vector(40626, 16),
47071 => conv_std_logic_vector(40809, 16),
47072 => conv_std_logic_vector(40992, 16),
47073 => conv_std_logic_vector(41175, 16),
47074 => conv_std_logic_vector(41358, 16),
47075 => conv_std_logic_vector(41541, 16),
47076 => conv_std_logic_vector(41724, 16),
47077 => conv_std_logic_vector(41907, 16),
47078 => conv_std_logic_vector(42090, 16),
47079 => conv_std_logic_vector(42273, 16),
47080 => conv_std_logic_vector(42456, 16),
47081 => conv_std_logic_vector(42639, 16),
47082 => conv_std_logic_vector(42822, 16),
47083 => conv_std_logic_vector(43005, 16),
47084 => conv_std_logic_vector(43188, 16),
47085 => conv_std_logic_vector(43371, 16),
47086 => conv_std_logic_vector(43554, 16),
47087 => conv_std_logic_vector(43737, 16),
47088 => conv_std_logic_vector(43920, 16),
47089 => conv_std_logic_vector(44103, 16),
47090 => conv_std_logic_vector(44286, 16),
47091 => conv_std_logic_vector(44469, 16),
47092 => conv_std_logic_vector(44652, 16),
47093 => conv_std_logic_vector(44835, 16),
47094 => conv_std_logic_vector(45018, 16),
47095 => conv_std_logic_vector(45201, 16),
47096 => conv_std_logic_vector(45384, 16),
47097 => conv_std_logic_vector(45567, 16),
47098 => conv_std_logic_vector(45750, 16),
47099 => conv_std_logic_vector(45933, 16),
47100 => conv_std_logic_vector(46116, 16),
47101 => conv_std_logic_vector(46299, 16),
47102 => conv_std_logic_vector(46482, 16),
47103 => conv_std_logic_vector(46665, 16),
47104 => conv_std_logic_vector(0, 16),
47105 => conv_std_logic_vector(184, 16),
47106 => conv_std_logic_vector(368, 16),
47107 => conv_std_logic_vector(552, 16),
47108 => conv_std_logic_vector(736, 16),
47109 => conv_std_logic_vector(920, 16),
47110 => conv_std_logic_vector(1104, 16),
47111 => conv_std_logic_vector(1288, 16),
47112 => conv_std_logic_vector(1472, 16),
47113 => conv_std_logic_vector(1656, 16),
47114 => conv_std_logic_vector(1840, 16),
47115 => conv_std_logic_vector(2024, 16),
47116 => conv_std_logic_vector(2208, 16),
47117 => conv_std_logic_vector(2392, 16),
47118 => conv_std_logic_vector(2576, 16),
47119 => conv_std_logic_vector(2760, 16),
47120 => conv_std_logic_vector(2944, 16),
47121 => conv_std_logic_vector(3128, 16),
47122 => conv_std_logic_vector(3312, 16),
47123 => conv_std_logic_vector(3496, 16),
47124 => conv_std_logic_vector(3680, 16),
47125 => conv_std_logic_vector(3864, 16),
47126 => conv_std_logic_vector(4048, 16),
47127 => conv_std_logic_vector(4232, 16),
47128 => conv_std_logic_vector(4416, 16),
47129 => conv_std_logic_vector(4600, 16),
47130 => conv_std_logic_vector(4784, 16),
47131 => conv_std_logic_vector(4968, 16),
47132 => conv_std_logic_vector(5152, 16),
47133 => conv_std_logic_vector(5336, 16),
47134 => conv_std_logic_vector(5520, 16),
47135 => conv_std_logic_vector(5704, 16),
47136 => conv_std_logic_vector(5888, 16),
47137 => conv_std_logic_vector(6072, 16),
47138 => conv_std_logic_vector(6256, 16),
47139 => conv_std_logic_vector(6440, 16),
47140 => conv_std_logic_vector(6624, 16),
47141 => conv_std_logic_vector(6808, 16),
47142 => conv_std_logic_vector(6992, 16),
47143 => conv_std_logic_vector(7176, 16),
47144 => conv_std_logic_vector(7360, 16),
47145 => conv_std_logic_vector(7544, 16),
47146 => conv_std_logic_vector(7728, 16),
47147 => conv_std_logic_vector(7912, 16),
47148 => conv_std_logic_vector(8096, 16),
47149 => conv_std_logic_vector(8280, 16),
47150 => conv_std_logic_vector(8464, 16),
47151 => conv_std_logic_vector(8648, 16),
47152 => conv_std_logic_vector(8832, 16),
47153 => conv_std_logic_vector(9016, 16),
47154 => conv_std_logic_vector(9200, 16),
47155 => conv_std_logic_vector(9384, 16),
47156 => conv_std_logic_vector(9568, 16),
47157 => conv_std_logic_vector(9752, 16),
47158 => conv_std_logic_vector(9936, 16),
47159 => conv_std_logic_vector(10120, 16),
47160 => conv_std_logic_vector(10304, 16),
47161 => conv_std_logic_vector(10488, 16),
47162 => conv_std_logic_vector(10672, 16),
47163 => conv_std_logic_vector(10856, 16),
47164 => conv_std_logic_vector(11040, 16),
47165 => conv_std_logic_vector(11224, 16),
47166 => conv_std_logic_vector(11408, 16),
47167 => conv_std_logic_vector(11592, 16),
47168 => conv_std_logic_vector(11776, 16),
47169 => conv_std_logic_vector(11960, 16),
47170 => conv_std_logic_vector(12144, 16),
47171 => conv_std_logic_vector(12328, 16),
47172 => conv_std_logic_vector(12512, 16),
47173 => conv_std_logic_vector(12696, 16),
47174 => conv_std_logic_vector(12880, 16),
47175 => conv_std_logic_vector(13064, 16),
47176 => conv_std_logic_vector(13248, 16),
47177 => conv_std_logic_vector(13432, 16),
47178 => conv_std_logic_vector(13616, 16),
47179 => conv_std_logic_vector(13800, 16),
47180 => conv_std_logic_vector(13984, 16),
47181 => conv_std_logic_vector(14168, 16),
47182 => conv_std_logic_vector(14352, 16),
47183 => conv_std_logic_vector(14536, 16),
47184 => conv_std_logic_vector(14720, 16),
47185 => conv_std_logic_vector(14904, 16),
47186 => conv_std_logic_vector(15088, 16),
47187 => conv_std_logic_vector(15272, 16),
47188 => conv_std_logic_vector(15456, 16),
47189 => conv_std_logic_vector(15640, 16),
47190 => conv_std_logic_vector(15824, 16),
47191 => conv_std_logic_vector(16008, 16),
47192 => conv_std_logic_vector(16192, 16),
47193 => conv_std_logic_vector(16376, 16),
47194 => conv_std_logic_vector(16560, 16),
47195 => conv_std_logic_vector(16744, 16),
47196 => conv_std_logic_vector(16928, 16),
47197 => conv_std_logic_vector(17112, 16),
47198 => conv_std_logic_vector(17296, 16),
47199 => conv_std_logic_vector(17480, 16),
47200 => conv_std_logic_vector(17664, 16),
47201 => conv_std_logic_vector(17848, 16),
47202 => conv_std_logic_vector(18032, 16),
47203 => conv_std_logic_vector(18216, 16),
47204 => conv_std_logic_vector(18400, 16),
47205 => conv_std_logic_vector(18584, 16),
47206 => conv_std_logic_vector(18768, 16),
47207 => conv_std_logic_vector(18952, 16),
47208 => conv_std_logic_vector(19136, 16),
47209 => conv_std_logic_vector(19320, 16),
47210 => conv_std_logic_vector(19504, 16),
47211 => conv_std_logic_vector(19688, 16),
47212 => conv_std_logic_vector(19872, 16),
47213 => conv_std_logic_vector(20056, 16),
47214 => conv_std_logic_vector(20240, 16),
47215 => conv_std_logic_vector(20424, 16),
47216 => conv_std_logic_vector(20608, 16),
47217 => conv_std_logic_vector(20792, 16),
47218 => conv_std_logic_vector(20976, 16),
47219 => conv_std_logic_vector(21160, 16),
47220 => conv_std_logic_vector(21344, 16),
47221 => conv_std_logic_vector(21528, 16),
47222 => conv_std_logic_vector(21712, 16),
47223 => conv_std_logic_vector(21896, 16),
47224 => conv_std_logic_vector(22080, 16),
47225 => conv_std_logic_vector(22264, 16),
47226 => conv_std_logic_vector(22448, 16),
47227 => conv_std_logic_vector(22632, 16),
47228 => conv_std_logic_vector(22816, 16),
47229 => conv_std_logic_vector(23000, 16),
47230 => conv_std_logic_vector(23184, 16),
47231 => conv_std_logic_vector(23368, 16),
47232 => conv_std_logic_vector(23552, 16),
47233 => conv_std_logic_vector(23736, 16),
47234 => conv_std_logic_vector(23920, 16),
47235 => conv_std_logic_vector(24104, 16),
47236 => conv_std_logic_vector(24288, 16),
47237 => conv_std_logic_vector(24472, 16),
47238 => conv_std_logic_vector(24656, 16),
47239 => conv_std_logic_vector(24840, 16),
47240 => conv_std_logic_vector(25024, 16),
47241 => conv_std_logic_vector(25208, 16),
47242 => conv_std_logic_vector(25392, 16),
47243 => conv_std_logic_vector(25576, 16),
47244 => conv_std_logic_vector(25760, 16),
47245 => conv_std_logic_vector(25944, 16),
47246 => conv_std_logic_vector(26128, 16),
47247 => conv_std_logic_vector(26312, 16),
47248 => conv_std_logic_vector(26496, 16),
47249 => conv_std_logic_vector(26680, 16),
47250 => conv_std_logic_vector(26864, 16),
47251 => conv_std_logic_vector(27048, 16),
47252 => conv_std_logic_vector(27232, 16),
47253 => conv_std_logic_vector(27416, 16),
47254 => conv_std_logic_vector(27600, 16),
47255 => conv_std_logic_vector(27784, 16),
47256 => conv_std_logic_vector(27968, 16),
47257 => conv_std_logic_vector(28152, 16),
47258 => conv_std_logic_vector(28336, 16),
47259 => conv_std_logic_vector(28520, 16),
47260 => conv_std_logic_vector(28704, 16),
47261 => conv_std_logic_vector(28888, 16),
47262 => conv_std_logic_vector(29072, 16),
47263 => conv_std_logic_vector(29256, 16),
47264 => conv_std_logic_vector(29440, 16),
47265 => conv_std_logic_vector(29624, 16),
47266 => conv_std_logic_vector(29808, 16),
47267 => conv_std_logic_vector(29992, 16),
47268 => conv_std_logic_vector(30176, 16),
47269 => conv_std_logic_vector(30360, 16),
47270 => conv_std_logic_vector(30544, 16),
47271 => conv_std_logic_vector(30728, 16),
47272 => conv_std_logic_vector(30912, 16),
47273 => conv_std_logic_vector(31096, 16),
47274 => conv_std_logic_vector(31280, 16),
47275 => conv_std_logic_vector(31464, 16),
47276 => conv_std_logic_vector(31648, 16),
47277 => conv_std_logic_vector(31832, 16),
47278 => conv_std_logic_vector(32016, 16),
47279 => conv_std_logic_vector(32200, 16),
47280 => conv_std_logic_vector(32384, 16),
47281 => conv_std_logic_vector(32568, 16),
47282 => conv_std_logic_vector(32752, 16),
47283 => conv_std_logic_vector(32936, 16),
47284 => conv_std_logic_vector(33120, 16),
47285 => conv_std_logic_vector(33304, 16),
47286 => conv_std_logic_vector(33488, 16),
47287 => conv_std_logic_vector(33672, 16),
47288 => conv_std_logic_vector(33856, 16),
47289 => conv_std_logic_vector(34040, 16),
47290 => conv_std_logic_vector(34224, 16),
47291 => conv_std_logic_vector(34408, 16),
47292 => conv_std_logic_vector(34592, 16),
47293 => conv_std_logic_vector(34776, 16),
47294 => conv_std_logic_vector(34960, 16),
47295 => conv_std_logic_vector(35144, 16),
47296 => conv_std_logic_vector(35328, 16),
47297 => conv_std_logic_vector(35512, 16),
47298 => conv_std_logic_vector(35696, 16),
47299 => conv_std_logic_vector(35880, 16),
47300 => conv_std_logic_vector(36064, 16),
47301 => conv_std_logic_vector(36248, 16),
47302 => conv_std_logic_vector(36432, 16),
47303 => conv_std_logic_vector(36616, 16),
47304 => conv_std_logic_vector(36800, 16),
47305 => conv_std_logic_vector(36984, 16),
47306 => conv_std_logic_vector(37168, 16),
47307 => conv_std_logic_vector(37352, 16),
47308 => conv_std_logic_vector(37536, 16),
47309 => conv_std_logic_vector(37720, 16),
47310 => conv_std_logic_vector(37904, 16),
47311 => conv_std_logic_vector(38088, 16),
47312 => conv_std_logic_vector(38272, 16),
47313 => conv_std_logic_vector(38456, 16),
47314 => conv_std_logic_vector(38640, 16),
47315 => conv_std_logic_vector(38824, 16),
47316 => conv_std_logic_vector(39008, 16),
47317 => conv_std_logic_vector(39192, 16),
47318 => conv_std_logic_vector(39376, 16),
47319 => conv_std_logic_vector(39560, 16),
47320 => conv_std_logic_vector(39744, 16),
47321 => conv_std_logic_vector(39928, 16),
47322 => conv_std_logic_vector(40112, 16),
47323 => conv_std_logic_vector(40296, 16),
47324 => conv_std_logic_vector(40480, 16),
47325 => conv_std_logic_vector(40664, 16),
47326 => conv_std_logic_vector(40848, 16),
47327 => conv_std_logic_vector(41032, 16),
47328 => conv_std_logic_vector(41216, 16),
47329 => conv_std_logic_vector(41400, 16),
47330 => conv_std_logic_vector(41584, 16),
47331 => conv_std_logic_vector(41768, 16),
47332 => conv_std_logic_vector(41952, 16),
47333 => conv_std_logic_vector(42136, 16),
47334 => conv_std_logic_vector(42320, 16),
47335 => conv_std_logic_vector(42504, 16),
47336 => conv_std_logic_vector(42688, 16),
47337 => conv_std_logic_vector(42872, 16),
47338 => conv_std_logic_vector(43056, 16),
47339 => conv_std_logic_vector(43240, 16),
47340 => conv_std_logic_vector(43424, 16),
47341 => conv_std_logic_vector(43608, 16),
47342 => conv_std_logic_vector(43792, 16),
47343 => conv_std_logic_vector(43976, 16),
47344 => conv_std_logic_vector(44160, 16),
47345 => conv_std_logic_vector(44344, 16),
47346 => conv_std_logic_vector(44528, 16),
47347 => conv_std_logic_vector(44712, 16),
47348 => conv_std_logic_vector(44896, 16),
47349 => conv_std_logic_vector(45080, 16),
47350 => conv_std_logic_vector(45264, 16),
47351 => conv_std_logic_vector(45448, 16),
47352 => conv_std_logic_vector(45632, 16),
47353 => conv_std_logic_vector(45816, 16),
47354 => conv_std_logic_vector(46000, 16),
47355 => conv_std_logic_vector(46184, 16),
47356 => conv_std_logic_vector(46368, 16),
47357 => conv_std_logic_vector(46552, 16),
47358 => conv_std_logic_vector(46736, 16),
47359 => conv_std_logic_vector(46920, 16),
47360 => conv_std_logic_vector(0, 16),
47361 => conv_std_logic_vector(185, 16),
47362 => conv_std_logic_vector(370, 16),
47363 => conv_std_logic_vector(555, 16),
47364 => conv_std_logic_vector(740, 16),
47365 => conv_std_logic_vector(925, 16),
47366 => conv_std_logic_vector(1110, 16),
47367 => conv_std_logic_vector(1295, 16),
47368 => conv_std_logic_vector(1480, 16),
47369 => conv_std_logic_vector(1665, 16),
47370 => conv_std_logic_vector(1850, 16),
47371 => conv_std_logic_vector(2035, 16),
47372 => conv_std_logic_vector(2220, 16),
47373 => conv_std_logic_vector(2405, 16),
47374 => conv_std_logic_vector(2590, 16),
47375 => conv_std_logic_vector(2775, 16),
47376 => conv_std_logic_vector(2960, 16),
47377 => conv_std_logic_vector(3145, 16),
47378 => conv_std_logic_vector(3330, 16),
47379 => conv_std_logic_vector(3515, 16),
47380 => conv_std_logic_vector(3700, 16),
47381 => conv_std_logic_vector(3885, 16),
47382 => conv_std_logic_vector(4070, 16),
47383 => conv_std_logic_vector(4255, 16),
47384 => conv_std_logic_vector(4440, 16),
47385 => conv_std_logic_vector(4625, 16),
47386 => conv_std_logic_vector(4810, 16),
47387 => conv_std_logic_vector(4995, 16),
47388 => conv_std_logic_vector(5180, 16),
47389 => conv_std_logic_vector(5365, 16),
47390 => conv_std_logic_vector(5550, 16),
47391 => conv_std_logic_vector(5735, 16),
47392 => conv_std_logic_vector(5920, 16),
47393 => conv_std_logic_vector(6105, 16),
47394 => conv_std_logic_vector(6290, 16),
47395 => conv_std_logic_vector(6475, 16),
47396 => conv_std_logic_vector(6660, 16),
47397 => conv_std_logic_vector(6845, 16),
47398 => conv_std_logic_vector(7030, 16),
47399 => conv_std_logic_vector(7215, 16),
47400 => conv_std_logic_vector(7400, 16),
47401 => conv_std_logic_vector(7585, 16),
47402 => conv_std_logic_vector(7770, 16),
47403 => conv_std_logic_vector(7955, 16),
47404 => conv_std_logic_vector(8140, 16),
47405 => conv_std_logic_vector(8325, 16),
47406 => conv_std_logic_vector(8510, 16),
47407 => conv_std_logic_vector(8695, 16),
47408 => conv_std_logic_vector(8880, 16),
47409 => conv_std_logic_vector(9065, 16),
47410 => conv_std_logic_vector(9250, 16),
47411 => conv_std_logic_vector(9435, 16),
47412 => conv_std_logic_vector(9620, 16),
47413 => conv_std_logic_vector(9805, 16),
47414 => conv_std_logic_vector(9990, 16),
47415 => conv_std_logic_vector(10175, 16),
47416 => conv_std_logic_vector(10360, 16),
47417 => conv_std_logic_vector(10545, 16),
47418 => conv_std_logic_vector(10730, 16),
47419 => conv_std_logic_vector(10915, 16),
47420 => conv_std_logic_vector(11100, 16),
47421 => conv_std_logic_vector(11285, 16),
47422 => conv_std_logic_vector(11470, 16),
47423 => conv_std_logic_vector(11655, 16),
47424 => conv_std_logic_vector(11840, 16),
47425 => conv_std_logic_vector(12025, 16),
47426 => conv_std_logic_vector(12210, 16),
47427 => conv_std_logic_vector(12395, 16),
47428 => conv_std_logic_vector(12580, 16),
47429 => conv_std_logic_vector(12765, 16),
47430 => conv_std_logic_vector(12950, 16),
47431 => conv_std_logic_vector(13135, 16),
47432 => conv_std_logic_vector(13320, 16),
47433 => conv_std_logic_vector(13505, 16),
47434 => conv_std_logic_vector(13690, 16),
47435 => conv_std_logic_vector(13875, 16),
47436 => conv_std_logic_vector(14060, 16),
47437 => conv_std_logic_vector(14245, 16),
47438 => conv_std_logic_vector(14430, 16),
47439 => conv_std_logic_vector(14615, 16),
47440 => conv_std_logic_vector(14800, 16),
47441 => conv_std_logic_vector(14985, 16),
47442 => conv_std_logic_vector(15170, 16),
47443 => conv_std_logic_vector(15355, 16),
47444 => conv_std_logic_vector(15540, 16),
47445 => conv_std_logic_vector(15725, 16),
47446 => conv_std_logic_vector(15910, 16),
47447 => conv_std_logic_vector(16095, 16),
47448 => conv_std_logic_vector(16280, 16),
47449 => conv_std_logic_vector(16465, 16),
47450 => conv_std_logic_vector(16650, 16),
47451 => conv_std_logic_vector(16835, 16),
47452 => conv_std_logic_vector(17020, 16),
47453 => conv_std_logic_vector(17205, 16),
47454 => conv_std_logic_vector(17390, 16),
47455 => conv_std_logic_vector(17575, 16),
47456 => conv_std_logic_vector(17760, 16),
47457 => conv_std_logic_vector(17945, 16),
47458 => conv_std_logic_vector(18130, 16),
47459 => conv_std_logic_vector(18315, 16),
47460 => conv_std_logic_vector(18500, 16),
47461 => conv_std_logic_vector(18685, 16),
47462 => conv_std_logic_vector(18870, 16),
47463 => conv_std_logic_vector(19055, 16),
47464 => conv_std_logic_vector(19240, 16),
47465 => conv_std_logic_vector(19425, 16),
47466 => conv_std_logic_vector(19610, 16),
47467 => conv_std_logic_vector(19795, 16),
47468 => conv_std_logic_vector(19980, 16),
47469 => conv_std_logic_vector(20165, 16),
47470 => conv_std_logic_vector(20350, 16),
47471 => conv_std_logic_vector(20535, 16),
47472 => conv_std_logic_vector(20720, 16),
47473 => conv_std_logic_vector(20905, 16),
47474 => conv_std_logic_vector(21090, 16),
47475 => conv_std_logic_vector(21275, 16),
47476 => conv_std_logic_vector(21460, 16),
47477 => conv_std_logic_vector(21645, 16),
47478 => conv_std_logic_vector(21830, 16),
47479 => conv_std_logic_vector(22015, 16),
47480 => conv_std_logic_vector(22200, 16),
47481 => conv_std_logic_vector(22385, 16),
47482 => conv_std_logic_vector(22570, 16),
47483 => conv_std_logic_vector(22755, 16),
47484 => conv_std_logic_vector(22940, 16),
47485 => conv_std_logic_vector(23125, 16),
47486 => conv_std_logic_vector(23310, 16),
47487 => conv_std_logic_vector(23495, 16),
47488 => conv_std_logic_vector(23680, 16),
47489 => conv_std_logic_vector(23865, 16),
47490 => conv_std_logic_vector(24050, 16),
47491 => conv_std_logic_vector(24235, 16),
47492 => conv_std_logic_vector(24420, 16),
47493 => conv_std_logic_vector(24605, 16),
47494 => conv_std_logic_vector(24790, 16),
47495 => conv_std_logic_vector(24975, 16),
47496 => conv_std_logic_vector(25160, 16),
47497 => conv_std_logic_vector(25345, 16),
47498 => conv_std_logic_vector(25530, 16),
47499 => conv_std_logic_vector(25715, 16),
47500 => conv_std_logic_vector(25900, 16),
47501 => conv_std_logic_vector(26085, 16),
47502 => conv_std_logic_vector(26270, 16),
47503 => conv_std_logic_vector(26455, 16),
47504 => conv_std_logic_vector(26640, 16),
47505 => conv_std_logic_vector(26825, 16),
47506 => conv_std_logic_vector(27010, 16),
47507 => conv_std_logic_vector(27195, 16),
47508 => conv_std_logic_vector(27380, 16),
47509 => conv_std_logic_vector(27565, 16),
47510 => conv_std_logic_vector(27750, 16),
47511 => conv_std_logic_vector(27935, 16),
47512 => conv_std_logic_vector(28120, 16),
47513 => conv_std_logic_vector(28305, 16),
47514 => conv_std_logic_vector(28490, 16),
47515 => conv_std_logic_vector(28675, 16),
47516 => conv_std_logic_vector(28860, 16),
47517 => conv_std_logic_vector(29045, 16),
47518 => conv_std_logic_vector(29230, 16),
47519 => conv_std_logic_vector(29415, 16),
47520 => conv_std_logic_vector(29600, 16),
47521 => conv_std_logic_vector(29785, 16),
47522 => conv_std_logic_vector(29970, 16),
47523 => conv_std_logic_vector(30155, 16),
47524 => conv_std_logic_vector(30340, 16),
47525 => conv_std_logic_vector(30525, 16),
47526 => conv_std_logic_vector(30710, 16),
47527 => conv_std_logic_vector(30895, 16),
47528 => conv_std_logic_vector(31080, 16),
47529 => conv_std_logic_vector(31265, 16),
47530 => conv_std_logic_vector(31450, 16),
47531 => conv_std_logic_vector(31635, 16),
47532 => conv_std_logic_vector(31820, 16),
47533 => conv_std_logic_vector(32005, 16),
47534 => conv_std_logic_vector(32190, 16),
47535 => conv_std_logic_vector(32375, 16),
47536 => conv_std_logic_vector(32560, 16),
47537 => conv_std_logic_vector(32745, 16),
47538 => conv_std_logic_vector(32930, 16),
47539 => conv_std_logic_vector(33115, 16),
47540 => conv_std_logic_vector(33300, 16),
47541 => conv_std_logic_vector(33485, 16),
47542 => conv_std_logic_vector(33670, 16),
47543 => conv_std_logic_vector(33855, 16),
47544 => conv_std_logic_vector(34040, 16),
47545 => conv_std_logic_vector(34225, 16),
47546 => conv_std_logic_vector(34410, 16),
47547 => conv_std_logic_vector(34595, 16),
47548 => conv_std_logic_vector(34780, 16),
47549 => conv_std_logic_vector(34965, 16),
47550 => conv_std_logic_vector(35150, 16),
47551 => conv_std_logic_vector(35335, 16),
47552 => conv_std_logic_vector(35520, 16),
47553 => conv_std_logic_vector(35705, 16),
47554 => conv_std_logic_vector(35890, 16),
47555 => conv_std_logic_vector(36075, 16),
47556 => conv_std_logic_vector(36260, 16),
47557 => conv_std_logic_vector(36445, 16),
47558 => conv_std_logic_vector(36630, 16),
47559 => conv_std_logic_vector(36815, 16),
47560 => conv_std_logic_vector(37000, 16),
47561 => conv_std_logic_vector(37185, 16),
47562 => conv_std_logic_vector(37370, 16),
47563 => conv_std_logic_vector(37555, 16),
47564 => conv_std_logic_vector(37740, 16),
47565 => conv_std_logic_vector(37925, 16),
47566 => conv_std_logic_vector(38110, 16),
47567 => conv_std_logic_vector(38295, 16),
47568 => conv_std_logic_vector(38480, 16),
47569 => conv_std_logic_vector(38665, 16),
47570 => conv_std_logic_vector(38850, 16),
47571 => conv_std_logic_vector(39035, 16),
47572 => conv_std_logic_vector(39220, 16),
47573 => conv_std_logic_vector(39405, 16),
47574 => conv_std_logic_vector(39590, 16),
47575 => conv_std_logic_vector(39775, 16),
47576 => conv_std_logic_vector(39960, 16),
47577 => conv_std_logic_vector(40145, 16),
47578 => conv_std_logic_vector(40330, 16),
47579 => conv_std_logic_vector(40515, 16),
47580 => conv_std_logic_vector(40700, 16),
47581 => conv_std_logic_vector(40885, 16),
47582 => conv_std_logic_vector(41070, 16),
47583 => conv_std_logic_vector(41255, 16),
47584 => conv_std_logic_vector(41440, 16),
47585 => conv_std_logic_vector(41625, 16),
47586 => conv_std_logic_vector(41810, 16),
47587 => conv_std_logic_vector(41995, 16),
47588 => conv_std_logic_vector(42180, 16),
47589 => conv_std_logic_vector(42365, 16),
47590 => conv_std_logic_vector(42550, 16),
47591 => conv_std_logic_vector(42735, 16),
47592 => conv_std_logic_vector(42920, 16),
47593 => conv_std_logic_vector(43105, 16),
47594 => conv_std_logic_vector(43290, 16),
47595 => conv_std_logic_vector(43475, 16),
47596 => conv_std_logic_vector(43660, 16),
47597 => conv_std_logic_vector(43845, 16),
47598 => conv_std_logic_vector(44030, 16),
47599 => conv_std_logic_vector(44215, 16),
47600 => conv_std_logic_vector(44400, 16),
47601 => conv_std_logic_vector(44585, 16),
47602 => conv_std_logic_vector(44770, 16),
47603 => conv_std_logic_vector(44955, 16),
47604 => conv_std_logic_vector(45140, 16),
47605 => conv_std_logic_vector(45325, 16),
47606 => conv_std_logic_vector(45510, 16),
47607 => conv_std_logic_vector(45695, 16),
47608 => conv_std_logic_vector(45880, 16),
47609 => conv_std_logic_vector(46065, 16),
47610 => conv_std_logic_vector(46250, 16),
47611 => conv_std_logic_vector(46435, 16),
47612 => conv_std_logic_vector(46620, 16),
47613 => conv_std_logic_vector(46805, 16),
47614 => conv_std_logic_vector(46990, 16),
47615 => conv_std_logic_vector(47175, 16),
47616 => conv_std_logic_vector(0, 16),
47617 => conv_std_logic_vector(186, 16),
47618 => conv_std_logic_vector(372, 16),
47619 => conv_std_logic_vector(558, 16),
47620 => conv_std_logic_vector(744, 16),
47621 => conv_std_logic_vector(930, 16),
47622 => conv_std_logic_vector(1116, 16),
47623 => conv_std_logic_vector(1302, 16),
47624 => conv_std_logic_vector(1488, 16),
47625 => conv_std_logic_vector(1674, 16),
47626 => conv_std_logic_vector(1860, 16),
47627 => conv_std_logic_vector(2046, 16),
47628 => conv_std_logic_vector(2232, 16),
47629 => conv_std_logic_vector(2418, 16),
47630 => conv_std_logic_vector(2604, 16),
47631 => conv_std_logic_vector(2790, 16),
47632 => conv_std_logic_vector(2976, 16),
47633 => conv_std_logic_vector(3162, 16),
47634 => conv_std_logic_vector(3348, 16),
47635 => conv_std_logic_vector(3534, 16),
47636 => conv_std_logic_vector(3720, 16),
47637 => conv_std_logic_vector(3906, 16),
47638 => conv_std_logic_vector(4092, 16),
47639 => conv_std_logic_vector(4278, 16),
47640 => conv_std_logic_vector(4464, 16),
47641 => conv_std_logic_vector(4650, 16),
47642 => conv_std_logic_vector(4836, 16),
47643 => conv_std_logic_vector(5022, 16),
47644 => conv_std_logic_vector(5208, 16),
47645 => conv_std_logic_vector(5394, 16),
47646 => conv_std_logic_vector(5580, 16),
47647 => conv_std_logic_vector(5766, 16),
47648 => conv_std_logic_vector(5952, 16),
47649 => conv_std_logic_vector(6138, 16),
47650 => conv_std_logic_vector(6324, 16),
47651 => conv_std_logic_vector(6510, 16),
47652 => conv_std_logic_vector(6696, 16),
47653 => conv_std_logic_vector(6882, 16),
47654 => conv_std_logic_vector(7068, 16),
47655 => conv_std_logic_vector(7254, 16),
47656 => conv_std_logic_vector(7440, 16),
47657 => conv_std_logic_vector(7626, 16),
47658 => conv_std_logic_vector(7812, 16),
47659 => conv_std_logic_vector(7998, 16),
47660 => conv_std_logic_vector(8184, 16),
47661 => conv_std_logic_vector(8370, 16),
47662 => conv_std_logic_vector(8556, 16),
47663 => conv_std_logic_vector(8742, 16),
47664 => conv_std_logic_vector(8928, 16),
47665 => conv_std_logic_vector(9114, 16),
47666 => conv_std_logic_vector(9300, 16),
47667 => conv_std_logic_vector(9486, 16),
47668 => conv_std_logic_vector(9672, 16),
47669 => conv_std_logic_vector(9858, 16),
47670 => conv_std_logic_vector(10044, 16),
47671 => conv_std_logic_vector(10230, 16),
47672 => conv_std_logic_vector(10416, 16),
47673 => conv_std_logic_vector(10602, 16),
47674 => conv_std_logic_vector(10788, 16),
47675 => conv_std_logic_vector(10974, 16),
47676 => conv_std_logic_vector(11160, 16),
47677 => conv_std_logic_vector(11346, 16),
47678 => conv_std_logic_vector(11532, 16),
47679 => conv_std_logic_vector(11718, 16),
47680 => conv_std_logic_vector(11904, 16),
47681 => conv_std_logic_vector(12090, 16),
47682 => conv_std_logic_vector(12276, 16),
47683 => conv_std_logic_vector(12462, 16),
47684 => conv_std_logic_vector(12648, 16),
47685 => conv_std_logic_vector(12834, 16),
47686 => conv_std_logic_vector(13020, 16),
47687 => conv_std_logic_vector(13206, 16),
47688 => conv_std_logic_vector(13392, 16),
47689 => conv_std_logic_vector(13578, 16),
47690 => conv_std_logic_vector(13764, 16),
47691 => conv_std_logic_vector(13950, 16),
47692 => conv_std_logic_vector(14136, 16),
47693 => conv_std_logic_vector(14322, 16),
47694 => conv_std_logic_vector(14508, 16),
47695 => conv_std_logic_vector(14694, 16),
47696 => conv_std_logic_vector(14880, 16),
47697 => conv_std_logic_vector(15066, 16),
47698 => conv_std_logic_vector(15252, 16),
47699 => conv_std_logic_vector(15438, 16),
47700 => conv_std_logic_vector(15624, 16),
47701 => conv_std_logic_vector(15810, 16),
47702 => conv_std_logic_vector(15996, 16),
47703 => conv_std_logic_vector(16182, 16),
47704 => conv_std_logic_vector(16368, 16),
47705 => conv_std_logic_vector(16554, 16),
47706 => conv_std_logic_vector(16740, 16),
47707 => conv_std_logic_vector(16926, 16),
47708 => conv_std_logic_vector(17112, 16),
47709 => conv_std_logic_vector(17298, 16),
47710 => conv_std_logic_vector(17484, 16),
47711 => conv_std_logic_vector(17670, 16),
47712 => conv_std_logic_vector(17856, 16),
47713 => conv_std_logic_vector(18042, 16),
47714 => conv_std_logic_vector(18228, 16),
47715 => conv_std_logic_vector(18414, 16),
47716 => conv_std_logic_vector(18600, 16),
47717 => conv_std_logic_vector(18786, 16),
47718 => conv_std_logic_vector(18972, 16),
47719 => conv_std_logic_vector(19158, 16),
47720 => conv_std_logic_vector(19344, 16),
47721 => conv_std_logic_vector(19530, 16),
47722 => conv_std_logic_vector(19716, 16),
47723 => conv_std_logic_vector(19902, 16),
47724 => conv_std_logic_vector(20088, 16),
47725 => conv_std_logic_vector(20274, 16),
47726 => conv_std_logic_vector(20460, 16),
47727 => conv_std_logic_vector(20646, 16),
47728 => conv_std_logic_vector(20832, 16),
47729 => conv_std_logic_vector(21018, 16),
47730 => conv_std_logic_vector(21204, 16),
47731 => conv_std_logic_vector(21390, 16),
47732 => conv_std_logic_vector(21576, 16),
47733 => conv_std_logic_vector(21762, 16),
47734 => conv_std_logic_vector(21948, 16),
47735 => conv_std_logic_vector(22134, 16),
47736 => conv_std_logic_vector(22320, 16),
47737 => conv_std_logic_vector(22506, 16),
47738 => conv_std_logic_vector(22692, 16),
47739 => conv_std_logic_vector(22878, 16),
47740 => conv_std_logic_vector(23064, 16),
47741 => conv_std_logic_vector(23250, 16),
47742 => conv_std_logic_vector(23436, 16),
47743 => conv_std_logic_vector(23622, 16),
47744 => conv_std_logic_vector(23808, 16),
47745 => conv_std_logic_vector(23994, 16),
47746 => conv_std_logic_vector(24180, 16),
47747 => conv_std_logic_vector(24366, 16),
47748 => conv_std_logic_vector(24552, 16),
47749 => conv_std_logic_vector(24738, 16),
47750 => conv_std_logic_vector(24924, 16),
47751 => conv_std_logic_vector(25110, 16),
47752 => conv_std_logic_vector(25296, 16),
47753 => conv_std_logic_vector(25482, 16),
47754 => conv_std_logic_vector(25668, 16),
47755 => conv_std_logic_vector(25854, 16),
47756 => conv_std_logic_vector(26040, 16),
47757 => conv_std_logic_vector(26226, 16),
47758 => conv_std_logic_vector(26412, 16),
47759 => conv_std_logic_vector(26598, 16),
47760 => conv_std_logic_vector(26784, 16),
47761 => conv_std_logic_vector(26970, 16),
47762 => conv_std_logic_vector(27156, 16),
47763 => conv_std_logic_vector(27342, 16),
47764 => conv_std_logic_vector(27528, 16),
47765 => conv_std_logic_vector(27714, 16),
47766 => conv_std_logic_vector(27900, 16),
47767 => conv_std_logic_vector(28086, 16),
47768 => conv_std_logic_vector(28272, 16),
47769 => conv_std_logic_vector(28458, 16),
47770 => conv_std_logic_vector(28644, 16),
47771 => conv_std_logic_vector(28830, 16),
47772 => conv_std_logic_vector(29016, 16),
47773 => conv_std_logic_vector(29202, 16),
47774 => conv_std_logic_vector(29388, 16),
47775 => conv_std_logic_vector(29574, 16),
47776 => conv_std_logic_vector(29760, 16),
47777 => conv_std_logic_vector(29946, 16),
47778 => conv_std_logic_vector(30132, 16),
47779 => conv_std_logic_vector(30318, 16),
47780 => conv_std_logic_vector(30504, 16),
47781 => conv_std_logic_vector(30690, 16),
47782 => conv_std_logic_vector(30876, 16),
47783 => conv_std_logic_vector(31062, 16),
47784 => conv_std_logic_vector(31248, 16),
47785 => conv_std_logic_vector(31434, 16),
47786 => conv_std_logic_vector(31620, 16),
47787 => conv_std_logic_vector(31806, 16),
47788 => conv_std_logic_vector(31992, 16),
47789 => conv_std_logic_vector(32178, 16),
47790 => conv_std_logic_vector(32364, 16),
47791 => conv_std_logic_vector(32550, 16),
47792 => conv_std_logic_vector(32736, 16),
47793 => conv_std_logic_vector(32922, 16),
47794 => conv_std_logic_vector(33108, 16),
47795 => conv_std_logic_vector(33294, 16),
47796 => conv_std_logic_vector(33480, 16),
47797 => conv_std_logic_vector(33666, 16),
47798 => conv_std_logic_vector(33852, 16),
47799 => conv_std_logic_vector(34038, 16),
47800 => conv_std_logic_vector(34224, 16),
47801 => conv_std_logic_vector(34410, 16),
47802 => conv_std_logic_vector(34596, 16),
47803 => conv_std_logic_vector(34782, 16),
47804 => conv_std_logic_vector(34968, 16),
47805 => conv_std_logic_vector(35154, 16),
47806 => conv_std_logic_vector(35340, 16),
47807 => conv_std_logic_vector(35526, 16),
47808 => conv_std_logic_vector(35712, 16),
47809 => conv_std_logic_vector(35898, 16),
47810 => conv_std_logic_vector(36084, 16),
47811 => conv_std_logic_vector(36270, 16),
47812 => conv_std_logic_vector(36456, 16),
47813 => conv_std_logic_vector(36642, 16),
47814 => conv_std_logic_vector(36828, 16),
47815 => conv_std_logic_vector(37014, 16),
47816 => conv_std_logic_vector(37200, 16),
47817 => conv_std_logic_vector(37386, 16),
47818 => conv_std_logic_vector(37572, 16),
47819 => conv_std_logic_vector(37758, 16),
47820 => conv_std_logic_vector(37944, 16),
47821 => conv_std_logic_vector(38130, 16),
47822 => conv_std_logic_vector(38316, 16),
47823 => conv_std_logic_vector(38502, 16),
47824 => conv_std_logic_vector(38688, 16),
47825 => conv_std_logic_vector(38874, 16),
47826 => conv_std_logic_vector(39060, 16),
47827 => conv_std_logic_vector(39246, 16),
47828 => conv_std_logic_vector(39432, 16),
47829 => conv_std_logic_vector(39618, 16),
47830 => conv_std_logic_vector(39804, 16),
47831 => conv_std_logic_vector(39990, 16),
47832 => conv_std_logic_vector(40176, 16),
47833 => conv_std_logic_vector(40362, 16),
47834 => conv_std_logic_vector(40548, 16),
47835 => conv_std_logic_vector(40734, 16),
47836 => conv_std_logic_vector(40920, 16),
47837 => conv_std_logic_vector(41106, 16),
47838 => conv_std_logic_vector(41292, 16),
47839 => conv_std_logic_vector(41478, 16),
47840 => conv_std_logic_vector(41664, 16),
47841 => conv_std_logic_vector(41850, 16),
47842 => conv_std_logic_vector(42036, 16),
47843 => conv_std_logic_vector(42222, 16),
47844 => conv_std_logic_vector(42408, 16),
47845 => conv_std_logic_vector(42594, 16),
47846 => conv_std_logic_vector(42780, 16),
47847 => conv_std_logic_vector(42966, 16),
47848 => conv_std_logic_vector(43152, 16),
47849 => conv_std_logic_vector(43338, 16),
47850 => conv_std_logic_vector(43524, 16),
47851 => conv_std_logic_vector(43710, 16),
47852 => conv_std_logic_vector(43896, 16),
47853 => conv_std_logic_vector(44082, 16),
47854 => conv_std_logic_vector(44268, 16),
47855 => conv_std_logic_vector(44454, 16),
47856 => conv_std_logic_vector(44640, 16),
47857 => conv_std_logic_vector(44826, 16),
47858 => conv_std_logic_vector(45012, 16),
47859 => conv_std_logic_vector(45198, 16),
47860 => conv_std_logic_vector(45384, 16),
47861 => conv_std_logic_vector(45570, 16),
47862 => conv_std_logic_vector(45756, 16),
47863 => conv_std_logic_vector(45942, 16),
47864 => conv_std_logic_vector(46128, 16),
47865 => conv_std_logic_vector(46314, 16),
47866 => conv_std_logic_vector(46500, 16),
47867 => conv_std_logic_vector(46686, 16),
47868 => conv_std_logic_vector(46872, 16),
47869 => conv_std_logic_vector(47058, 16),
47870 => conv_std_logic_vector(47244, 16),
47871 => conv_std_logic_vector(47430, 16),
47872 => conv_std_logic_vector(0, 16),
47873 => conv_std_logic_vector(187, 16),
47874 => conv_std_logic_vector(374, 16),
47875 => conv_std_logic_vector(561, 16),
47876 => conv_std_logic_vector(748, 16),
47877 => conv_std_logic_vector(935, 16),
47878 => conv_std_logic_vector(1122, 16),
47879 => conv_std_logic_vector(1309, 16),
47880 => conv_std_logic_vector(1496, 16),
47881 => conv_std_logic_vector(1683, 16),
47882 => conv_std_logic_vector(1870, 16),
47883 => conv_std_logic_vector(2057, 16),
47884 => conv_std_logic_vector(2244, 16),
47885 => conv_std_logic_vector(2431, 16),
47886 => conv_std_logic_vector(2618, 16),
47887 => conv_std_logic_vector(2805, 16),
47888 => conv_std_logic_vector(2992, 16),
47889 => conv_std_logic_vector(3179, 16),
47890 => conv_std_logic_vector(3366, 16),
47891 => conv_std_logic_vector(3553, 16),
47892 => conv_std_logic_vector(3740, 16),
47893 => conv_std_logic_vector(3927, 16),
47894 => conv_std_logic_vector(4114, 16),
47895 => conv_std_logic_vector(4301, 16),
47896 => conv_std_logic_vector(4488, 16),
47897 => conv_std_logic_vector(4675, 16),
47898 => conv_std_logic_vector(4862, 16),
47899 => conv_std_logic_vector(5049, 16),
47900 => conv_std_logic_vector(5236, 16),
47901 => conv_std_logic_vector(5423, 16),
47902 => conv_std_logic_vector(5610, 16),
47903 => conv_std_logic_vector(5797, 16),
47904 => conv_std_logic_vector(5984, 16),
47905 => conv_std_logic_vector(6171, 16),
47906 => conv_std_logic_vector(6358, 16),
47907 => conv_std_logic_vector(6545, 16),
47908 => conv_std_logic_vector(6732, 16),
47909 => conv_std_logic_vector(6919, 16),
47910 => conv_std_logic_vector(7106, 16),
47911 => conv_std_logic_vector(7293, 16),
47912 => conv_std_logic_vector(7480, 16),
47913 => conv_std_logic_vector(7667, 16),
47914 => conv_std_logic_vector(7854, 16),
47915 => conv_std_logic_vector(8041, 16),
47916 => conv_std_logic_vector(8228, 16),
47917 => conv_std_logic_vector(8415, 16),
47918 => conv_std_logic_vector(8602, 16),
47919 => conv_std_logic_vector(8789, 16),
47920 => conv_std_logic_vector(8976, 16),
47921 => conv_std_logic_vector(9163, 16),
47922 => conv_std_logic_vector(9350, 16),
47923 => conv_std_logic_vector(9537, 16),
47924 => conv_std_logic_vector(9724, 16),
47925 => conv_std_logic_vector(9911, 16),
47926 => conv_std_logic_vector(10098, 16),
47927 => conv_std_logic_vector(10285, 16),
47928 => conv_std_logic_vector(10472, 16),
47929 => conv_std_logic_vector(10659, 16),
47930 => conv_std_logic_vector(10846, 16),
47931 => conv_std_logic_vector(11033, 16),
47932 => conv_std_logic_vector(11220, 16),
47933 => conv_std_logic_vector(11407, 16),
47934 => conv_std_logic_vector(11594, 16),
47935 => conv_std_logic_vector(11781, 16),
47936 => conv_std_logic_vector(11968, 16),
47937 => conv_std_logic_vector(12155, 16),
47938 => conv_std_logic_vector(12342, 16),
47939 => conv_std_logic_vector(12529, 16),
47940 => conv_std_logic_vector(12716, 16),
47941 => conv_std_logic_vector(12903, 16),
47942 => conv_std_logic_vector(13090, 16),
47943 => conv_std_logic_vector(13277, 16),
47944 => conv_std_logic_vector(13464, 16),
47945 => conv_std_logic_vector(13651, 16),
47946 => conv_std_logic_vector(13838, 16),
47947 => conv_std_logic_vector(14025, 16),
47948 => conv_std_logic_vector(14212, 16),
47949 => conv_std_logic_vector(14399, 16),
47950 => conv_std_logic_vector(14586, 16),
47951 => conv_std_logic_vector(14773, 16),
47952 => conv_std_logic_vector(14960, 16),
47953 => conv_std_logic_vector(15147, 16),
47954 => conv_std_logic_vector(15334, 16),
47955 => conv_std_logic_vector(15521, 16),
47956 => conv_std_logic_vector(15708, 16),
47957 => conv_std_logic_vector(15895, 16),
47958 => conv_std_logic_vector(16082, 16),
47959 => conv_std_logic_vector(16269, 16),
47960 => conv_std_logic_vector(16456, 16),
47961 => conv_std_logic_vector(16643, 16),
47962 => conv_std_logic_vector(16830, 16),
47963 => conv_std_logic_vector(17017, 16),
47964 => conv_std_logic_vector(17204, 16),
47965 => conv_std_logic_vector(17391, 16),
47966 => conv_std_logic_vector(17578, 16),
47967 => conv_std_logic_vector(17765, 16),
47968 => conv_std_logic_vector(17952, 16),
47969 => conv_std_logic_vector(18139, 16),
47970 => conv_std_logic_vector(18326, 16),
47971 => conv_std_logic_vector(18513, 16),
47972 => conv_std_logic_vector(18700, 16),
47973 => conv_std_logic_vector(18887, 16),
47974 => conv_std_logic_vector(19074, 16),
47975 => conv_std_logic_vector(19261, 16),
47976 => conv_std_logic_vector(19448, 16),
47977 => conv_std_logic_vector(19635, 16),
47978 => conv_std_logic_vector(19822, 16),
47979 => conv_std_logic_vector(20009, 16),
47980 => conv_std_logic_vector(20196, 16),
47981 => conv_std_logic_vector(20383, 16),
47982 => conv_std_logic_vector(20570, 16),
47983 => conv_std_logic_vector(20757, 16),
47984 => conv_std_logic_vector(20944, 16),
47985 => conv_std_logic_vector(21131, 16),
47986 => conv_std_logic_vector(21318, 16),
47987 => conv_std_logic_vector(21505, 16),
47988 => conv_std_logic_vector(21692, 16),
47989 => conv_std_logic_vector(21879, 16),
47990 => conv_std_logic_vector(22066, 16),
47991 => conv_std_logic_vector(22253, 16),
47992 => conv_std_logic_vector(22440, 16),
47993 => conv_std_logic_vector(22627, 16),
47994 => conv_std_logic_vector(22814, 16),
47995 => conv_std_logic_vector(23001, 16),
47996 => conv_std_logic_vector(23188, 16),
47997 => conv_std_logic_vector(23375, 16),
47998 => conv_std_logic_vector(23562, 16),
47999 => conv_std_logic_vector(23749, 16),
48000 => conv_std_logic_vector(23936, 16),
48001 => conv_std_logic_vector(24123, 16),
48002 => conv_std_logic_vector(24310, 16),
48003 => conv_std_logic_vector(24497, 16),
48004 => conv_std_logic_vector(24684, 16),
48005 => conv_std_logic_vector(24871, 16),
48006 => conv_std_logic_vector(25058, 16),
48007 => conv_std_logic_vector(25245, 16),
48008 => conv_std_logic_vector(25432, 16),
48009 => conv_std_logic_vector(25619, 16),
48010 => conv_std_logic_vector(25806, 16),
48011 => conv_std_logic_vector(25993, 16),
48012 => conv_std_logic_vector(26180, 16),
48013 => conv_std_logic_vector(26367, 16),
48014 => conv_std_logic_vector(26554, 16),
48015 => conv_std_logic_vector(26741, 16),
48016 => conv_std_logic_vector(26928, 16),
48017 => conv_std_logic_vector(27115, 16),
48018 => conv_std_logic_vector(27302, 16),
48019 => conv_std_logic_vector(27489, 16),
48020 => conv_std_logic_vector(27676, 16),
48021 => conv_std_logic_vector(27863, 16),
48022 => conv_std_logic_vector(28050, 16),
48023 => conv_std_logic_vector(28237, 16),
48024 => conv_std_logic_vector(28424, 16),
48025 => conv_std_logic_vector(28611, 16),
48026 => conv_std_logic_vector(28798, 16),
48027 => conv_std_logic_vector(28985, 16),
48028 => conv_std_logic_vector(29172, 16),
48029 => conv_std_logic_vector(29359, 16),
48030 => conv_std_logic_vector(29546, 16),
48031 => conv_std_logic_vector(29733, 16),
48032 => conv_std_logic_vector(29920, 16),
48033 => conv_std_logic_vector(30107, 16),
48034 => conv_std_logic_vector(30294, 16),
48035 => conv_std_logic_vector(30481, 16),
48036 => conv_std_logic_vector(30668, 16),
48037 => conv_std_logic_vector(30855, 16),
48038 => conv_std_logic_vector(31042, 16),
48039 => conv_std_logic_vector(31229, 16),
48040 => conv_std_logic_vector(31416, 16),
48041 => conv_std_logic_vector(31603, 16),
48042 => conv_std_logic_vector(31790, 16),
48043 => conv_std_logic_vector(31977, 16),
48044 => conv_std_logic_vector(32164, 16),
48045 => conv_std_logic_vector(32351, 16),
48046 => conv_std_logic_vector(32538, 16),
48047 => conv_std_logic_vector(32725, 16),
48048 => conv_std_logic_vector(32912, 16),
48049 => conv_std_logic_vector(33099, 16),
48050 => conv_std_logic_vector(33286, 16),
48051 => conv_std_logic_vector(33473, 16),
48052 => conv_std_logic_vector(33660, 16),
48053 => conv_std_logic_vector(33847, 16),
48054 => conv_std_logic_vector(34034, 16),
48055 => conv_std_logic_vector(34221, 16),
48056 => conv_std_logic_vector(34408, 16),
48057 => conv_std_logic_vector(34595, 16),
48058 => conv_std_logic_vector(34782, 16),
48059 => conv_std_logic_vector(34969, 16),
48060 => conv_std_logic_vector(35156, 16),
48061 => conv_std_logic_vector(35343, 16),
48062 => conv_std_logic_vector(35530, 16),
48063 => conv_std_logic_vector(35717, 16),
48064 => conv_std_logic_vector(35904, 16),
48065 => conv_std_logic_vector(36091, 16),
48066 => conv_std_logic_vector(36278, 16),
48067 => conv_std_logic_vector(36465, 16),
48068 => conv_std_logic_vector(36652, 16),
48069 => conv_std_logic_vector(36839, 16),
48070 => conv_std_logic_vector(37026, 16),
48071 => conv_std_logic_vector(37213, 16),
48072 => conv_std_logic_vector(37400, 16),
48073 => conv_std_logic_vector(37587, 16),
48074 => conv_std_logic_vector(37774, 16),
48075 => conv_std_logic_vector(37961, 16),
48076 => conv_std_logic_vector(38148, 16),
48077 => conv_std_logic_vector(38335, 16),
48078 => conv_std_logic_vector(38522, 16),
48079 => conv_std_logic_vector(38709, 16),
48080 => conv_std_logic_vector(38896, 16),
48081 => conv_std_logic_vector(39083, 16),
48082 => conv_std_logic_vector(39270, 16),
48083 => conv_std_logic_vector(39457, 16),
48084 => conv_std_logic_vector(39644, 16),
48085 => conv_std_logic_vector(39831, 16),
48086 => conv_std_logic_vector(40018, 16),
48087 => conv_std_logic_vector(40205, 16),
48088 => conv_std_logic_vector(40392, 16),
48089 => conv_std_logic_vector(40579, 16),
48090 => conv_std_logic_vector(40766, 16),
48091 => conv_std_logic_vector(40953, 16),
48092 => conv_std_logic_vector(41140, 16),
48093 => conv_std_logic_vector(41327, 16),
48094 => conv_std_logic_vector(41514, 16),
48095 => conv_std_logic_vector(41701, 16),
48096 => conv_std_logic_vector(41888, 16),
48097 => conv_std_logic_vector(42075, 16),
48098 => conv_std_logic_vector(42262, 16),
48099 => conv_std_logic_vector(42449, 16),
48100 => conv_std_logic_vector(42636, 16),
48101 => conv_std_logic_vector(42823, 16),
48102 => conv_std_logic_vector(43010, 16),
48103 => conv_std_logic_vector(43197, 16),
48104 => conv_std_logic_vector(43384, 16),
48105 => conv_std_logic_vector(43571, 16),
48106 => conv_std_logic_vector(43758, 16),
48107 => conv_std_logic_vector(43945, 16),
48108 => conv_std_logic_vector(44132, 16),
48109 => conv_std_logic_vector(44319, 16),
48110 => conv_std_logic_vector(44506, 16),
48111 => conv_std_logic_vector(44693, 16),
48112 => conv_std_logic_vector(44880, 16),
48113 => conv_std_logic_vector(45067, 16),
48114 => conv_std_logic_vector(45254, 16),
48115 => conv_std_logic_vector(45441, 16),
48116 => conv_std_logic_vector(45628, 16),
48117 => conv_std_logic_vector(45815, 16),
48118 => conv_std_logic_vector(46002, 16),
48119 => conv_std_logic_vector(46189, 16),
48120 => conv_std_logic_vector(46376, 16),
48121 => conv_std_logic_vector(46563, 16),
48122 => conv_std_logic_vector(46750, 16),
48123 => conv_std_logic_vector(46937, 16),
48124 => conv_std_logic_vector(47124, 16),
48125 => conv_std_logic_vector(47311, 16),
48126 => conv_std_logic_vector(47498, 16),
48127 => conv_std_logic_vector(47685, 16),
48128 => conv_std_logic_vector(0, 16),
48129 => conv_std_logic_vector(188, 16),
48130 => conv_std_logic_vector(376, 16),
48131 => conv_std_logic_vector(564, 16),
48132 => conv_std_logic_vector(752, 16),
48133 => conv_std_logic_vector(940, 16),
48134 => conv_std_logic_vector(1128, 16),
48135 => conv_std_logic_vector(1316, 16),
48136 => conv_std_logic_vector(1504, 16),
48137 => conv_std_logic_vector(1692, 16),
48138 => conv_std_logic_vector(1880, 16),
48139 => conv_std_logic_vector(2068, 16),
48140 => conv_std_logic_vector(2256, 16),
48141 => conv_std_logic_vector(2444, 16),
48142 => conv_std_logic_vector(2632, 16),
48143 => conv_std_logic_vector(2820, 16),
48144 => conv_std_logic_vector(3008, 16),
48145 => conv_std_logic_vector(3196, 16),
48146 => conv_std_logic_vector(3384, 16),
48147 => conv_std_logic_vector(3572, 16),
48148 => conv_std_logic_vector(3760, 16),
48149 => conv_std_logic_vector(3948, 16),
48150 => conv_std_logic_vector(4136, 16),
48151 => conv_std_logic_vector(4324, 16),
48152 => conv_std_logic_vector(4512, 16),
48153 => conv_std_logic_vector(4700, 16),
48154 => conv_std_logic_vector(4888, 16),
48155 => conv_std_logic_vector(5076, 16),
48156 => conv_std_logic_vector(5264, 16),
48157 => conv_std_logic_vector(5452, 16),
48158 => conv_std_logic_vector(5640, 16),
48159 => conv_std_logic_vector(5828, 16),
48160 => conv_std_logic_vector(6016, 16),
48161 => conv_std_logic_vector(6204, 16),
48162 => conv_std_logic_vector(6392, 16),
48163 => conv_std_logic_vector(6580, 16),
48164 => conv_std_logic_vector(6768, 16),
48165 => conv_std_logic_vector(6956, 16),
48166 => conv_std_logic_vector(7144, 16),
48167 => conv_std_logic_vector(7332, 16),
48168 => conv_std_logic_vector(7520, 16),
48169 => conv_std_logic_vector(7708, 16),
48170 => conv_std_logic_vector(7896, 16),
48171 => conv_std_logic_vector(8084, 16),
48172 => conv_std_logic_vector(8272, 16),
48173 => conv_std_logic_vector(8460, 16),
48174 => conv_std_logic_vector(8648, 16),
48175 => conv_std_logic_vector(8836, 16),
48176 => conv_std_logic_vector(9024, 16),
48177 => conv_std_logic_vector(9212, 16),
48178 => conv_std_logic_vector(9400, 16),
48179 => conv_std_logic_vector(9588, 16),
48180 => conv_std_logic_vector(9776, 16),
48181 => conv_std_logic_vector(9964, 16),
48182 => conv_std_logic_vector(10152, 16),
48183 => conv_std_logic_vector(10340, 16),
48184 => conv_std_logic_vector(10528, 16),
48185 => conv_std_logic_vector(10716, 16),
48186 => conv_std_logic_vector(10904, 16),
48187 => conv_std_logic_vector(11092, 16),
48188 => conv_std_logic_vector(11280, 16),
48189 => conv_std_logic_vector(11468, 16),
48190 => conv_std_logic_vector(11656, 16),
48191 => conv_std_logic_vector(11844, 16),
48192 => conv_std_logic_vector(12032, 16),
48193 => conv_std_logic_vector(12220, 16),
48194 => conv_std_logic_vector(12408, 16),
48195 => conv_std_logic_vector(12596, 16),
48196 => conv_std_logic_vector(12784, 16),
48197 => conv_std_logic_vector(12972, 16),
48198 => conv_std_logic_vector(13160, 16),
48199 => conv_std_logic_vector(13348, 16),
48200 => conv_std_logic_vector(13536, 16),
48201 => conv_std_logic_vector(13724, 16),
48202 => conv_std_logic_vector(13912, 16),
48203 => conv_std_logic_vector(14100, 16),
48204 => conv_std_logic_vector(14288, 16),
48205 => conv_std_logic_vector(14476, 16),
48206 => conv_std_logic_vector(14664, 16),
48207 => conv_std_logic_vector(14852, 16),
48208 => conv_std_logic_vector(15040, 16),
48209 => conv_std_logic_vector(15228, 16),
48210 => conv_std_logic_vector(15416, 16),
48211 => conv_std_logic_vector(15604, 16),
48212 => conv_std_logic_vector(15792, 16),
48213 => conv_std_logic_vector(15980, 16),
48214 => conv_std_logic_vector(16168, 16),
48215 => conv_std_logic_vector(16356, 16),
48216 => conv_std_logic_vector(16544, 16),
48217 => conv_std_logic_vector(16732, 16),
48218 => conv_std_logic_vector(16920, 16),
48219 => conv_std_logic_vector(17108, 16),
48220 => conv_std_logic_vector(17296, 16),
48221 => conv_std_logic_vector(17484, 16),
48222 => conv_std_logic_vector(17672, 16),
48223 => conv_std_logic_vector(17860, 16),
48224 => conv_std_logic_vector(18048, 16),
48225 => conv_std_logic_vector(18236, 16),
48226 => conv_std_logic_vector(18424, 16),
48227 => conv_std_logic_vector(18612, 16),
48228 => conv_std_logic_vector(18800, 16),
48229 => conv_std_logic_vector(18988, 16),
48230 => conv_std_logic_vector(19176, 16),
48231 => conv_std_logic_vector(19364, 16),
48232 => conv_std_logic_vector(19552, 16),
48233 => conv_std_logic_vector(19740, 16),
48234 => conv_std_logic_vector(19928, 16),
48235 => conv_std_logic_vector(20116, 16),
48236 => conv_std_logic_vector(20304, 16),
48237 => conv_std_logic_vector(20492, 16),
48238 => conv_std_logic_vector(20680, 16),
48239 => conv_std_logic_vector(20868, 16),
48240 => conv_std_logic_vector(21056, 16),
48241 => conv_std_logic_vector(21244, 16),
48242 => conv_std_logic_vector(21432, 16),
48243 => conv_std_logic_vector(21620, 16),
48244 => conv_std_logic_vector(21808, 16),
48245 => conv_std_logic_vector(21996, 16),
48246 => conv_std_logic_vector(22184, 16),
48247 => conv_std_logic_vector(22372, 16),
48248 => conv_std_logic_vector(22560, 16),
48249 => conv_std_logic_vector(22748, 16),
48250 => conv_std_logic_vector(22936, 16),
48251 => conv_std_logic_vector(23124, 16),
48252 => conv_std_logic_vector(23312, 16),
48253 => conv_std_logic_vector(23500, 16),
48254 => conv_std_logic_vector(23688, 16),
48255 => conv_std_logic_vector(23876, 16),
48256 => conv_std_logic_vector(24064, 16),
48257 => conv_std_logic_vector(24252, 16),
48258 => conv_std_logic_vector(24440, 16),
48259 => conv_std_logic_vector(24628, 16),
48260 => conv_std_logic_vector(24816, 16),
48261 => conv_std_logic_vector(25004, 16),
48262 => conv_std_logic_vector(25192, 16),
48263 => conv_std_logic_vector(25380, 16),
48264 => conv_std_logic_vector(25568, 16),
48265 => conv_std_logic_vector(25756, 16),
48266 => conv_std_logic_vector(25944, 16),
48267 => conv_std_logic_vector(26132, 16),
48268 => conv_std_logic_vector(26320, 16),
48269 => conv_std_logic_vector(26508, 16),
48270 => conv_std_logic_vector(26696, 16),
48271 => conv_std_logic_vector(26884, 16),
48272 => conv_std_logic_vector(27072, 16),
48273 => conv_std_logic_vector(27260, 16),
48274 => conv_std_logic_vector(27448, 16),
48275 => conv_std_logic_vector(27636, 16),
48276 => conv_std_logic_vector(27824, 16),
48277 => conv_std_logic_vector(28012, 16),
48278 => conv_std_logic_vector(28200, 16),
48279 => conv_std_logic_vector(28388, 16),
48280 => conv_std_logic_vector(28576, 16),
48281 => conv_std_logic_vector(28764, 16),
48282 => conv_std_logic_vector(28952, 16),
48283 => conv_std_logic_vector(29140, 16),
48284 => conv_std_logic_vector(29328, 16),
48285 => conv_std_logic_vector(29516, 16),
48286 => conv_std_logic_vector(29704, 16),
48287 => conv_std_logic_vector(29892, 16),
48288 => conv_std_logic_vector(30080, 16),
48289 => conv_std_logic_vector(30268, 16),
48290 => conv_std_logic_vector(30456, 16),
48291 => conv_std_logic_vector(30644, 16),
48292 => conv_std_logic_vector(30832, 16),
48293 => conv_std_logic_vector(31020, 16),
48294 => conv_std_logic_vector(31208, 16),
48295 => conv_std_logic_vector(31396, 16),
48296 => conv_std_logic_vector(31584, 16),
48297 => conv_std_logic_vector(31772, 16),
48298 => conv_std_logic_vector(31960, 16),
48299 => conv_std_logic_vector(32148, 16),
48300 => conv_std_logic_vector(32336, 16),
48301 => conv_std_logic_vector(32524, 16),
48302 => conv_std_logic_vector(32712, 16),
48303 => conv_std_logic_vector(32900, 16),
48304 => conv_std_logic_vector(33088, 16),
48305 => conv_std_logic_vector(33276, 16),
48306 => conv_std_logic_vector(33464, 16),
48307 => conv_std_logic_vector(33652, 16),
48308 => conv_std_logic_vector(33840, 16),
48309 => conv_std_logic_vector(34028, 16),
48310 => conv_std_logic_vector(34216, 16),
48311 => conv_std_logic_vector(34404, 16),
48312 => conv_std_logic_vector(34592, 16),
48313 => conv_std_logic_vector(34780, 16),
48314 => conv_std_logic_vector(34968, 16),
48315 => conv_std_logic_vector(35156, 16),
48316 => conv_std_logic_vector(35344, 16),
48317 => conv_std_logic_vector(35532, 16),
48318 => conv_std_logic_vector(35720, 16),
48319 => conv_std_logic_vector(35908, 16),
48320 => conv_std_logic_vector(36096, 16),
48321 => conv_std_logic_vector(36284, 16),
48322 => conv_std_logic_vector(36472, 16),
48323 => conv_std_logic_vector(36660, 16),
48324 => conv_std_logic_vector(36848, 16),
48325 => conv_std_logic_vector(37036, 16),
48326 => conv_std_logic_vector(37224, 16),
48327 => conv_std_logic_vector(37412, 16),
48328 => conv_std_logic_vector(37600, 16),
48329 => conv_std_logic_vector(37788, 16),
48330 => conv_std_logic_vector(37976, 16),
48331 => conv_std_logic_vector(38164, 16),
48332 => conv_std_logic_vector(38352, 16),
48333 => conv_std_logic_vector(38540, 16),
48334 => conv_std_logic_vector(38728, 16),
48335 => conv_std_logic_vector(38916, 16),
48336 => conv_std_logic_vector(39104, 16),
48337 => conv_std_logic_vector(39292, 16),
48338 => conv_std_logic_vector(39480, 16),
48339 => conv_std_logic_vector(39668, 16),
48340 => conv_std_logic_vector(39856, 16),
48341 => conv_std_logic_vector(40044, 16),
48342 => conv_std_logic_vector(40232, 16),
48343 => conv_std_logic_vector(40420, 16),
48344 => conv_std_logic_vector(40608, 16),
48345 => conv_std_logic_vector(40796, 16),
48346 => conv_std_logic_vector(40984, 16),
48347 => conv_std_logic_vector(41172, 16),
48348 => conv_std_logic_vector(41360, 16),
48349 => conv_std_logic_vector(41548, 16),
48350 => conv_std_logic_vector(41736, 16),
48351 => conv_std_logic_vector(41924, 16),
48352 => conv_std_logic_vector(42112, 16),
48353 => conv_std_logic_vector(42300, 16),
48354 => conv_std_logic_vector(42488, 16),
48355 => conv_std_logic_vector(42676, 16),
48356 => conv_std_logic_vector(42864, 16),
48357 => conv_std_logic_vector(43052, 16),
48358 => conv_std_logic_vector(43240, 16),
48359 => conv_std_logic_vector(43428, 16),
48360 => conv_std_logic_vector(43616, 16),
48361 => conv_std_logic_vector(43804, 16),
48362 => conv_std_logic_vector(43992, 16),
48363 => conv_std_logic_vector(44180, 16),
48364 => conv_std_logic_vector(44368, 16),
48365 => conv_std_logic_vector(44556, 16),
48366 => conv_std_logic_vector(44744, 16),
48367 => conv_std_logic_vector(44932, 16),
48368 => conv_std_logic_vector(45120, 16),
48369 => conv_std_logic_vector(45308, 16),
48370 => conv_std_logic_vector(45496, 16),
48371 => conv_std_logic_vector(45684, 16),
48372 => conv_std_logic_vector(45872, 16),
48373 => conv_std_logic_vector(46060, 16),
48374 => conv_std_logic_vector(46248, 16),
48375 => conv_std_logic_vector(46436, 16),
48376 => conv_std_logic_vector(46624, 16),
48377 => conv_std_logic_vector(46812, 16),
48378 => conv_std_logic_vector(47000, 16),
48379 => conv_std_logic_vector(47188, 16),
48380 => conv_std_logic_vector(47376, 16),
48381 => conv_std_logic_vector(47564, 16),
48382 => conv_std_logic_vector(47752, 16),
48383 => conv_std_logic_vector(47940, 16),
48384 => conv_std_logic_vector(0, 16),
48385 => conv_std_logic_vector(189, 16),
48386 => conv_std_logic_vector(378, 16),
48387 => conv_std_logic_vector(567, 16),
48388 => conv_std_logic_vector(756, 16),
48389 => conv_std_logic_vector(945, 16),
48390 => conv_std_logic_vector(1134, 16),
48391 => conv_std_logic_vector(1323, 16),
48392 => conv_std_logic_vector(1512, 16),
48393 => conv_std_logic_vector(1701, 16),
48394 => conv_std_logic_vector(1890, 16),
48395 => conv_std_logic_vector(2079, 16),
48396 => conv_std_logic_vector(2268, 16),
48397 => conv_std_logic_vector(2457, 16),
48398 => conv_std_logic_vector(2646, 16),
48399 => conv_std_logic_vector(2835, 16),
48400 => conv_std_logic_vector(3024, 16),
48401 => conv_std_logic_vector(3213, 16),
48402 => conv_std_logic_vector(3402, 16),
48403 => conv_std_logic_vector(3591, 16),
48404 => conv_std_logic_vector(3780, 16),
48405 => conv_std_logic_vector(3969, 16),
48406 => conv_std_logic_vector(4158, 16),
48407 => conv_std_logic_vector(4347, 16),
48408 => conv_std_logic_vector(4536, 16),
48409 => conv_std_logic_vector(4725, 16),
48410 => conv_std_logic_vector(4914, 16),
48411 => conv_std_logic_vector(5103, 16),
48412 => conv_std_logic_vector(5292, 16),
48413 => conv_std_logic_vector(5481, 16),
48414 => conv_std_logic_vector(5670, 16),
48415 => conv_std_logic_vector(5859, 16),
48416 => conv_std_logic_vector(6048, 16),
48417 => conv_std_logic_vector(6237, 16),
48418 => conv_std_logic_vector(6426, 16),
48419 => conv_std_logic_vector(6615, 16),
48420 => conv_std_logic_vector(6804, 16),
48421 => conv_std_logic_vector(6993, 16),
48422 => conv_std_logic_vector(7182, 16),
48423 => conv_std_logic_vector(7371, 16),
48424 => conv_std_logic_vector(7560, 16),
48425 => conv_std_logic_vector(7749, 16),
48426 => conv_std_logic_vector(7938, 16),
48427 => conv_std_logic_vector(8127, 16),
48428 => conv_std_logic_vector(8316, 16),
48429 => conv_std_logic_vector(8505, 16),
48430 => conv_std_logic_vector(8694, 16),
48431 => conv_std_logic_vector(8883, 16),
48432 => conv_std_logic_vector(9072, 16),
48433 => conv_std_logic_vector(9261, 16),
48434 => conv_std_logic_vector(9450, 16),
48435 => conv_std_logic_vector(9639, 16),
48436 => conv_std_logic_vector(9828, 16),
48437 => conv_std_logic_vector(10017, 16),
48438 => conv_std_logic_vector(10206, 16),
48439 => conv_std_logic_vector(10395, 16),
48440 => conv_std_logic_vector(10584, 16),
48441 => conv_std_logic_vector(10773, 16),
48442 => conv_std_logic_vector(10962, 16),
48443 => conv_std_logic_vector(11151, 16),
48444 => conv_std_logic_vector(11340, 16),
48445 => conv_std_logic_vector(11529, 16),
48446 => conv_std_logic_vector(11718, 16),
48447 => conv_std_logic_vector(11907, 16),
48448 => conv_std_logic_vector(12096, 16),
48449 => conv_std_logic_vector(12285, 16),
48450 => conv_std_logic_vector(12474, 16),
48451 => conv_std_logic_vector(12663, 16),
48452 => conv_std_logic_vector(12852, 16),
48453 => conv_std_logic_vector(13041, 16),
48454 => conv_std_logic_vector(13230, 16),
48455 => conv_std_logic_vector(13419, 16),
48456 => conv_std_logic_vector(13608, 16),
48457 => conv_std_logic_vector(13797, 16),
48458 => conv_std_logic_vector(13986, 16),
48459 => conv_std_logic_vector(14175, 16),
48460 => conv_std_logic_vector(14364, 16),
48461 => conv_std_logic_vector(14553, 16),
48462 => conv_std_logic_vector(14742, 16),
48463 => conv_std_logic_vector(14931, 16),
48464 => conv_std_logic_vector(15120, 16),
48465 => conv_std_logic_vector(15309, 16),
48466 => conv_std_logic_vector(15498, 16),
48467 => conv_std_logic_vector(15687, 16),
48468 => conv_std_logic_vector(15876, 16),
48469 => conv_std_logic_vector(16065, 16),
48470 => conv_std_logic_vector(16254, 16),
48471 => conv_std_logic_vector(16443, 16),
48472 => conv_std_logic_vector(16632, 16),
48473 => conv_std_logic_vector(16821, 16),
48474 => conv_std_logic_vector(17010, 16),
48475 => conv_std_logic_vector(17199, 16),
48476 => conv_std_logic_vector(17388, 16),
48477 => conv_std_logic_vector(17577, 16),
48478 => conv_std_logic_vector(17766, 16),
48479 => conv_std_logic_vector(17955, 16),
48480 => conv_std_logic_vector(18144, 16),
48481 => conv_std_logic_vector(18333, 16),
48482 => conv_std_logic_vector(18522, 16),
48483 => conv_std_logic_vector(18711, 16),
48484 => conv_std_logic_vector(18900, 16),
48485 => conv_std_logic_vector(19089, 16),
48486 => conv_std_logic_vector(19278, 16),
48487 => conv_std_logic_vector(19467, 16),
48488 => conv_std_logic_vector(19656, 16),
48489 => conv_std_logic_vector(19845, 16),
48490 => conv_std_logic_vector(20034, 16),
48491 => conv_std_logic_vector(20223, 16),
48492 => conv_std_logic_vector(20412, 16),
48493 => conv_std_logic_vector(20601, 16),
48494 => conv_std_logic_vector(20790, 16),
48495 => conv_std_logic_vector(20979, 16),
48496 => conv_std_logic_vector(21168, 16),
48497 => conv_std_logic_vector(21357, 16),
48498 => conv_std_logic_vector(21546, 16),
48499 => conv_std_logic_vector(21735, 16),
48500 => conv_std_logic_vector(21924, 16),
48501 => conv_std_logic_vector(22113, 16),
48502 => conv_std_logic_vector(22302, 16),
48503 => conv_std_logic_vector(22491, 16),
48504 => conv_std_logic_vector(22680, 16),
48505 => conv_std_logic_vector(22869, 16),
48506 => conv_std_logic_vector(23058, 16),
48507 => conv_std_logic_vector(23247, 16),
48508 => conv_std_logic_vector(23436, 16),
48509 => conv_std_logic_vector(23625, 16),
48510 => conv_std_logic_vector(23814, 16),
48511 => conv_std_logic_vector(24003, 16),
48512 => conv_std_logic_vector(24192, 16),
48513 => conv_std_logic_vector(24381, 16),
48514 => conv_std_logic_vector(24570, 16),
48515 => conv_std_logic_vector(24759, 16),
48516 => conv_std_logic_vector(24948, 16),
48517 => conv_std_logic_vector(25137, 16),
48518 => conv_std_logic_vector(25326, 16),
48519 => conv_std_logic_vector(25515, 16),
48520 => conv_std_logic_vector(25704, 16),
48521 => conv_std_logic_vector(25893, 16),
48522 => conv_std_logic_vector(26082, 16),
48523 => conv_std_logic_vector(26271, 16),
48524 => conv_std_logic_vector(26460, 16),
48525 => conv_std_logic_vector(26649, 16),
48526 => conv_std_logic_vector(26838, 16),
48527 => conv_std_logic_vector(27027, 16),
48528 => conv_std_logic_vector(27216, 16),
48529 => conv_std_logic_vector(27405, 16),
48530 => conv_std_logic_vector(27594, 16),
48531 => conv_std_logic_vector(27783, 16),
48532 => conv_std_logic_vector(27972, 16),
48533 => conv_std_logic_vector(28161, 16),
48534 => conv_std_logic_vector(28350, 16),
48535 => conv_std_logic_vector(28539, 16),
48536 => conv_std_logic_vector(28728, 16),
48537 => conv_std_logic_vector(28917, 16),
48538 => conv_std_logic_vector(29106, 16),
48539 => conv_std_logic_vector(29295, 16),
48540 => conv_std_logic_vector(29484, 16),
48541 => conv_std_logic_vector(29673, 16),
48542 => conv_std_logic_vector(29862, 16),
48543 => conv_std_logic_vector(30051, 16),
48544 => conv_std_logic_vector(30240, 16),
48545 => conv_std_logic_vector(30429, 16),
48546 => conv_std_logic_vector(30618, 16),
48547 => conv_std_logic_vector(30807, 16),
48548 => conv_std_logic_vector(30996, 16),
48549 => conv_std_logic_vector(31185, 16),
48550 => conv_std_logic_vector(31374, 16),
48551 => conv_std_logic_vector(31563, 16),
48552 => conv_std_logic_vector(31752, 16),
48553 => conv_std_logic_vector(31941, 16),
48554 => conv_std_logic_vector(32130, 16),
48555 => conv_std_logic_vector(32319, 16),
48556 => conv_std_logic_vector(32508, 16),
48557 => conv_std_logic_vector(32697, 16),
48558 => conv_std_logic_vector(32886, 16),
48559 => conv_std_logic_vector(33075, 16),
48560 => conv_std_logic_vector(33264, 16),
48561 => conv_std_logic_vector(33453, 16),
48562 => conv_std_logic_vector(33642, 16),
48563 => conv_std_logic_vector(33831, 16),
48564 => conv_std_logic_vector(34020, 16),
48565 => conv_std_logic_vector(34209, 16),
48566 => conv_std_logic_vector(34398, 16),
48567 => conv_std_logic_vector(34587, 16),
48568 => conv_std_logic_vector(34776, 16),
48569 => conv_std_logic_vector(34965, 16),
48570 => conv_std_logic_vector(35154, 16),
48571 => conv_std_logic_vector(35343, 16),
48572 => conv_std_logic_vector(35532, 16),
48573 => conv_std_logic_vector(35721, 16),
48574 => conv_std_logic_vector(35910, 16),
48575 => conv_std_logic_vector(36099, 16),
48576 => conv_std_logic_vector(36288, 16),
48577 => conv_std_logic_vector(36477, 16),
48578 => conv_std_logic_vector(36666, 16),
48579 => conv_std_logic_vector(36855, 16),
48580 => conv_std_logic_vector(37044, 16),
48581 => conv_std_logic_vector(37233, 16),
48582 => conv_std_logic_vector(37422, 16),
48583 => conv_std_logic_vector(37611, 16),
48584 => conv_std_logic_vector(37800, 16),
48585 => conv_std_logic_vector(37989, 16),
48586 => conv_std_logic_vector(38178, 16),
48587 => conv_std_logic_vector(38367, 16),
48588 => conv_std_logic_vector(38556, 16),
48589 => conv_std_logic_vector(38745, 16),
48590 => conv_std_logic_vector(38934, 16),
48591 => conv_std_logic_vector(39123, 16),
48592 => conv_std_logic_vector(39312, 16),
48593 => conv_std_logic_vector(39501, 16),
48594 => conv_std_logic_vector(39690, 16),
48595 => conv_std_logic_vector(39879, 16),
48596 => conv_std_logic_vector(40068, 16),
48597 => conv_std_logic_vector(40257, 16),
48598 => conv_std_logic_vector(40446, 16),
48599 => conv_std_logic_vector(40635, 16),
48600 => conv_std_logic_vector(40824, 16),
48601 => conv_std_logic_vector(41013, 16),
48602 => conv_std_logic_vector(41202, 16),
48603 => conv_std_logic_vector(41391, 16),
48604 => conv_std_logic_vector(41580, 16),
48605 => conv_std_logic_vector(41769, 16),
48606 => conv_std_logic_vector(41958, 16),
48607 => conv_std_logic_vector(42147, 16),
48608 => conv_std_logic_vector(42336, 16),
48609 => conv_std_logic_vector(42525, 16),
48610 => conv_std_logic_vector(42714, 16),
48611 => conv_std_logic_vector(42903, 16),
48612 => conv_std_logic_vector(43092, 16),
48613 => conv_std_logic_vector(43281, 16),
48614 => conv_std_logic_vector(43470, 16),
48615 => conv_std_logic_vector(43659, 16),
48616 => conv_std_logic_vector(43848, 16),
48617 => conv_std_logic_vector(44037, 16),
48618 => conv_std_logic_vector(44226, 16),
48619 => conv_std_logic_vector(44415, 16),
48620 => conv_std_logic_vector(44604, 16),
48621 => conv_std_logic_vector(44793, 16),
48622 => conv_std_logic_vector(44982, 16),
48623 => conv_std_logic_vector(45171, 16),
48624 => conv_std_logic_vector(45360, 16),
48625 => conv_std_logic_vector(45549, 16),
48626 => conv_std_logic_vector(45738, 16),
48627 => conv_std_logic_vector(45927, 16),
48628 => conv_std_logic_vector(46116, 16),
48629 => conv_std_logic_vector(46305, 16),
48630 => conv_std_logic_vector(46494, 16),
48631 => conv_std_logic_vector(46683, 16),
48632 => conv_std_logic_vector(46872, 16),
48633 => conv_std_logic_vector(47061, 16),
48634 => conv_std_logic_vector(47250, 16),
48635 => conv_std_logic_vector(47439, 16),
48636 => conv_std_logic_vector(47628, 16),
48637 => conv_std_logic_vector(47817, 16),
48638 => conv_std_logic_vector(48006, 16),
48639 => conv_std_logic_vector(48195, 16),
48640 => conv_std_logic_vector(0, 16),
48641 => conv_std_logic_vector(190, 16),
48642 => conv_std_logic_vector(380, 16),
48643 => conv_std_logic_vector(570, 16),
48644 => conv_std_logic_vector(760, 16),
48645 => conv_std_logic_vector(950, 16),
48646 => conv_std_logic_vector(1140, 16),
48647 => conv_std_logic_vector(1330, 16),
48648 => conv_std_logic_vector(1520, 16),
48649 => conv_std_logic_vector(1710, 16),
48650 => conv_std_logic_vector(1900, 16),
48651 => conv_std_logic_vector(2090, 16),
48652 => conv_std_logic_vector(2280, 16),
48653 => conv_std_logic_vector(2470, 16),
48654 => conv_std_logic_vector(2660, 16),
48655 => conv_std_logic_vector(2850, 16),
48656 => conv_std_logic_vector(3040, 16),
48657 => conv_std_logic_vector(3230, 16),
48658 => conv_std_logic_vector(3420, 16),
48659 => conv_std_logic_vector(3610, 16),
48660 => conv_std_logic_vector(3800, 16),
48661 => conv_std_logic_vector(3990, 16),
48662 => conv_std_logic_vector(4180, 16),
48663 => conv_std_logic_vector(4370, 16),
48664 => conv_std_logic_vector(4560, 16),
48665 => conv_std_logic_vector(4750, 16),
48666 => conv_std_logic_vector(4940, 16),
48667 => conv_std_logic_vector(5130, 16),
48668 => conv_std_logic_vector(5320, 16),
48669 => conv_std_logic_vector(5510, 16),
48670 => conv_std_logic_vector(5700, 16),
48671 => conv_std_logic_vector(5890, 16),
48672 => conv_std_logic_vector(6080, 16),
48673 => conv_std_logic_vector(6270, 16),
48674 => conv_std_logic_vector(6460, 16),
48675 => conv_std_logic_vector(6650, 16),
48676 => conv_std_logic_vector(6840, 16),
48677 => conv_std_logic_vector(7030, 16),
48678 => conv_std_logic_vector(7220, 16),
48679 => conv_std_logic_vector(7410, 16),
48680 => conv_std_logic_vector(7600, 16),
48681 => conv_std_logic_vector(7790, 16),
48682 => conv_std_logic_vector(7980, 16),
48683 => conv_std_logic_vector(8170, 16),
48684 => conv_std_logic_vector(8360, 16),
48685 => conv_std_logic_vector(8550, 16),
48686 => conv_std_logic_vector(8740, 16),
48687 => conv_std_logic_vector(8930, 16),
48688 => conv_std_logic_vector(9120, 16),
48689 => conv_std_logic_vector(9310, 16),
48690 => conv_std_logic_vector(9500, 16),
48691 => conv_std_logic_vector(9690, 16),
48692 => conv_std_logic_vector(9880, 16),
48693 => conv_std_logic_vector(10070, 16),
48694 => conv_std_logic_vector(10260, 16),
48695 => conv_std_logic_vector(10450, 16),
48696 => conv_std_logic_vector(10640, 16),
48697 => conv_std_logic_vector(10830, 16),
48698 => conv_std_logic_vector(11020, 16),
48699 => conv_std_logic_vector(11210, 16),
48700 => conv_std_logic_vector(11400, 16),
48701 => conv_std_logic_vector(11590, 16),
48702 => conv_std_logic_vector(11780, 16),
48703 => conv_std_logic_vector(11970, 16),
48704 => conv_std_logic_vector(12160, 16),
48705 => conv_std_logic_vector(12350, 16),
48706 => conv_std_logic_vector(12540, 16),
48707 => conv_std_logic_vector(12730, 16),
48708 => conv_std_logic_vector(12920, 16),
48709 => conv_std_logic_vector(13110, 16),
48710 => conv_std_logic_vector(13300, 16),
48711 => conv_std_logic_vector(13490, 16),
48712 => conv_std_logic_vector(13680, 16),
48713 => conv_std_logic_vector(13870, 16),
48714 => conv_std_logic_vector(14060, 16),
48715 => conv_std_logic_vector(14250, 16),
48716 => conv_std_logic_vector(14440, 16),
48717 => conv_std_logic_vector(14630, 16),
48718 => conv_std_logic_vector(14820, 16),
48719 => conv_std_logic_vector(15010, 16),
48720 => conv_std_logic_vector(15200, 16),
48721 => conv_std_logic_vector(15390, 16),
48722 => conv_std_logic_vector(15580, 16),
48723 => conv_std_logic_vector(15770, 16),
48724 => conv_std_logic_vector(15960, 16),
48725 => conv_std_logic_vector(16150, 16),
48726 => conv_std_logic_vector(16340, 16),
48727 => conv_std_logic_vector(16530, 16),
48728 => conv_std_logic_vector(16720, 16),
48729 => conv_std_logic_vector(16910, 16),
48730 => conv_std_logic_vector(17100, 16),
48731 => conv_std_logic_vector(17290, 16),
48732 => conv_std_logic_vector(17480, 16),
48733 => conv_std_logic_vector(17670, 16),
48734 => conv_std_logic_vector(17860, 16),
48735 => conv_std_logic_vector(18050, 16),
48736 => conv_std_logic_vector(18240, 16),
48737 => conv_std_logic_vector(18430, 16),
48738 => conv_std_logic_vector(18620, 16),
48739 => conv_std_logic_vector(18810, 16),
48740 => conv_std_logic_vector(19000, 16),
48741 => conv_std_logic_vector(19190, 16),
48742 => conv_std_logic_vector(19380, 16),
48743 => conv_std_logic_vector(19570, 16),
48744 => conv_std_logic_vector(19760, 16),
48745 => conv_std_logic_vector(19950, 16),
48746 => conv_std_logic_vector(20140, 16),
48747 => conv_std_logic_vector(20330, 16),
48748 => conv_std_logic_vector(20520, 16),
48749 => conv_std_logic_vector(20710, 16),
48750 => conv_std_logic_vector(20900, 16),
48751 => conv_std_logic_vector(21090, 16),
48752 => conv_std_logic_vector(21280, 16),
48753 => conv_std_logic_vector(21470, 16),
48754 => conv_std_logic_vector(21660, 16),
48755 => conv_std_logic_vector(21850, 16),
48756 => conv_std_logic_vector(22040, 16),
48757 => conv_std_logic_vector(22230, 16),
48758 => conv_std_logic_vector(22420, 16),
48759 => conv_std_logic_vector(22610, 16),
48760 => conv_std_logic_vector(22800, 16),
48761 => conv_std_logic_vector(22990, 16),
48762 => conv_std_logic_vector(23180, 16),
48763 => conv_std_logic_vector(23370, 16),
48764 => conv_std_logic_vector(23560, 16),
48765 => conv_std_logic_vector(23750, 16),
48766 => conv_std_logic_vector(23940, 16),
48767 => conv_std_logic_vector(24130, 16),
48768 => conv_std_logic_vector(24320, 16),
48769 => conv_std_logic_vector(24510, 16),
48770 => conv_std_logic_vector(24700, 16),
48771 => conv_std_logic_vector(24890, 16),
48772 => conv_std_logic_vector(25080, 16),
48773 => conv_std_logic_vector(25270, 16),
48774 => conv_std_logic_vector(25460, 16),
48775 => conv_std_logic_vector(25650, 16),
48776 => conv_std_logic_vector(25840, 16),
48777 => conv_std_logic_vector(26030, 16),
48778 => conv_std_logic_vector(26220, 16),
48779 => conv_std_logic_vector(26410, 16),
48780 => conv_std_logic_vector(26600, 16),
48781 => conv_std_logic_vector(26790, 16),
48782 => conv_std_logic_vector(26980, 16),
48783 => conv_std_logic_vector(27170, 16),
48784 => conv_std_logic_vector(27360, 16),
48785 => conv_std_logic_vector(27550, 16),
48786 => conv_std_logic_vector(27740, 16),
48787 => conv_std_logic_vector(27930, 16),
48788 => conv_std_logic_vector(28120, 16),
48789 => conv_std_logic_vector(28310, 16),
48790 => conv_std_logic_vector(28500, 16),
48791 => conv_std_logic_vector(28690, 16),
48792 => conv_std_logic_vector(28880, 16),
48793 => conv_std_logic_vector(29070, 16),
48794 => conv_std_logic_vector(29260, 16),
48795 => conv_std_logic_vector(29450, 16),
48796 => conv_std_logic_vector(29640, 16),
48797 => conv_std_logic_vector(29830, 16),
48798 => conv_std_logic_vector(30020, 16),
48799 => conv_std_logic_vector(30210, 16),
48800 => conv_std_logic_vector(30400, 16),
48801 => conv_std_logic_vector(30590, 16),
48802 => conv_std_logic_vector(30780, 16),
48803 => conv_std_logic_vector(30970, 16),
48804 => conv_std_logic_vector(31160, 16),
48805 => conv_std_logic_vector(31350, 16),
48806 => conv_std_logic_vector(31540, 16),
48807 => conv_std_logic_vector(31730, 16),
48808 => conv_std_logic_vector(31920, 16),
48809 => conv_std_logic_vector(32110, 16),
48810 => conv_std_logic_vector(32300, 16),
48811 => conv_std_logic_vector(32490, 16),
48812 => conv_std_logic_vector(32680, 16),
48813 => conv_std_logic_vector(32870, 16),
48814 => conv_std_logic_vector(33060, 16),
48815 => conv_std_logic_vector(33250, 16),
48816 => conv_std_logic_vector(33440, 16),
48817 => conv_std_logic_vector(33630, 16),
48818 => conv_std_logic_vector(33820, 16),
48819 => conv_std_logic_vector(34010, 16),
48820 => conv_std_logic_vector(34200, 16),
48821 => conv_std_logic_vector(34390, 16),
48822 => conv_std_logic_vector(34580, 16),
48823 => conv_std_logic_vector(34770, 16),
48824 => conv_std_logic_vector(34960, 16),
48825 => conv_std_logic_vector(35150, 16),
48826 => conv_std_logic_vector(35340, 16),
48827 => conv_std_logic_vector(35530, 16),
48828 => conv_std_logic_vector(35720, 16),
48829 => conv_std_logic_vector(35910, 16),
48830 => conv_std_logic_vector(36100, 16),
48831 => conv_std_logic_vector(36290, 16),
48832 => conv_std_logic_vector(36480, 16),
48833 => conv_std_logic_vector(36670, 16),
48834 => conv_std_logic_vector(36860, 16),
48835 => conv_std_logic_vector(37050, 16),
48836 => conv_std_logic_vector(37240, 16),
48837 => conv_std_logic_vector(37430, 16),
48838 => conv_std_logic_vector(37620, 16),
48839 => conv_std_logic_vector(37810, 16),
48840 => conv_std_logic_vector(38000, 16),
48841 => conv_std_logic_vector(38190, 16),
48842 => conv_std_logic_vector(38380, 16),
48843 => conv_std_logic_vector(38570, 16),
48844 => conv_std_logic_vector(38760, 16),
48845 => conv_std_logic_vector(38950, 16),
48846 => conv_std_logic_vector(39140, 16),
48847 => conv_std_logic_vector(39330, 16),
48848 => conv_std_logic_vector(39520, 16),
48849 => conv_std_logic_vector(39710, 16),
48850 => conv_std_logic_vector(39900, 16),
48851 => conv_std_logic_vector(40090, 16),
48852 => conv_std_logic_vector(40280, 16),
48853 => conv_std_logic_vector(40470, 16),
48854 => conv_std_logic_vector(40660, 16),
48855 => conv_std_logic_vector(40850, 16),
48856 => conv_std_logic_vector(41040, 16),
48857 => conv_std_logic_vector(41230, 16),
48858 => conv_std_logic_vector(41420, 16),
48859 => conv_std_logic_vector(41610, 16),
48860 => conv_std_logic_vector(41800, 16),
48861 => conv_std_logic_vector(41990, 16),
48862 => conv_std_logic_vector(42180, 16),
48863 => conv_std_logic_vector(42370, 16),
48864 => conv_std_logic_vector(42560, 16),
48865 => conv_std_logic_vector(42750, 16),
48866 => conv_std_logic_vector(42940, 16),
48867 => conv_std_logic_vector(43130, 16),
48868 => conv_std_logic_vector(43320, 16),
48869 => conv_std_logic_vector(43510, 16),
48870 => conv_std_logic_vector(43700, 16),
48871 => conv_std_logic_vector(43890, 16),
48872 => conv_std_logic_vector(44080, 16),
48873 => conv_std_logic_vector(44270, 16),
48874 => conv_std_logic_vector(44460, 16),
48875 => conv_std_logic_vector(44650, 16),
48876 => conv_std_logic_vector(44840, 16),
48877 => conv_std_logic_vector(45030, 16),
48878 => conv_std_logic_vector(45220, 16),
48879 => conv_std_logic_vector(45410, 16),
48880 => conv_std_logic_vector(45600, 16),
48881 => conv_std_logic_vector(45790, 16),
48882 => conv_std_logic_vector(45980, 16),
48883 => conv_std_logic_vector(46170, 16),
48884 => conv_std_logic_vector(46360, 16),
48885 => conv_std_logic_vector(46550, 16),
48886 => conv_std_logic_vector(46740, 16),
48887 => conv_std_logic_vector(46930, 16),
48888 => conv_std_logic_vector(47120, 16),
48889 => conv_std_logic_vector(47310, 16),
48890 => conv_std_logic_vector(47500, 16),
48891 => conv_std_logic_vector(47690, 16),
48892 => conv_std_logic_vector(47880, 16),
48893 => conv_std_logic_vector(48070, 16),
48894 => conv_std_logic_vector(48260, 16),
48895 => conv_std_logic_vector(48450, 16),
48896 => conv_std_logic_vector(0, 16),
48897 => conv_std_logic_vector(191, 16),
48898 => conv_std_logic_vector(382, 16),
48899 => conv_std_logic_vector(573, 16),
48900 => conv_std_logic_vector(764, 16),
48901 => conv_std_logic_vector(955, 16),
48902 => conv_std_logic_vector(1146, 16),
48903 => conv_std_logic_vector(1337, 16),
48904 => conv_std_logic_vector(1528, 16),
48905 => conv_std_logic_vector(1719, 16),
48906 => conv_std_logic_vector(1910, 16),
48907 => conv_std_logic_vector(2101, 16),
48908 => conv_std_logic_vector(2292, 16),
48909 => conv_std_logic_vector(2483, 16),
48910 => conv_std_logic_vector(2674, 16),
48911 => conv_std_logic_vector(2865, 16),
48912 => conv_std_logic_vector(3056, 16),
48913 => conv_std_logic_vector(3247, 16),
48914 => conv_std_logic_vector(3438, 16),
48915 => conv_std_logic_vector(3629, 16),
48916 => conv_std_logic_vector(3820, 16),
48917 => conv_std_logic_vector(4011, 16),
48918 => conv_std_logic_vector(4202, 16),
48919 => conv_std_logic_vector(4393, 16),
48920 => conv_std_logic_vector(4584, 16),
48921 => conv_std_logic_vector(4775, 16),
48922 => conv_std_logic_vector(4966, 16),
48923 => conv_std_logic_vector(5157, 16),
48924 => conv_std_logic_vector(5348, 16),
48925 => conv_std_logic_vector(5539, 16),
48926 => conv_std_logic_vector(5730, 16),
48927 => conv_std_logic_vector(5921, 16),
48928 => conv_std_logic_vector(6112, 16),
48929 => conv_std_logic_vector(6303, 16),
48930 => conv_std_logic_vector(6494, 16),
48931 => conv_std_logic_vector(6685, 16),
48932 => conv_std_logic_vector(6876, 16),
48933 => conv_std_logic_vector(7067, 16),
48934 => conv_std_logic_vector(7258, 16),
48935 => conv_std_logic_vector(7449, 16),
48936 => conv_std_logic_vector(7640, 16),
48937 => conv_std_logic_vector(7831, 16),
48938 => conv_std_logic_vector(8022, 16),
48939 => conv_std_logic_vector(8213, 16),
48940 => conv_std_logic_vector(8404, 16),
48941 => conv_std_logic_vector(8595, 16),
48942 => conv_std_logic_vector(8786, 16),
48943 => conv_std_logic_vector(8977, 16),
48944 => conv_std_logic_vector(9168, 16),
48945 => conv_std_logic_vector(9359, 16),
48946 => conv_std_logic_vector(9550, 16),
48947 => conv_std_logic_vector(9741, 16),
48948 => conv_std_logic_vector(9932, 16),
48949 => conv_std_logic_vector(10123, 16),
48950 => conv_std_logic_vector(10314, 16),
48951 => conv_std_logic_vector(10505, 16),
48952 => conv_std_logic_vector(10696, 16),
48953 => conv_std_logic_vector(10887, 16),
48954 => conv_std_logic_vector(11078, 16),
48955 => conv_std_logic_vector(11269, 16),
48956 => conv_std_logic_vector(11460, 16),
48957 => conv_std_logic_vector(11651, 16),
48958 => conv_std_logic_vector(11842, 16),
48959 => conv_std_logic_vector(12033, 16),
48960 => conv_std_logic_vector(12224, 16),
48961 => conv_std_logic_vector(12415, 16),
48962 => conv_std_logic_vector(12606, 16),
48963 => conv_std_logic_vector(12797, 16),
48964 => conv_std_logic_vector(12988, 16),
48965 => conv_std_logic_vector(13179, 16),
48966 => conv_std_logic_vector(13370, 16),
48967 => conv_std_logic_vector(13561, 16),
48968 => conv_std_logic_vector(13752, 16),
48969 => conv_std_logic_vector(13943, 16),
48970 => conv_std_logic_vector(14134, 16),
48971 => conv_std_logic_vector(14325, 16),
48972 => conv_std_logic_vector(14516, 16),
48973 => conv_std_logic_vector(14707, 16),
48974 => conv_std_logic_vector(14898, 16),
48975 => conv_std_logic_vector(15089, 16),
48976 => conv_std_logic_vector(15280, 16),
48977 => conv_std_logic_vector(15471, 16),
48978 => conv_std_logic_vector(15662, 16),
48979 => conv_std_logic_vector(15853, 16),
48980 => conv_std_logic_vector(16044, 16),
48981 => conv_std_logic_vector(16235, 16),
48982 => conv_std_logic_vector(16426, 16),
48983 => conv_std_logic_vector(16617, 16),
48984 => conv_std_logic_vector(16808, 16),
48985 => conv_std_logic_vector(16999, 16),
48986 => conv_std_logic_vector(17190, 16),
48987 => conv_std_logic_vector(17381, 16),
48988 => conv_std_logic_vector(17572, 16),
48989 => conv_std_logic_vector(17763, 16),
48990 => conv_std_logic_vector(17954, 16),
48991 => conv_std_logic_vector(18145, 16),
48992 => conv_std_logic_vector(18336, 16),
48993 => conv_std_logic_vector(18527, 16),
48994 => conv_std_logic_vector(18718, 16),
48995 => conv_std_logic_vector(18909, 16),
48996 => conv_std_logic_vector(19100, 16),
48997 => conv_std_logic_vector(19291, 16),
48998 => conv_std_logic_vector(19482, 16),
48999 => conv_std_logic_vector(19673, 16),
49000 => conv_std_logic_vector(19864, 16),
49001 => conv_std_logic_vector(20055, 16),
49002 => conv_std_logic_vector(20246, 16),
49003 => conv_std_logic_vector(20437, 16),
49004 => conv_std_logic_vector(20628, 16),
49005 => conv_std_logic_vector(20819, 16),
49006 => conv_std_logic_vector(21010, 16),
49007 => conv_std_logic_vector(21201, 16),
49008 => conv_std_logic_vector(21392, 16),
49009 => conv_std_logic_vector(21583, 16),
49010 => conv_std_logic_vector(21774, 16),
49011 => conv_std_logic_vector(21965, 16),
49012 => conv_std_logic_vector(22156, 16),
49013 => conv_std_logic_vector(22347, 16),
49014 => conv_std_logic_vector(22538, 16),
49015 => conv_std_logic_vector(22729, 16),
49016 => conv_std_logic_vector(22920, 16),
49017 => conv_std_logic_vector(23111, 16),
49018 => conv_std_logic_vector(23302, 16),
49019 => conv_std_logic_vector(23493, 16),
49020 => conv_std_logic_vector(23684, 16),
49021 => conv_std_logic_vector(23875, 16),
49022 => conv_std_logic_vector(24066, 16),
49023 => conv_std_logic_vector(24257, 16),
49024 => conv_std_logic_vector(24448, 16),
49025 => conv_std_logic_vector(24639, 16),
49026 => conv_std_logic_vector(24830, 16),
49027 => conv_std_logic_vector(25021, 16),
49028 => conv_std_logic_vector(25212, 16),
49029 => conv_std_logic_vector(25403, 16),
49030 => conv_std_logic_vector(25594, 16),
49031 => conv_std_logic_vector(25785, 16),
49032 => conv_std_logic_vector(25976, 16),
49033 => conv_std_logic_vector(26167, 16),
49034 => conv_std_logic_vector(26358, 16),
49035 => conv_std_logic_vector(26549, 16),
49036 => conv_std_logic_vector(26740, 16),
49037 => conv_std_logic_vector(26931, 16),
49038 => conv_std_logic_vector(27122, 16),
49039 => conv_std_logic_vector(27313, 16),
49040 => conv_std_logic_vector(27504, 16),
49041 => conv_std_logic_vector(27695, 16),
49042 => conv_std_logic_vector(27886, 16),
49043 => conv_std_logic_vector(28077, 16),
49044 => conv_std_logic_vector(28268, 16),
49045 => conv_std_logic_vector(28459, 16),
49046 => conv_std_logic_vector(28650, 16),
49047 => conv_std_logic_vector(28841, 16),
49048 => conv_std_logic_vector(29032, 16),
49049 => conv_std_logic_vector(29223, 16),
49050 => conv_std_logic_vector(29414, 16),
49051 => conv_std_logic_vector(29605, 16),
49052 => conv_std_logic_vector(29796, 16),
49053 => conv_std_logic_vector(29987, 16),
49054 => conv_std_logic_vector(30178, 16),
49055 => conv_std_logic_vector(30369, 16),
49056 => conv_std_logic_vector(30560, 16),
49057 => conv_std_logic_vector(30751, 16),
49058 => conv_std_logic_vector(30942, 16),
49059 => conv_std_logic_vector(31133, 16),
49060 => conv_std_logic_vector(31324, 16),
49061 => conv_std_logic_vector(31515, 16),
49062 => conv_std_logic_vector(31706, 16),
49063 => conv_std_logic_vector(31897, 16),
49064 => conv_std_logic_vector(32088, 16),
49065 => conv_std_logic_vector(32279, 16),
49066 => conv_std_logic_vector(32470, 16),
49067 => conv_std_logic_vector(32661, 16),
49068 => conv_std_logic_vector(32852, 16),
49069 => conv_std_logic_vector(33043, 16),
49070 => conv_std_logic_vector(33234, 16),
49071 => conv_std_logic_vector(33425, 16),
49072 => conv_std_logic_vector(33616, 16),
49073 => conv_std_logic_vector(33807, 16),
49074 => conv_std_logic_vector(33998, 16),
49075 => conv_std_logic_vector(34189, 16),
49076 => conv_std_logic_vector(34380, 16),
49077 => conv_std_logic_vector(34571, 16),
49078 => conv_std_logic_vector(34762, 16),
49079 => conv_std_logic_vector(34953, 16),
49080 => conv_std_logic_vector(35144, 16),
49081 => conv_std_logic_vector(35335, 16),
49082 => conv_std_logic_vector(35526, 16),
49083 => conv_std_logic_vector(35717, 16),
49084 => conv_std_logic_vector(35908, 16),
49085 => conv_std_logic_vector(36099, 16),
49086 => conv_std_logic_vector(36290, 16),
49087 => conv_std_logic_vector(36481, 16),
49088 => conv_std_logic_vector(36672, 16),
49089 => conv_std_logic_vector(36863, 16),
49090 => conv_std_logic_vector(37054, 16),
49091 => conv_std_logic_vector(37245, 16),
49092 => conv_std_logic_vector(37436, 16),
49093 => conv_std_logic_vector(37627, 16),
49094 => conv_std_logic_vector(37818, 16),
49095 => conv_std_logic_vector(38009, 16),
49096 => conv_std_logic_vector(38200, 16),
49097 => conv_std_logic_vector(38391, 16),
49098 => conv_std_logic_vector(38582, 16),
49099 => conv_std_logic_vector(38773, 16),
49100 => conv_std_logic_vector(38964, 16),
49101 => conv_std_logic_vector(39155, 16),
49102 => conv_std_logic_vector(39346, 16),
49103 => conv_std_logic_vector(39537, 16),
49104 => conv_std_logic_vector(39728, 16),
49105 => conv_std_logic_vector(39919, 16),
49106 => conv_std_logic_vector(40110, 16),
49107 => conv_std_logic_vector(40301, 16),
49108 => conv_std_logic_vector(40492, 16),
49109 => conv_std_logic_vector(40683, 16),
49110 => conv_std_logic_vector(40874, 16),
49111 => conv_std_logic_vector(41065, 16),
49112 => conv_std_logic_vector(41256, 16),
49113 => conv_std_logic_vector(41447, 16),
49114 => conv_std_logic_vector(41638, 16),
49115 => conv_std_logic_vector(41829, 16),
49116 => conv_std_logic_vector(42020, 16),
49117 => conv_std_logic_vector(42211, 16),
49118 => conv_std_logic_vector(42402, 16),
49119 => conv_std_logic_vector(42593, 16),
49120 => conv_std_logic_vector(42784, 16),
49121 => conv_std_logic_vector(42975, 16),
49122 => conv_std_logic_vector(43166, 16),
49123 => conv_std_logic_vector(43357, 16),
49124 => conv_std_logic_vector(43548, 16),
49125 => conv_std_logic_vector(43739, 16),
49126 => conv_std_logic_vector(43930, 16),
49127 => conv_std_logic_vector(44121, 16),
49128 => conv_std_logic_vector(44312, 16),
49129 => conv_std_logic_vector(44503, 16),
49130 => conv_std_logic_vector(44694, 16),
49131 => conv_std_logic_vector(44885, 16),
49132 => conv_std_logic_vector(45076, 16),
49133 => conv_std_logic_vector(45267, 16),
49134 => conv_std_logic_vector(45458, 16),
49135 => conv_std_logic_vector(45649, 16),
49136 => conv_std_logic_vector(45840, 16),
49137 => conv_std_logic_vector(46031, 16),
49138 => conv_std_logic_vector(46222, 16),
49139 => conv_std_logic_vector(46413, 16),
49140 => conv_std_logic_vector(46604, 16),
49141 => conv_std_logic_vector(46795, 16),
49142 => conv_std_logic_vector(46986, 16),
49143 => conv_std_logic_vector(47177, 16),
49144 => conv_std_logic_vector(47368, 16),
49145 => conv_std_logic_vector(47559, 16),
49146 => conv_std_logic_vector(47750, 16),
49147 => conv_std_logic_vector(47941, 16),
49148 => conv_std_logic_vector(48132, 16),
49149 => conv_std_logic_vector(48323, 16),
49150 => conv_std_logic_vector(48514, 16),
49151 => conv_std_logic_vector(48705, 16),
49152 => conv_std_logic_vector(0, 16),
49153 => conv_std_logic_vector(192, 16),
49154 => conv_std_logic_vector(384, 16),
49155 => conv_std_logic_vector(576, 16),
49156 => conv_std_logic_vector(768, 16),
49157 => conv_std_logic_vector(960, 16),
49158 => conv_std_logic_vector(1152, 16),
49159 => conv_std_logic_vector(1344, 16),
49160 => conv_std_logic_vector(1536, 16),
49161 => conv_std_logic_vector(1728, 16),
49162 => conv_std_logic_vector(1920, 16),
49163 => conv_std_logic_vector(2112, 16),
49164 => conv_std_logic_vector(2304, 16),
49165 => conv_std_logic_vector(2496, 16),
49166 => conv_std_logic_vector(2688, 16),
49167 => conv_std_logic_vector(2880, 16),
49168 => conv_std_logic_vector(3072, 16),
49169 => conv_std_logic_vector(3264, 16),
49170 => conv_std_logic_vector(3456, 16),
49171 => conv_std_logic_vector(3648, 16),
49172 => conv_std_logic_vector(3840, 16),
49173 => conv_std_logic_vector(4032, 16),
49174 => conv_std_logic_vector(4224, 16),
49175 => conv_std_logic_vector(4416, 16),
49176 => conv_std_logic_vector(4608, 16),
49177 => conv_std_logic_vector(4800, 16),
49178 => conv_std_logic_vector(4992, 16),
49179 => conv_std_logic_vector(5184, 16),
49180 => conv_std_logic_vector(5376, 16),
49181 => conv_std_logic_vector(5568, 16),
49182 => conv_std_logic_vector(5760, 16),
49183 => conv_std_logic_vector(5952, 16),
49184 => conv_std_logic_vector(6144, 16),
49185 => conv_std_logic_vector(6336, 16),
49186 => conv_std_logic_vector(6528, 16),
49187 => conv_std_logic_vector(6720, 16),
49188 => conv_std_logic_vector(6912, 16),
49189 => conv_std_logic_vector(7104, 16),
49190 => conv_std_logic_vector(7296, 16),
49191 => conv_std_logic_vector(7488, 16),
49192 => conv_std_logic_vector(7680, 16),
49193 => conv_std_logic_vector(7872, 16),
49194 => conv_std_logic_vector(8064, 16),
49195 => conv_std_logic_vector(8256, 16),
49196 => conv_std_logic_vector(8448, 16),
49197 => conv_std_logic_vector(8640, 16),
49198 => conv_std_logic_vector(8832, 16),
49199 => conv_std_logic_vector(9024, 16),
49200 => conv_std_logic_vector(9216, 16),
49201 => conv_std_logic_vector(9408, 16),
49202 => conv_std_logic_vector(9600, 16),
49203 => conv_std_logic_vector(9792, 16),
49204 => conv_std_logic_vector(9984, 16),
49205 => conv_std_logic_vector(10176, 16),
49206 => conv_std_logic_vector(10368, 16),
49207 => conv_std_logic_vector(10560, 16),
49208 => conv_std_logic_vector(10752, 16),
49209 => conv_std_logic_vector(10944, 16),
49210 => conv_std_logic_vector(11136, 16),
49211 => conv_std_logic_vector(11328, 16),
49212 => conv_std_logic_vector(11520, 16),
49213 => conv_std_logic_vector(11712, 16),
49214 => conv_std_logic_vector(11904, 16),
49215 => conv_std_logic_vector(12096, 16),
49216 => conv_std_logic_vector(12288, 16),
49217 => conv_std_logic_vector(12480, 16),
49218 => conv_std_logic_vector(12672, 16),
49219 => conv_std_logic_vector(12864, 16),
49220 => conv_std_logic_vector(13056, 16),
49221 => conv_std_logic_vector(13248, 16),
49222 => conv_std_logic_vector(13440, 16),
49223 => conv_std_logic_vector(13632, 16),
49224 => conv_std_logic_vector(13824, 16),
49225 => conv_std_logic_vector(14016, 16),
49226 => conv_std_logic_vector(14208, 16),
49227 => conv_std_logic_vector(14400, 16),
49228 => conv_std_logic_vector(14592, 16),
49229 => conv_std_logic_vector(14784, 16),
49230 => conv_std_logic_vector(14976, 16),
49231 => conv_std_logic_vector(15168, 16),
49232 => conv_std_logic_vector(15360, 16),
49233 => conv_std_logic_vector(15552, 16),
49234 => conv_std_logic_vector(15744, 16),
49235 => conv_std_logic_vector(15936, 16),
49236 => conv_std_logic_vector(16128, 16),
49237 => conv_std_logic_vector(16320, 16),
49238 => conv_std_logic_vector(16512, 16),
49239 => conv_std_logic_vector(16704, 16),
49240 => conv_std_logic_vector(16896, 16),
49241 => conv_std_logic_vector(17088, 16),
49242 => conv_std_logic_vector(17280, 16),
49243 => conv_std_logic_vector(17472, 16),
49244 => conv_std_logic_vector(17664, 16),
49245 => conv_std_logic_vector(17856, 16),
49246 => conv_std_logic_vector(18048, 16),
49247 => conv_std_logic_vector(18240, 16),
49248 => conv_std_logic_vector(18432, 16),
49249 => conv_std_logic_vector(18624, 16),
49250 => conv_std_logic_vector(18816, 16),
49251 => conv_std_logic_vector(19008, 16),
49252 => conv_std_logic_vector(19200, 16),
49253 => conv_std_logic_vector(19392, 16),
49254 => conv_std_logic_vector(19584, 16),
49255 => conv_std_logic_vector(19776, 16),
49256 => conv_std_logic_vector(19968, 16),
49257 => conv_std_logic_vector(20160, 16),
49258 => conv_std_logic_vector(20352, 16),
49259 => conv_std_logic_vector(20544, 16),
49260 => conv_std_logic_vector(20736, 16),
49261 => conv_std_logic_vector(20928, 16),
49262 => conv_std_logic_vector(21120, 16),
49263 => conv_std_logic_vector(21312, 16),
49264 => conv_std_logic_vector(21504, 16),
49265 => conv_std_logic_vector(21696, 16),
49266 => conv_std_logic_vector(21888, 16),
49267 => conv_std_logic_vector(22080, 16),
49268 => conv_std_logic_vector(22272, 16),
49269 => conv_std_logic_vector(22464, 16),
49270 => conv_std_logic_vector(22656, 16),
49271 => conv_std_logic_vector(22848, 16),
49272 => conv_std_logic_vector(23040, 16),
49273 => conv_std_logic_vector(23232, 16),
49274 => conv_std_logic_vector(23424, 16),
49275 => conv_std_logic_vector(23616, 16),
49276 => conv_std_logic_vector(23808, 16),
49277 => conv_std_logic_vector(24000, 16),
49278 => conv_std_logic_vector(24192, 16),
49279 => conv_std_logic_vector(24384, 16),
49280 => conv_std_logic_vector(24576, 16),
49281 => conv_std_logic_vector(24768, 16),
49282 => conv_std_logic_vector(24960, 16),
49283 => conv_std_logic_vector(25152, 16),
49284 => conv_std_logic_vector(25344, 16),
49285 => conv_std_logic_vector(25536, 16),
49286 => conv_std_logic_vector(25728, 16),
49287 => conv_std_logic_vector(25920, 16),
49288 => conv_std_logic_vector(26112, 16),
49289 => conv_std_logic_vector(26304, 16),
49290 => conv_std_logic_vector(26496, 16),
49291 => conv_std_logic_vector(26688, 16),
49292 => conv_std_logic_vector(26880, 16),
49293 => conv_std_logic_vector(27072, 16),
49294 => conv_std_logic_vector(27264, 16),
49295 => conv_std_logic_vector(27456, 16),
49296 => conv_std_logic_vector(27648, 16),
49297 => conv_std_logic_vector(27840, 16),
49298 => conv_std_logic_vector(28032, 16),
49299 => conv_std_logic_vector(28224, 16),
49300 => conv_std_logic_vector(28416, 16),
49301 => conv_std_logic_vector(28608, 16),
49302 => conv_std_logic_vector(28800, 16),
49303 => conv_std_logic_vector(28992, 16),
49304 => conv_std_logic_vector(29184, 16),
49305 => conv_std_logic_vector(29376, 16),
49306 => conv_std_logic_vector(29568, 16),
49307 => conv_std_logic_vector(29760, 16),
49308 => conv_std_logic_vector(29952, 16),
49309 => conv_std_logic_vector(30144, 16),
49310 => conv_std_logic_vector(30336, 16),
49311 => conv_std_logic_vector(30528, 16),
49312 => conv_std_logic_vector(30720, 16),
49313 => conv_std_logic_vector(30912, 16),
49314 => conv_std_logic_vector(31104, 16),
49315 => conv_std_logic_vector(31296, 16),
49316 => conv_std_logic_vector(31488, 16),
49317 => conv_std_logic_vector(31680, 16),
49318 => conv_std_logic_vector(31872, 16),
49319 => conv_std_logic_vector(32064, 16),
49320 => conv_std_logic_vector(32256, 16),
49321 => conv_std_logic_vector(32448, 16),
49322 => conv_std_logic_vector(32640, 16),
49323 => conv_std_logic_vector(32832, 16),
49324 => conv_std_logic_vector(33024, 16),
49325 => conv_std_logic_vector(33216, 16),
49326 => conv_std_logic_vector(33408, 16),
49327 => conv_std_logic_vector(33600, 16),
49328 => conv_std_logic_vector(33792, 16),
49329 => conv_std_logic_vector(33984, 16),
49330 => conv_std_logic_vector(34176, 16),
49331 => conv_std_logic_vector(34368, 16),
49332 => conv_std_logic_vector(34560, 16),
49333 => conv_std_logic_vector(34752, 16),
49334 => conv_std_logic_vector(34944, 16),
49335 => conv_std_logic_vector(35136, 16),
49336 => conv_std_logic_vector(35328, 16),
49337 => conv_std_logic_vector(35520, 16),
49338 => conv_std_logic_vector(35712, 16),
49339 => conv_std_logic_vector(35904, 16),
49340 => conv_std_logic_vector(36096, 16),
49341 => conv_std_logic_vector(36288, 16),
49342 => conv_std_logic_vector(36480, 16),
49343 => conv_std_logic_vector(36672, 16),
49344 => conv_std_logic_vector(36864, 16),
49345 => conv_std_logic_vector(37056, 16),
49346 => conv_std_logic_vector(37248, 16),
49347 => conv_std_logic_vector(37440, 16),
49348 => conv_std_logic_vector(37632, 16),
49349 => conv_std_logic_vector(37824, 16),
49350 => conv_std_logic_vector(38016, 16),
49351 => conv_std_logic_vector(38208, 16),
49352 => conv_std_logic_vector(38400, 16),
49353 => conv_std_logic_vector(38592, 16),
49354 => conv_std_logic_vector(38784, 16),
49355 => conv_std_logic_vector(38976, 16),
49356 => conv_std_logic_vector(39168, 16),
49357 => conv_std_logic_vector(39360, 16),
49358 => conv_std_logic_vector(39552, 16),
49359 => conv_std_logic_vector(39744, 16),
49360 => conv_std_logic_vector(39936, 16),
49361 => conv_std_logic_vector(40128, 16),
49362 => conv_std_logic_vector(40320, 16),
49363 => conv_std_logic_vector(40512, 16),
49364 => conv_std_logic_vector(40704, 16),
49365 => conv_std_logic_vector(40896, 16),
49366 => conv_std_logic_vector(41088, 16),
49367 => conv_std_logic_vector(41280, 16),
49368 => conv_std_logic_vector(41472, 16),
49369 => conv_std_logic_vector(41664, 16),
49370 => conv_std_logic_vector(41856, 16),
49371 => conv_std_logic_vector(42048, 16),
49372 => conv_std_logic_vector(42240, 16),
49373 => conv_std_logic_vector(42432, 16),
49374 => conv_std_logic_vector(42624, 16),
49375 => conv_std_logic_vector(42816, 16),
49376 => conv_std_logic_vector(43008, 16),
49377 => conv_std_logic_vector(43200, 16),
49378 => conv_std_logic_vector(43392, 16),
49379 => conv_std_logic_vector(43584, 16),
49380 => conv_std_logic_vector(43776, 16),
49381 => conv_std_logic_vector(43968, 16),
49382 => conv_std_logic_vector(44160, 16),
49383 => conv_std_logic_vector(44352, 16),
49384 => conv_std_logic_vector(44544, 16),
49385 => conv_std_logic_vector(44736, 16),
49386 => conv_std_logic_vector(44928, 16),
49387 => conv_std_logic_vector(45120, 16),
49388 => conv_std_logic_vector(45312, 16),
49389 => conv_std_logic_vector(45504, 16),
49390 => conv_std_logic_vector(45696, 16),
49391 => conv_std_logic_vector(45888, 16),
49392 => conv_std_logic_vector(46080, 16),
49393 => conv_std_logic_vector(46272, 16),
49394 => conv_std_logic_vector(46464, 16),
49395 => conv_std_logic_vector(46656, 16),
49396 => conv_std_logic_vector(46848, 16),
49397 => conv_std_logic_vector(47040, 16),
49398 => conv_std_logic_vector(47232, 16),
49399 => conv_std_logic_vector(47424, 16),
49400 => conv_std_logic_vector(47616, 16),
49401 => conv_std_logic_vector(47808, 16),
49402 => conv_std_logic_vector(48000, 16),
49403 => conv_std_logic_vector(48192, 16),
49404 => conv_std_logic_vector(48384, 16),
49405 => conv_std_logic_vector(48576, 16),
49406 => conv_std_logic_vector(48768, 16),
49407 => conv_std_logic_vector(48960, 16),
49408 => conv_std_logic_vector(0, 16),
49409 => conv_std_logic_vector(193, 16),
49410 => conv_std_logic_vector(386, 16),
49411 => conv_std_logic_vector(579, 16),
49412 => conv_std_logic_vector(772, 16),
49413 => conv_std_logic_vector(965, 16),
49414 => conv_std_logic_vector(1158, 16),
49415 => conv_std_logic_vector(1351, 16),
49416 => conv_std_logic_vector(1544, 16),
49417 => conv_std_logic_vector(1737, 16),
49418 => conv_std_logic_vector(1930, 16),
49419 => conv_std_logic_vector(2123, 16),
49420 => conv_std_logic_vector(2316, 16),
49421 => conv_std_logic_vector(2509, 16),
49422 => conv_std_logic_vector(2702, 16),
49423 => conv_std_logic_vector(2895, 16),
49424 => conv_std_logic_vector(3088, 16),
49425 => conv_std_logic_vector(3281, 16),
49426 => conv_std_logic_vector(3474, 16),
49427 => conv_std_logic_vector(3667, 16),
49428 => conv_std_logic_vector(3860, 16),
49429 => conv_std_logic_vector(4053, 16),
49430 => conv_std_logic_vector(4246, 16),
49431 => conv_std_logic_vector(4439, 16),
49432 => conv_std_logic_vector(4632, 16),
49433 => conv_std_logic_vector(4825, 16),
49434 => conv_std_logic_vector(5018, 16),
49435 => conv_std_logic_vector(5211, 16),
49436 => conv_std_logic_vector(5404, 16),
49437 => conv_std_logic_vector(5597, 16),
49438 => conv_std_logic_vector(5790, 16),
49439 => conv_std_logic_vector(5983, 16),
49440 => conv_std_logic_vector(6176, 16),
49441 => conv_std_logic_vector(6369, 16),
49442 => conv_std_logic_vector(6562, 16),
49443 => conv_std_logic_vector(6755, 16),
49444 => conv_std_logic_vector(6948, 16),
49445 => conv_std_logic_vector(7141, 16),
49446 => conv_std_logic_vector(7334, 16),
49447 => conv_std_logic_vector(7527, 16),
49448 => conv_std_logic_vector(7720, 16),
49449 => conv_std_logic_vector(7913, 16),
49450 => conv_std_logic_vector(8106, 16),
49451 => conv_std_logic_vector(8299, 16),
49452 => conv_std_logic_vector(8492, 16),
49453 => conv_std_logic_vector(8685, 16),
49454 => conv_std_logic_vector(8878, 16),
49455 => conv_std_logic_vector(9071, 16),
49456 => conv_std_logic_vector(9264, 16),
49457 => conv_std_logic_vector(9457, 16),
49458 => conv_std_logic_vector(9650, 16),
49459 => conv_std_logic_vector(9843, 16),
49460 => conv_std_logic_vector(10036, 16),
49461 => conv_std_logic_vector(10229, 16),
49462 => conv_std_logic_vector(10422, 16),
49463 => conv_std_logic_vector(10615, 16),
49464 => conv_std_logic_vector(10808, 16),
49465 => conv_std_logic_vector(11001, 16),
49466 => conv_std_logic_vector(11194, 16),
49467 => conv_std_logic_vector(11387, 16),
49468 => conv_std_logic_vector(11580, 16),
49469 => conv_std_logic_vector(11773, 16),
49470 => conv_std_logic_vector(11966, 16),
49471 => conv_std_logic_vector(12159, 16),
49472 => conv_std_logic_vector(12352, 16),
49473 => conv_std_logic_vector(12545, 16),
49474 => conv_std_logic_vector(12738, 16),
49475 => conv_std_logic_vector(12931, 16),
49476 => conv_std_logic_vector(13124, 16),
49477 => conv_std_logic_vector(13317, 16),
49478 => conv_std_logic_vector(13510, 16),
49479 => conv_std_logic_vector(13703, 16),
49480 => conv_std_logic_vector(13896, 16),
49481 => conv_std_logic_vector(14089, 16),
49482 => conv_std_logic_vector(14282, 16),
49483 => conv_std_logic_vector(14475, 16),
49484 => conv_std_logic_vector(14668, 16),
49485 => conv_std_logic_vector(14861, 16),
49486 => conv_std_logic_vector(15054, 16),
49487 => conv_std_logic_vector(15247, 16),
49488 => conv_std_logic_vector(15440, 16),
49489 => conv_std_logic_vector(15633, 16),
49490 => conv_std_logic_vector(15826, 16),
49491 => conv_std_logic_vector(16019, 16),
49492 => conv_std_logic_vector(16212, 16),
49493 => conv_std_logic_vector(16405, 16),
49494 => conv_std_logic_vector(16598, 16),
49495 => conv_std_logic_vector(16791, 16),
49496 => conv_std_logic_vector(16984, 16),
49497 => conv_std_logic_vector(17177, 16),
49498 => conv_std_logic_vector(17370, 16),
49499 => conv_std_logic_vector(17563, 16),
49500 => conv_std_logic_vector(17756, 16),
49501 => conv_std_logic_vector(17949, 16),
49502 => conv_std_logic_vector(18142, 16),
49503 => conv_std_logic_vector(18335, 16),
49504 => conv_std_logic_vector(18528, 16),
49505 => conv_std_logic_vector(18721, 16),
49506 => conv_std_logic_vector(18914, 16),
49507 => conv_std_logic_vector(19107, 16),
49508 => conv_std_logic_vector(19300, 16),
49509 => conv_std_logic_vector(19493, 16),
49510 => conv_std_logic_vector(19686, 16),
49511 => conv_std_logic_vector(19879, 16),
49512 => conv_std_logic_vector(20072, 16),
49513 => conv_std_logic_vector(20265, 16),
49514 => conv_std_logic_vector(20458, 16),
49515 => conv_std_logic_vector(20651, 16),
49516 => conv_std_logic_vector(20844, 16),
49517 => conv_std_logic_vector(21037, 16),
49518 => conv_std_logic_vector(21230, 16),
49519 => conv_std_logic_vector(21423, 16),
49520 => conv_std_logic_vector(21616, 16),
49521 => conv_std_logic_vector(21809, 16),
49522 => conv_std_logic_vector(22002, 16),
49523 => conv_std_logic_vector(22195, 16),
49524 => conv_std_logic_vector(22388, 16),
49525 => conv_std_logic_vector(22581, 16),
49526 => conv_std_logic_vector(22774, 16),
49527 => conv_std_logic_vector(22967, 16),
49528 => conv_std_logic_vector(23160, 16),
49529 => conv_std_logic_vector(23353, 16),
49530 => conv_std_logic_vector(23546, 16),
49531 => conv_std_logic_vector(23739, 16),
49532 => conv_std_logic_vector(23932, 16),
49533 => conv_std_logic_vector(24125, 16),
49534 => conv_std_logic_vector(24318, 16),
49535 => conv_std_logic_vector(24511, 16),
49536 => conv_std_logic_vector(24704, 16),
49537 => conv_std_logic_vector(24897, 16),
49538 => conv_std_logic_vector(25090, 16),
49539 => conv_std_logic_vector(25283, 16),
49540 => conv_std_logic_vector(25476, 16),
49541 => conv_std_logic_vector(25669, 16),
49542 => conv_std_logic_vector(25862, 16),
49543 => conv_std_logic_vector(26055, 16),
49544 => conv_std_logic_vector(26248, 16),
49545 => conv_std_logic_vector(26441, 16),
49546 => conv_std_logic_vector(26634, 16),
49547 => conv_std_logic_vector(26827, 16),
49548 => conv_std_logic_vector(27020, 16),
49549 => conv_std_logic_vector(27213, 16),
49550 => conv_std_logic_vector(27406, 16),
49551 => conv_std_logic_vector(27599, 16),
49552 => conv_std_logic_vector(27792, 16),
49553 => conv_std_logic_vector(27985, 16),
49554 => conv_std_logic_vector(28178, 16),
49555 => conv_std_logic_vector(28371, 16),
49556 => conv_std_logic_vector(28564, 16),
49557 => conv_std_logic_vector(28757, 16),
49558 => conv_std_logic_vector(28950, 16),
49559 => conv_std_logic_vector(29143, 16),
49560 => conv_std_logic_vector(29336, 16),
49561 => conv_std_logic_vector(29529, 16),
49562 => conv_std_logic_vector(29722, 16),
49563 => conv_std_logic_vector(29915, 16),
49564 => conv_std_logic_vector(30108, 16),
49565 => conv_std_logic_vector(30301, 16),
49566 => conv_std_logic_vector(30494, 16),
49567 => conv_std_logic_vector(30687, 16),
49568 => conv_std_logic_vector(30880, 16),
49569 => conv_std_logic_vector(31073, 16),
49570 => conv_std_logic_vector(31266, 16),
49571 => conv_std_logic_vector(31459, 16),
49572 => conv_std_logic_vector(31652, 16),
49573 => conv_std_logic_vector(31845, 16),
49574 => conv_std_logic_vector(32038, 16),
49575 => conv_std_logic_vector(32231, 16),
49576 => conv_std_logic_vector(32424, 16),
49577 => conv_std_logic_vector(32617, 16),
49578 => conv_std_logic_vector(32810, 16),
49579 => conv_std_logic_vector(33003, 16),
49580 => conv_std_logic_vector(33196, 16),
49581 => conv_std_logic_vector(33389, 16),
49582 => conv_std_logic_vector(33582, 16),
49583 => conv_std_logic_vector(33775, 16),
49584 => conv_std_logic_vector(33968, 16),
49585 => conv_std_logic_vector(34161, 16),
49586 => conv_std_logic_vector(34354, 16),
49587 => conv_std_logic_vector(34547, 16),
49588 => conv_std_logic_vector(34740, 16),
49589 => conv_std_logic_vector(34933, 16),
49590 => conv_std_logic_vector(35126, 16),
49591 => conv_std_logic_vector(35319, 16),
49592 => conv_std_logic_vector(35512, 16),
49593 => conv_std_logic_vector(35705, 16),
49594 => conv_std_logic_vector(35898, 16),
49595 => conv_std_logic_vector(36091, 16),
49596 => conv_std_logic_vector(36284, 16),
49597 => conv_std_logic_vector(36477, 16),
49598 => conv_std_logic_vector(36670, 16),
49599 => conv_std_logic_vector(36863, 16),
49600 => conv_std_logic_vector(37056, 16),
49601 => conv_std_logic_vector(37249, 16),
49602 => conv_std_logic_vector(37442, 16),
49603 => conv_std_logic_vector(37635, 16),
49604 => conv_std_logic_vector(37828, 16),
49605 => conv_std_logic_vector(38021, 16),
49606 => conv_std_logic_vector(38214, 16),
49607 => conv_std_logic_vector(38407, 16),
49608 => conv_std_logic_vector(38600, 16),
49609 => conv_std_logic_vector(38793, 16),
49610 => conv_std_logic_vector(38986, 16),
49611 => conv_std_logic_vector(39179, 16),
49612 => conv_std_logic_vector(39372, 16),
49613 => conv_std_logic_vector(39565, 16),
49614 => conv_std_logic_vector(39758, 16),
49615 => conv_std_logic_vector(39951, 16),
49616 => conv_std_logic_vector(40144, 16),
49617 => conv_std_logic_vector(40337, 16),
49618 => conv_std_logic_vector(40530, 16),
49619 => conv_std_logic_vector(40723, 16),
49620 => conv_std_logic_vector(40916, 16),
49621 => conv_std_logic_vector(41109, 16),
49622 => conv_std_logic_vector(41302, 16),
49623 => conv_std_logic_vector(41495, 16),
49624 => conv_std_logic_vector(41688, 16),
49625 => conv_std_logic_vector(41881, 16),
49626 => conv_std_logic_vector(42074, 16),
49627 => conv_std_logic_vector(42267, 16),
49628 => conv_std_logic_vector(42460, 16),
49629 => conv_std_logic_vector(42653, 16),
49630 => conv_std_logic_vector(42846, 16),
49631 => conv_std_logic_vector(43039, 16),
49632 => conv_std_logic_vector(43232, 16),
49633 => conv_std_logic_vector(43425, 16),
49634 => conv_std_logic_vector(43618, 16),
49635 => conv_std_logic_vector(43811, 16),
49636 => conv_std_logic_vector(44004, 16),
49637 => conv_std_logic_vector(44197, 16),
49638 => conv_std_logic_vector(44390, 16),
49639 => conv_std_logic_vector(44583, 16),
49640 => conv_std_logic_vector(44776, 16),
49641 => conv_std_logic_vector(44969, 16),
49642 => conv_std_logic_vector(45162, 16),
49643 => conv_std_logic_vector(45355, 16),
49644 => conv_std_logic_vector(45548, 16),
49645 => conv_std_logic_vector(45741, 16),
49646 => conv_std_logic_vector(45934, 16),
49647 => conv_std_logic_vector(46127, 16),
49648 => conv_std_logic_vector(46320, 16),
49649 => conv_std_logic_vector(46513, 16),
49650 => conv_std_logic_vector(46706, 16),
49651 => conv_std_logic_vector(46899, 16),
49652 => conv_std_logic_vector(47092, 16),
49653 => conv_std_logic_vector(47285, 16),
49654 => conv_std_logic_vector(47478, 16),
49655 => conv_std_logic_vector(47671, 16),
49656 => conv_std_logic_vector(47864, 16),
49657 => conv_std_logic_vector(48057, 16),
49658 => conv_std_logic_vector(48250, 16),
49659 => conv_std_logic_vector(48443, 16),
49660 => conv_std_logic_vector(48636, 16),
49661 => conv_std_logic_vector(48829, 16),
49662 => conv_std_logic_vector(49022, 16),
49663 => conv_std_logic_vector(49215, 16),
49664 => conv_std_logic_vector(0, 16),
49665 => conv_std_logic_vector(194, 16),
49666 => conv_std_logic_vector(388, 16),
49667 => conv_std_logic_vector(582, 16),
49668 => conv_std_logic_vector(776, 16),
49669 => conv_std_logic_vector(970, 16),
49670 => conv_std_logic_vector(1164, 16),
49671 => conv_std_logic_vector(1358, 16),
49672 => conv_std_logic_vector(1552, 16),
49673 => conv_std_logic_vector(1746, 16),
49674 => conv_std_logic_vector(1940, 16),
49675 => conv_std_logic_vector(2134, 16),
49676 => conv_std_logic_vector(2328, 16),
49677 => conv_std_logic_vector(2522, 16),
49678 => conv_std_logic_vector(2716, 16),
49679 => conv_std_logic_vector(2910, 16),
49680 => conv_std_logic_vector(3104, 16),
49681 => conv_std_logic_vector(3298, 16),
49682 => conv_std_logic_vector(3492, 16),
49683 => conv_std_logic_vector(3686, 16),
49684 => conv_std_logic_vector(3880, 16),
49685 => conv_std_logic_vector(4074, 16),
49686 => conv_std_logic_vector(4268, 16),
49687 => conv_std_logic_vector(4462, 16),
49688 => conv_std_logic_vector(4656, 16),
49689 => conv_std_logic_vector(4850, 16),
49690 => conv_std_logic_vector(5044, 16),
49691 => conv_std_logic_vector(5238, 16),
49692 => conv_std_logic_vector(5432, 16),
49693 => conv_std_logic_vector(5626, 16),
49694 => conv_std_logic_vector(5820, 16),
49695 => conv_std_logic_vector(6014, 16),
49696 => conv_std_logic_vector(6208, 16),
49697 => conv_std_logic_vector(6402, 16),
49698 => conv_std_logic_vector(6596, 16),
49699 => conv_std_logic_vector(6790, 16),
49700 => conv_std_logic_vector(6984, 16),
49701 => conv_std_logic_vector(7178, 16),
49702 => conv_std_logic_vector(7372, 16),
49703 => conv_std_logic_vector(7566, 16),
49704 => conv_std_logic_vector(7760, 16),
49705 => conv_std_logic_vector(7954, 16),
49706 => conv_std_logic_vector(8148, 16),
49707 => conv_std_logic_vector(8342, 16),
49708 => conv_std_logic_vector(8536, 16),
49709 => conv_std_logic_vector(8730, 16),
49710 => conv_std_logic_vector(8924, 16),
49711 => conv_std_logic_vector(9118, 16),
49712 => conv_std_logic_vector(9312, 16),
49713 => conv_std_logic_vector(9506, 16),
49714 => conv_std_logic_vector(9700, 16),
49715 => conv_std_logic_vector(9894, 16),
49716 => conv_std_logic_vector(10088, 16),
49717 => conv_std_logic_vector(10282, 16),
49718 => conv_std_logic_vector(10476, 16),
49719 => conv_std_logic_vector(10670, 16),
49720 => conv_std_logic_vector(10864, 16),
49721 => conv_std_logic_vector(11058, 16),
49722 => conv_std_logic_vector(11252, 16),
49723 => conv_std_logic_vector(11446, 16),
49724 => conv_std_logic_vector(11640, 16),
49725 => conv_std_logic_vector(11834, 16),
49726 => conv_std_logic_vector(12028, 16),
49727 => conv_std_logic_vector(12222, 16),
49728 => conv_std_logic_vector(12416, 16),
49729 => conv_std_logic_vector(12610, 16),
49730 => conv_std_logic_vector(12804, 16),
49731 => conv_std_logic_vector(12998, 16),
49732 => conv_std_logic_vector(13192, 16),
49733 => conv_std_logic_vector(13386, 16),
49734 => conv_std_logic_vector(13580, 16),
49735 => conv_std_logic_vector(13774, 16),
49736 => conv_std_logic_vector(13968, 16),
49737 => conv_std_logic_vector(14162, 16),
49738 => conv_std_logic_vector(14356, 16),
49739 => conv_std_logic_vector(14550, 16),
49740 => conv_std_logic_vector(14744, 16),
49741 => conv_std_logic_vector(14938, 16),
49742 => conv_std_logic_vector(15132, 16),
49743 => conv_std_logic_vector(15326, 16),
49744 => conv_std_logic_vector(15520, 16),
49745 => conv_std_logic_vector(15714, 16),
49746 => conv_std_logic_vector(15908, 16),
49747 => conv_std_logic_vector(16102, 16),
49748 => conv_std_logic_vector(16296, 16),
49749 => conv_std_logic_vector(16490, 16),
49750 => conv_std_logic_vector(16684, 16),
49751 => conv_std_logic_vector(16878, 16),
49752 => conv_std_logic_vector(17072, 16),
49753 => conv_std_logic_vector(17266, 16),
49754 => conv_std_logic_vector(17460, 16),
49755 => conv_std_logic_vector(17654, 16),
49756 => conv_std_logic_vector(17848, 16),
49757 => conv_std_logic_vector(18042, 16),
49758 => conv_std_logic_vector(18236, 16),
49759 => conv_std_logic_vector(18430, 16),
49760 => conv_std_logic_vector(18624, 16),
49761 => conv_std_logic_vector(18818, 16),
49762 => conv_std_logic_vector(19012, 16),
49763 => conv_std_logic_vector(19206, 16),
49764 => conv_std_logic_vector(19400, 16),
49765 => conv_std_logic_vector(19594, 16),
49766 => conv_std_logic_vector(19788, 16),
49767 => conv_std_logic_vector(19982, 16),
49768 => conv_std_logic_vector(20176, 16),
49769 => conv_std_logic_vector(20370, 16),
49770 => conv_std_logic_vector(20564, 16),
49771 => conv_std_logic_vector(20758, 16),
49772 => conv_std_logic_vector(20952, 16),
49773 => conv_std_logic_vector(21146, 16),
49774 => conv_std_logic_vector(21340, 16),
49775 => conv_std_logic_vector(21534, 16),
49776 => conv_std_logic_vector(21728, 16),
49777 => conv_std_logic_vector(21922, 16),
49778 => conv_std_logic_vector(22116, 16),
49779 => conv_std_logic_vector(22310, 16),
49780 => conv_std_logic_vector(22504, 16),
49781 => conv_std_logic_vector(22698, 16),
49782 => conv_std_logic_vector(22892, 16),
49783 => conv_std_logic_vector(23086, 16),
49784 => conv_std_logic_vector(23280, 16),
49785 => conv_std_logic_vector(23474, 16),
49786 => conv_std_logic_vector(23668, 16),
49787 => conv_std_logic_vector(23862, 16),
49788 => conv_std_logic_vector(24056, 16),
49789 => conv_std_logic_vector(24250, 16),
49790 => conv_std_logic_vector(24444, 16),
49791 => conv_std_logic_vector(24638, 16),
49792 => conv_std_logic_vector(24832, 16),
49793 => conv_std_logic_vector(25026, 16),
49794 => conv_std_logic_vector(25220, 16),
49795 => conv_std_logic_vector(25414, 16),
49796 => conv_std_logic_vector(25608, 16),
49797 => conv_std_logic_vector(25802, 16),
49798 => conv_std_logic_vector(25996, 16),
49799 => conv_std_logic_vector(26190, 16),
49800 => conv_std_logic_vector(26384, 16),
49801 => conv_std_logic_vector(26578, 16),
49802 => conv_std_logic_vector(26772, 16),
49803 => conv_std_logic_vector(26966, 16),
49804 => conv_std_logic_vector(27160, 16),
49805 => conv_std_logic_vector(27354, 16),
49806 => conv_std_logic_vector(27548, 16),
49807 => conv_std_logic_vector(27742, 16),
49808 => conv_std_logic_vector(27936, 16),
49809 => conv_std_logic_vector(28130, 16),
49810 => conv_std_logic_vector(28324, 16),
49811 => conv_std_logic_vector(28518, 16),
49812 => conv_std_logic_vector(28712, 16),
49813 => conv_std_logic_vector(28906, 16),
49814 => conv_std_logic_vector(29100, 16),
49815 => conv_std_logic_vector(29294, 16),
49816 => conv_std_logic_vector(29488, 16),
49817 => conv_std_logic_vector(29682, 16),
49818 => conv_std_logic_vector(29876, 16),
49819 => conv_std_logic_vector(30070, 16),
49820 => conv_std_logic_vector(30264, 16),
49821 => conv_std_logic_vector(30458, 16),
49822 => conv_std_logic_vector(30652, 16),
49823 => conv_std_logic_vector(30846, 16),
49824 => conv_std_logic_vector(31040, 16),
49825 => conv_std_logic_vector(31234, 16),
49826 => conv_std_logic_vector(31428, 16),
49827 => conv_std_logic_vector(31622, 16),
49828 => conv_std_logic_vector(31816, 16),
49829 => conv_std_logic_vector(32010, 16),
49830 => conv_std_logic_vector(32204, 16),
49831 => conv_std_logic_vector(32398, 16),
49832 => conv_std_logic_vector(32592, 16),
49833 => conv_std_logic_vector(32786, 16),
49834 => conv_std_logic_vector(32980, 16),
49835 => conv_std_logic_vector(33174, 16),
49836 => conv_std_logic_vector(33368, 16),
49837 => conv_std_logic_vector(33562, 16),
49838 => conv_std_logic_vector(33756, 16),
49839 => conv_std_logic_vector(33950, 16),
49840 => conv_std_logic_vector(34144, 16),
49841 => conv_std_logic_vector(34338, 16),
49842 => conv_std_logic_vector(34532, 16),
49843 => conv_std_logic_vector(34726, 16),
49844 => conv_std_logic_vector(34920, 16),
49845 => conv_std_logic_vector(35114, 16),
49846 => conv_std_logic_vector(35308, 16),
49847 => conv_std_logic_vector(35502, 16),
49848 => conv_std_logic_vector(35696, 16),
49849 => conv_std_logic_vector(35890, 16),
49850 => conv_std_logic_vector(36084, 16),
49851 => conv_std_logic_vector(36278, 16),
49852 => conv_std_logic_vector(36472, 16),
49853 => conv_std_logic_vector(36666, 16),
49854 => conv_std_logic_vector(36860, 16),
49855 => conv_std_logic_vector(37054, 16),
49856 => conv_std_logic_vector(37248, 16),
49857 => conv_std_logic_vector(37442, 16),
49858 => conv_std_logic_vector(37636, 16),
49859 => conv_std_logic_vector(37830, 16),
49860 => conv_std_logic_vector(38024, 16),
49861 => conv_std_logic_vector(38218, 16),
49862 => conv_std_logic_vector(38412, 16),
49863 => conv_std_logic_vector(38606, 16),
49864 => conv_std_logic_vector(38800, 16),
49865 => conv_std_logic_vector(38994, 16),
49866 => conv_std_logic_vector(39188, 16),
49867 => conv_std_logic_vector(39382, 16),
49868 => conv_std_logic_vector(39576, 16),
49869 => conv_std_logic_vector(39770, 16),
49870 => conv_std_logic_vector(39964, 16),
49871 => conv_std_logic_vector(40158, 16),
49872 => conv_std_logic_vector(40352, 16),
49873 => conv_std_logic_vector(40546, 16),
49874 => conv_std_logic_vector(40740, 16),
49875 => conv_std_logic_vector(40934, 16),
49876 => conv_std_logic_vector(41128, 16),
49877 => conv_std_logic_vector(41322, 16),
49878 => conv_std_logic_vector(41516, 16),
49879 => conv_std_logic_vector(41710, 16),
49880 => conv_std_logic_vector(41904, 16),
49881 => conv_std_logic_vector(42098, 16),
49882 => conv_std_logic_vector(42292, 16),
49883 => conv_std_logic_vector(42486, 16),
49884 => conv_std_logic_vector(42680, 16),
49885 => conv_std_logic_vector(42874, 16),
49886 => conv_std_logic_vector(43068, 16),
49887 => conv_std_logic_vector(43262, 16),
49888 => conv_std_logic_vector(43456, 16),
49889 => conv_std_logic_vector(43650, 16),
49890 => conv_std_logic_vector(43844, 16),
49891 => conv_std_logic_vector(44038, 16),
49892 => conv_std_logic_vector(44232, 16),
49893 => conv_std_logic_vector(44426, 16),
49894 => conv_std_logic_vector(44620, 16),
49895 => conv_std_logic_vector(44814, 16),
49896 => conv_std_logic_vector(45008, 16),
49897 => conv_std_logic_vector(45202, 16),
49898 => conv_std_logic_vector(45396, 16),
49899 => conv_std_logic_vector(45590, 16),
49900 => conv_std_logic_vector(45784, 16),
49901 => conv_std_logic_vector(45978, 16),
49902 => conv_std_logic_vector(46172, 16),
49903 => conv_std_logic_vector(46366, 16),
49904 => conv_std_logic_vector(46560, 16),
49905 => conv_std_logic_vector(46754, 16),
49906 => conv_std_logic_vector(46948, 16),
49907 => conv_std_logic_vector(47142, 16),
49908 => conv_std_logic_vector(47336, 16),
49909 => conv_std_logic_vector(47530, 16),
49910 => conv_std_logic_vector(47724, 16),
49911 => conv_std_logic_vector(47918, 16),
49912 => conv_std_logic_vector(48112, 16),
49913 => conv_std_logic_vector(48306, 16),
49914 => conv_std_logic_vector(48500, 16),
49915 => conv_std_logic_vector(48694, 16),
49916 => conv_std_logic_vector(48888, 16),
49917 => conv_std_logic_vector(49082, 16),
49918 => conv_std_logic_vector(49276, 16),
49919 => conv_std_logic_vector(49470, 16),
49920 => conv_std_logic_vector(0, 16),
49921 => conv_std_logic_vector(195, 16),
49922 => conv_std_logic_vector(390, 16),
49923 => conv_std_logic_vector(585, 16),
49924 => conv_std_logic_vector(780, 16),
49925 => conv_std_logic_vector(975, 16),
49926 => conv_std_logic_vector(1170, 16),
49927 => conv_std_logic_vector(1365, 16),
49928 => conv_std_logic_vector(1560, 16),
49929 => conv_std_logic_vector(1755, 16),
49930 => conv_std_logic_vector(1950, 16),
49931 => conv_std_logic_vector(2145, 16),
49932 => conv_std_logic_vector(2340, 16),
49933 => conv_std_logic_vector(2535, 16),
49934 => conv_std_logic_vector(2730, 16),
49935 => conv_std_logic_vector(2925, 16),
49936 => conv_std_logic_vector(3120, 16),
49937 => conv_std_logic_vector(3315, 16),
49938 => conv_std_logic_vector(3510, 16),
49939 => conv_std_logic_vector(3705, 16),
49940 => conv_std_logic_vector(3900, 16),
49941 => conv_std_logic_vector(4095, 16),
49942 => conv_std_logic_vector(4290, 16),
49943 => conv_std_logic_vector(4485, 16),
49944 => conv_std_logic_vector(4680, 16),
49945 => conv_std_logic_vector(4875, 16),
49946 => conv_std_logic_vector(5070, 16),
49947 => conv_std_logic_vector(5265, 16),
49948 => conv_std_logic_vector(5460, 16),
49949 => conv_std_logic_vector(5655, 16),
49950 => conv_std_logic_vector(5850, 16),
49951 => conv_std_logic_vector(6045, 16),
49952 => conv_std_logic_vector(6240, 16),
49953 => conv_std_logic_vector(6435, 16),
49954 => conv_std_logic_vector(6630, 16),
49955 => conv_std_logic_vector(6825, 16),
49956 => conv_std_logic_vector(7020, 16),
49957 => conv_std_logic_vector(7215, 16),
49958 => conv_std_logic_vector(7410, 16),
49959 => conv_std_logic_vector(7605, 16),
49960 => conv_std_logic_vector(7800, 16),
49961 => conv_std_logic_vector(7995, 16),
49962 => conv_std_logic_vector(8190, 16),
49963 => conv_std_logic_vector(8385, 16),
49964 => conv_std_logic_vector(8580, 16),
49965 => conv_std_logic_vector(8775, 16),
49966 => conv_std_logic_vector(8970, 16),
49967 => conv_std_logic_vector(9165, 16),
49968 => conv_std_logic_vector(9360, 16),
49969 => conv_std_logic_vector(9555, 16),
49970 => conv_std_logic_vector(9750, 16),
49971 => conv_std_logic_vector(9945, 16),
49972 => conv_std_logic_vector(10140, 16),
49973 => conv_std_logic_vector(10335, 16),
49974 => conv_std_logic_vector(10530, 16),
49975 => conv_std_logic_vector(10725, 16),
49976 => conv_std_logic_vector(10920, 16),
49977 => conv_std_logic_vector(11115, 16),
49978 => conv_std_logic_vector(11310, 16),
49979 => conv_std_logic_vector(11505, 16),
49980 => conv_std_logic_vector(11700, 16),
49981 => conv_std_logic_vector(11895, 16),
49982 => conv_std_logic_vector(12090, 16),
49983 => conv_std_logic_vector(12285, 16),
49984 => conv_std_logic_vector(12480, 16),
49985 => conv_std_logic_vector(12675, 16),
49986 => conv_std_logic_vector(12870, 16),
49987 => conv_std_logic_vector(13065, 16),
49988 => conv_std_logic_vector(13260, 16),
49989 => conv_std_logic_vector(13455, 16),
49990 => conv_std_logic_vector(13650, 16),
49991 => conv_std_logic_vector(13845, 16),
49992 => conv_std_logic_vector(14040, 16),
49993 => conv_std_logic_vector(14235, 16),
49994 => conv_std_logic_vector(14430, 16),
49995 => conv_std_logic_vector(14625, 16),
49996 => conv_std_logic_vector(14820, 16),
49997 => conv_std_logic_vector(15015, 16),
49998 => conv_std_logic_vector(15210, 16),
49999 => conv_std_logic_vector(15405, 16),
50000 => conv_std_logic_vector(15600, 16),
50001 => conv_std_logic_vector(15795, 16),
50002 => conv_std_logic_vector(15990, 16),
50003 => conv_std_logic_vector(16185, 16),
50004 => conv_std_logic_vector(16380, 16),
50005 => conv_std_logic_vector(16575, 16),
50006 => conv_std_logic_vector(16770, 16),
50007 => conv_std_logic_vector(16965, 16),
50008 => conv_std_logic_vector(17160, 16),
50009 => conv_std_logic_vector(17355, 16),
50010 => conv_std_logic_vector(17550, 16),
50011 => conv_std_logic_vector(17745, 16),
50012 => conv_std_logic_vector(17940, 16),
50013 => conv_std_logic_vector(18135, 16),
50014 => conv_std_logic_vector(18330, 16),
50015 => conv_std_logic_vector(18525, 16),
50016 => conv_std_logic_vector(18720, 16),
50017 => conv_std_logic_vector(18915, 16),
50018 => conv_std_logic_vector(19110, 16),
50019 => conv_std_logic_vector(19305, 16),
50020 => conv_std_logic_vector(19500, 16),
50021 => conv_std_logic_vector(19695, 16),
50022 => conv_std_logic_vector(19890, 16),
50023 => conv_std_logic_vector(20085, 16),
50024 => conv_std_logic_vector(20280, 16),
50025 => conv_std_logic_vector(20475, 16),
50026 => conv_std_logic_vector(20670, 16),
50027 => conv_std_logic_vector(20865, 16),
50028 => conv_std_logic_vector(21060, 16),
50029 => conv_std_logic_vector(21255, 16),
50030 => conv_std_logic_vector(21450, 16),
50031 => conv_std_logic_vector(21645, 16),
50032 => conv_std_logic_vector(21840, 16),
50033 => conv_std_logic_vector(22035, 16),
50034 => conv_std_logic_vector(22230, 16),
50035 => conv_std_logic_vector(22425, 16),
50036 => conv_std_logic_vector(22620, 16),
50037 => conv_std_logic_vector(22815, 16),
50038 => conv_std_logic_vector(23010, 16),
50039 => conv_std_logic_vector(23205, 16),
50040 => conv_std_logic_vector(23400, 16),
50041 => conv_std_logic_vector(23595, 16),
50042 => conv_std_logic_vector(23790, 16),
50043 => conv_std_logic_vector(23985, 16),
50044 => conv_std_logic_vector(24180, 16),
50045 => conv_std_logic_vector(24375, 16),
50046 => conv_std_logic_vector(24570, 16),
50047 => conv_std_logic_vector(24765, 16),
50048 => conv_std_logic_vector(24960, 16),
50049 => conv_std_logic_vector(25155, 16),
50050 => conv_std_logic_vector(25350, 16),
50051 => conv_std_logic_vector(25545, 16),
50052 => conv_std_logic_vector(25740, 16),
50053 => conv_std_logic_vector(25935, 16),
50054 => conv_std_logic_vector(26130, 16),
50055 => conv_std_logic_vector(26325, 16),
50056 => conv_std_logic_vector(26520, 16),
50057 => conv_std_logic_vector(26715, 16),
50058 => conv_std_logic_vector(26910, 16),
50059 => conv_std_logic_vector(27105, 16),
50060 => conv_std_logic_vector(27300, 16),
50061 => conv_std_logic_vector(27495, 16),
50062 => conv_std_logic_vector(27690, 16),
50063 => conv_std_logic_vector(27885, 16),
50064 => conv_std_logic_vector(28080, 16),
50065 => conv_std_logic_vector(28275, 16),
50066 => conv_std_logic_vector(28470, 16),
50067 => conv_std_logic_vector(28665, 16),
50068 => conv_std_logic_vector(28860, 16),
50069 => conv_std_logic_vector(29055, 16),
50070 => conv_std_logic_vector(29250, 16),
50071 => conv_std_logic_vector(29445, 16),
50072 => conv_std_logic_vector(29640, 16),
50073 => conv_std_logic_vector(29835, 16),
50074 => conv_std_logic_vector(30030, 16),
50075 => conv_std_logic_vector(30225, 16),
50076 => conv_std_logic_vector(30420, 16),
50077 => conv_std_logic_vector(30615, 16),
50078 => conv_std_logic_vector(30810, 16),
50079 => conv_std_logic_vector(31005, 16),
50080 => conv_std_logic_vector(31200, 16),
50081 => conv_std_logic_vector(31395, 16),
50082 => conv_std_logic_vector(31590, 16),
50083 => conv_std_logic_vector(31785, 16),
50084 => conv_std_logic_vector(31980, 16),
50085 => conv_std_logic_vector(32175, 16),
50086 => conv_std_logic_vector(32370, 16),
50087 => conv_std_logic_vector(32565, 16),
50088 => conv_std_logic_vector(32760, 16),
50089 => conv_std_logic_vector(32955, 16),
50090 => conv_std_logic_vector(33150, 16),
50091 => conv_std_logic_vector(33345, 16),
50092 => conv_std_logic_vector(33540, 16),
50093 => conv_std_logic_vector(33735, 16),
50094 => conv_std_logic_vector(33930, 16),
50095 => conv_std_logic_vector(34125, 16),
50096 => conv_std_logic_vector(34320, 16),
50097 => conv_std_logic_vector(34515, 16),
50098 => conv_std_logic_vector(34710, 16),
50099 => conv_std_logic_vector(34905, 16),
50100 => conv_std_logic_vector(35100, 16),
50101 => conv_std_logic_vector(35295, 16),
50102 => conv_std_logic_vector(35490, 16),
50103 => conv_std_logic_vector(35685, 16),
50104 => conv_std_logic_vector(35880, 16),
50105 => conv_std_logic_vector(36075, 16),
50106 => conv_std_logic_vector(36270, 16),
50107 => conv_std_logic_vector(36465, 16),
50108 => conv_std_logic_vector(36660, 16),
50109 => conv_std_logic_vector(36855, 16),
50110 => conv_std_logic_vector(37050, 16),
50111 => conv_std_logic_vector(37245, 16),
50112 => conv_std_logic_vector(37440, 16),
50113 => conv_std_logic_vector(37635, 16),
50114 => conv_std_logic_vector(37830, 16),
50115 => conv_std_logic_vector(38025, 16),
50116 => conv_std_logic_vector(38220, 16),
50117 => conv_std_logic_vector(38415, 16),
50118 => conv_std_logic_vector(38610, 16),
50119 => conv_std_logic_vector(38805, 16),
50120 => conv_std_logic_vector(39000, 16),
50121 => conv_std_logic_vector(39195, 16),
50122 => conv_std_logic_vector(39390, 16),
50123 => conv_std_logic_vector(39585, 16),
50124 => conv_std_logic_vector(39780, 16),
50125 => conv_std_logic_vector(39975, 16),
50126 => conv_std_logic_vector(40170, 16),
50127 => conv_std_logic_vector(40365, 16),
50128 => conv_std_logic_vector(40560, 16),
50129 => conv_std_logic_vector(40755, 16),
50130 => conv_std_logic_vector(40950, 16),
50131 => conv_std_logic_vector(41145, 16),
50132 => conv_std_logic_vector(41340, 16),
50133 => conv_std_logic_vector(41535, 16),
50134 => conv_std_logic_vector(41730, 16),
50135 => conv_std_logic_vector(41925, 16),
50136 => conv_std_logic_vector(42120, 16),
50137 => conv_std_logic_vector(42315, 16),
50138 => conv_std_logic_vector(42510, 16),
50139 => conv_std_logic_vector(42705, 16),
50140 => conv_std_logic_vector(42900, 16),
50141 => conv_std_logic_vector(43095, 16),
50142 => conv_std_logic_vector(43290, 16),
50143 => conv_std_logic_vector(43485, 16),
50144 => conv_std_logic_vector(43680, 16),
50145 => conv_std_logic_vector(43875, 16),
50146 => conv_std_logic_vector(44070, 16),
50147 => conv_std_logic_vector(44265, 16),
50148 => conv_std_logic_vector(44460, 16),
50149 => conv_std_logic_vector(44655, 16),
50150 => conv_std_logic_vector(44850, 16),
50151 => conv_std_logic_vector(45045, 16),
50152 => conv_std_logic_vector(45240, 16),
50153 => conv_std_logic_vector(45435, 16),
50154 => conv_std_logic_vector(45630, 16),
50155 => conv_std_logic_vector(45825, 16),
50156 => conv_std_logic_vector(46020, 16),
50157 => conv_std_logic_vector(46215, 16),
50158 => conv_std_logic_vector(46410, 16),
50159 => conv_std_logic_vector(46605, 16),
50160 => conv_std_logic_vector(46800, 16),
50161 => conv_std_logic_vector(46995, 16),
50162 => conv_std_logic_vector(47190, 16),
50163 => conv_std_logic_vector(47385, 16),
50164 => conv_std_logic_vector(47580, 16),
50165 => conv_std_logic_vector(47775, 16),
50166 => conv_std_logic_vector(47970, 16),
50167 => conv_std_logic_vector(48165, 16),
50168 => conv_std_logic_vector(48360, 16),
50169 => conv_std_logic_vector(48555, 16),
50170 => conv_std_logic_vector(48750, 16),
50171 => conv_std_logic_vector(48945, 16),
50172 => conv_std_logic_vector(49140, 16),
50173 => conv_std_logic_vector(49335, 16),
50174 => conv_std_logic_vector(49530, 16),
50175 => conv_std_logic_vector(49725, 16),
50176 => conv_std_logic_vector(0, 16),
50177 => conv_std_logic_vector(196, 16),
50178 => conv_std_logic_vector(392, 16),
50179 => conv_std_logic_vector(588, 16),
50180 => conv_std_logic_vector(784, 16),
50181 => conv_std_logic_vector(980, 16),
50182 => conv_std_logic_vector(1176, 16),
50183 => conv_std_logic_vector(1372, 16),
50184 => conv_std_logic_vector(1568, 16),
50185 => conv_std_logic_vector(1764, 16),
50186 => conv_std_logic_vector(1960, 16),
50187 => conv_std_logic_vector(2156, 16),
50188 => conv_std_logic_vector(2352, 16),
50189 => conv_std_logic_vector(2548, 16),
50190 => conv_std_logic_vector(2744, 16),
50191 => conv_std_logic_vector(2940, 16),
50192 => conv_std_logic_vector(3136, 16),
50193 => conv_std_logic_vector(3332, 16),
50194 => conv_std_logic_vector(3528, 16),
50195 => conv_std_logic_vector(3724, 16),
50196 => conv_std_logic_vector(3920, 16),
50197 => conv_std_logic_vector(4116, 16),
50198 => conv_std_logic_vector(4312, 16),
50199 => conv_std_logic_vector(4508, 16),
50200 => conv_std_logic_vector(4704, 16),
50201 => conv_std_logic_vector(4900, 16),
50202 => conv_std_logic_vector(5096, 16),
50203 => conv_std_logic_vector(5292, 16),
50204 => conv_std_logic_vector(5488, 16),
50205 => conv_std_logic_vector(5684, 16),
50206 => conv_std_logic_vector(5880, 16),
50207 => conv_std_logic_vector(6076, 16),
50208 => conv_std_logic_vector(6272, 16),
50209 => conv_std_logic_vector(6468, 16),
50210 => conv_std_logic_vector(6664, 16),
50211 => conv_std_logic_vector(6860, 16),
50212 => conv_std_logic_vector(7056, 16),
50213 => conv_std_logic_vector(7252, 16),
50214 => conv_std_logic_vector(7448, 16),
50215 => conv_std_logic_vector(7644, 16),
50216 => conv_std_logic_vector(7840, 16),
50217 => conv_std_logic_vector(8036, 16),
50218 => conv_std_logic_vector(8232, 16),
50219 => conv_std_logic_vector(8428, 16),
50220 => conv_std_logic_vector(8624, 16),
50221 => conv_std_logic_vector(8820, 16),
50222 => conv_std_logic_vector(9016, 16),
50223 => conv_std_logic_vector(9212, 16),
50224 => conv_std_logic_vector(9408, 16),
50225 => conv_std_logic_vector(9604, 16),
50226 => conv_std_logic_vector(9800, 16),
50227 => conv_std_logic_vector(9996, 16),
50228 => conv_std_logic_vector(10192, 16),
50229 => conv_std_logic_vector(10388, 16),
50230 => conv_std_logic_vector(10584, 16),
50231 => conv_std_logic_vector(10780, 16),
50232 => conv_std_logic_vector(10976, 16),
50233 => conv_std_logic_vector(11172, 16),
50234 => conv_std_logic_vector(11368, 16),
50235 => conv_std_logic_vector(11564, 16),
50236 => conv_std_logic_vector(11760, 16),
50237 => conv_std_logic_vector(11956, 16),
50238 => conv_std_logic_vector(12152, 16),
50239 => conv_std_logic_vector(12348, 16),
50240 => conv_std_logic_vector(12544, 16),
50241 => conv_std_logic_vector(12740, 16),
50242 => conv_std_logic_vector(12936, 16),
50243 => conv_std_logic_vector(13132, 16),
50244 => conv_std_logic_vector(13328, 16),
50245 => conv_std_logic_vector(13524, 16),
50246 => conv_std_logic_vector(13720, 16),
50247 => conv_std_logic_vector(13916, 16),
50248 => conv_std_logic_vector(14112, 16),
50249 => conv_std_logic_vector(14308, 16),
50250 => conv_std_logic_vector(14504, 16),
50251 => conv_std_logic_vector(14700, 16),
50252 => conv_std_logic_vector(14896, 16),
50253 => conv_std_logic_vector(15092, 16),
50254 => conv_std_logic_vector(15288, 16),
50255 => conv_std_logic_vector(15484, 16),
50256 => conv_std_logic_vector(15680, 16),
50257 => conv_std_logic_vector(15876, 16),
50258 => conv_std_logic_vector(16072, 16),
50259 => conv_std_logic_vector(16268, 16),
50260 => conv_std_logic_vector(16464, 16),
50261 => conv_std_logic_vector(16660, 16),
50262 => conv_std_logic_vector(16856, 16),
50263 => conv_std_logic_vector(17052, 16),
50264 => conv_std_logic_vector(17248, 16),
50265 => conv_std_logic_vector(17444, 16),
50266 => conv_std_logic_vector(17640, 16),
50267 => conv_std_logic_vector(17836, 16),
50268 => conv_std_logic_vector(18032, 16),
50269 => conv_std_logic_vector(18228, 16),
50270 => conv_std_logic_vector(18424, 16),
50271 => conv_std_logic_vector(18620, 16),
50272 => conv_std_logic_vector(18816, 16),
50273 => conv_std_logic_vector(19012, 16),
50274 => conv_std_logic_vector(19208, 16),
50275 => conv_std_logic_vector(19404, 16),
50276 => conv_std_logic_vector(19600, 16),
50277 => conv_std_logic_vector(19796, 16),
50278 => conv_std_logic_vector(19992, 16),
50279 => conv_std_logic_vector(20188, 16),
50280 => conv_std_logic_vector(20384, 16),
50281 => conv_std_logic_vector(20580, 16),
50282 => conv_std_logic_vector(20776, 16),
50283 => conv_std_logic_vector(20972, 16),
50284 => conv_std_logic_vector(21168, 16),
50285 => conv_std_logic_vector(21364, 16),
50286 => conv_std_logic_vector(21560, 16),
50287 => conv_std_logic_vector(21756, 16),
50288 => conv_std_logic_vector(21952, 16),
50289 => conv_std_logic_vector(22148, 16),
50290 => conv_std_logic_vector(22344, 16),
50291 => conv_std_logic_vector(22540, 16),
50292 => conv_std_logic_vector(22736, 16),
50293 => conv_std_logic_vector(22932, 16),
50294 => conv_std_logic_vector(23128, 16),
50295 => conv_std_logic_vector(23324, 16),
50296 => conv_std_logic_vector(23520, 16),
50297 => conv_std_logic_vector(23716, 16),
50298 => conv_std_logic_vector(23912, 16),
50299 => conv_std_logic_vector(24108, 16),
50300 => conv_std_logic_vector(24304, 16),
50301 => conv_std_logic_vector(24500, 16),
50302 => conv_std_logic_vector(24696, 16),
50303 => conv_std_logic_vector(24892, 16),
50304 => conv_std_logic_vector(25088, 16),
50305 => conv_std_logic_vector(25284, 16),
50306 => conv_std_logic_vector(25480, 16),
50307 => conv_std_logic_vector(25676, 16),
50308 => conv_std_logic_vector(25872, 16),
50309 => conv_std_logic_vector(26068, 16),
50310 => conv_std_logic_vector(26264, 16),
50311 => conv_std_logic_vector(26460, 16),
50312 => conv_std_logic_vector(26656, 16),
50313 => conv_std_logic_vector(26852, 16),
50314 => conv_std_logic_vector(27048, 16),
50315 => conv_std_logic_vector(27244, 16),
50316 => conv_std_logic_vector(27440, 16),
50317 => conv_std_logic_vector(27636, 16),
50318 => conv_std_logic_vector(27832, 16),
50319 => conv_std_logic_vector(28028, 16),
50320 => conv_std_logic_vector(28224, 16),
50321 => conv_std_logic_vector(28420, 16),
50322 => conv_std_logic_vector(28616, 16),
50323 => conv_std_logic_vector(28812, 16),
50324 => conv_std_logic_vector(29008, 16),
50325 => conv_std_logic_vector(29204, 16),
50326 => conv_std_logic_vector(29400, 16),
50327 => conv_std_logic_vector(29596, 16),
50328 => conv_std_logic_vector(29792, 16),
50329 => conv_std_logic_vector(29988, 16),
50330 => conv_std_logic_vector(30184, 16),
50331 => conv_std_logic_vector(30380, 16),
50332 => conv_std_logic_vector(30576, 16),
50333 => conv_std_logic_vector(30772, 16),
50334 => conv_std_logic_vector(30968, 16),
50335 => conv_std_logic_vector(31164, 16),
50336 => conv_std_logic_vector(31360, 16),
50337 => conv_std_logic_vector(31556, 16),
50338 => conv_std_logic_vector(31752, 16),
50339 => conv_std_logic_vector(31948, 16),
50340 => conv_std_logic_vector(32144, 16),
50341 => conv_std_logic_vector(32340, 16),
50342 => conv_std_logic_vector(32536, 16),
50343 => conv_std_logic_vector(32732, 16),
50344 => conv_std_logic_vector(32928, 16),
50345 => conv_std_logic_vector(33124, 16),
50346 => conv_std_logic_vector(33320, 16),
50347 => conv_std_logic_vector(33516, 16),
50348 => conv_std_logic_vector(33712, 16),
50349 => conv_std_logic_vector(33908, 16),
50350 => conv_std_logic_vector(34104, 16),
50351 => conv_std_logic_vector(34300, 16),
50352 => conv_std_logic_vector(34496, 16),
50353 => conv_std_logic_vector(34692, 16),
50354 => conv_std_logic_vector(34888, 16),
50355 => conv_std_logic_vector(35084, 16),
50356 => conv_std_logic_vector(35280, 16),
50357 => conv_std_logic_vector(35476, 16),
50358 => conv_std_logic_vector(35672, 16),
50359 => conv_std_logic_vector(35868, 16),
50360 => conv_std_logic_vector(36064, 16),
50361 => conv_std_logic_vector(36260, 16),
50362 => conv_std_logic_vector(36456, 16),
50363 => conv_std_logic_vector(36652, 16),
50364 => conv_std_logic_vector(36848, 16),
50365 => conv_std_logic_vector(37044, 16),
50366 => conv_std_logic_vector(37240, 16),
50367 => conv_std_logic_vector(37436, 16),
50368 => conv_std_logic_vector(37632, 16),
50369 => conv_std_logic_vector(37828, 16),
50370 => conv_std_logic_vector(38024, 16),
50371 => conv_std_logic_vector(38220, 16),
50372 => conv_std_logic_vector(38416, 16),
50373 => conv_std_logic_vector(38612, 16),
50374 => conv_std_logic_vector(38808, 16),
50375 => conv_std_logic_vector(39004, 16),
50376 => conv_std_logic_vector(39200, 16),
50377 => conv_std_logic_vector(39396, 16),
50378 => conv_std_logic_vector(39592, 16),
50379 => conv_std_logic_vector(39788, 16),
50380 => conv_std_logic_vector(39984, 16),
50381 => conv_std_logic_vector(40180, 16),
50382 => conv_std_logic_vector(40376, 16),
50383 => conv_std_logic_vector(40572, 16),
50384 => conv_std_logic_vector(40768, 16),
50385 => conv_std_logic_vector(40964, 16),
50386 => conv_std_logic_vector(41160, 16),
50387 => conv_std_logic_vector(41356, 16),
50388 => conv_std_logic_vector(41552, 16),
50389 => conv_std_logic_vector(41748, 16),
50390 => conv_std_logic_vector(41944, 16),
50391 => conv_std_logic_vector(42140, 16),
50392 => conv_std_logic_vector(42336, 16),
50393 => conv_std_logic_vector(42532, 16),
50394 => conv_std_logic_vector(42728, 16),
50395 => conv_std_logic_vector(42924, 16),
50396 => conv_std_logic_vector(43120, 16),
50397 => conv_std_logic_vector(43316, 16),
50398 => conv_std_logic_vector(43512, 16),
50399 => conv_std_logic_vector(43708, 16),
50400 => conv_std_logic_vector(43904, 16),
50401 => conv_std_logic_vector(44100, 16),
50402 => conv_std_logic_vector(44296, 16),
50403 => conv_std_logic_vector(44492, 16),
50404 => conv_std_logic_vector(44688, 16),
50405 => conv_std_logic_vector(44884, 16),
50406 => conv_std_logic_vector(45080, 16),
50407 => conv_std_logic_vector(45276, 16),
50408 => conv_std_logic_vector(45472, 16),
50409 => conv_std_logic_vector(45668, 16),
50410 => conv_std_logic_vector(45864, 16),
50411 => conv_std_logic_vector(46060, 16),
50412 => conv_std_logic_vector(46256, 16),
50413 => conv_std_logic_vector(46452, 16),
50414 => conv_std_logic_vector(46648, 16),
50415 => conv_std_logic_vector(46844, 16),
50416 => conv_std_logic_vector(47040, 16),
50417 => conv_std_logic_vector(47236, 16),
50418 => conv_std_logic_vector(47432, 16),
50419 => conv_std_logic_vector(47628, 16),
50420 => conv_std_logic_vector(47824, 16),
50421 => conv_std_logic_vector(48020, 16),
50422 => conv_std_logic_vector(48216, 16),
50423 => conv_std_logic_vector(48412, 16),
50424 => conv_std_logic_vector(48608, 16),
50425 => conv_std_logic_vector(48804, 16),
50426 => conv_std_logic_vector(49000, 16),
50427 => conv_std_logic_vector(49196, 16),
50428 => conv_std_logic_vector(49392, 16),
50429 => conv_std_logic_vector(49588, 16),
50430 => conv_std_logic_vector(49784, 16),
50431 => conv_std_logic_vector(49980, 16),
50432 => conv_std_logic_vector(0, 16),
50433 => conv_std_logic_vector(197, 16),
50434 => conv_std_logic_vector(394, 16),
50435 => conv_std_logic_vector(591, 16),
50436 => conv_std_logic_vector(788, 16),
50437 => conv_std_logic_vector(985, 16),
50438 => conv_std_logic_vector(1182, 16),
50439 => conv_std_logic_vector(1379, 16),
50440 => conv_std_logic_vector(1576, 16),
50441 => conv_std_logic_vector(1773, 16),
50442 => conv_std_logic_vector(1970, 16),
50443 => conv_std_logic_vector(2167, 16),
50444 => conv_std_logic_vector(2364, 16),
50445 => conv_std_logic_vector(2561, 16),
50446 => conv_std_logic_vector(2758, 16),
50447 => conv_std_logic_vector(2955, 16),
50448 => conv_std_logic_vector(3152, 16),
50449 => conv_std_logic_vector(3349, 16),
50450 => conv_std_logic_vector(3546, 16),
50451 => conv_std_logic_vector(3743, 16),
50452 => conv_std_logic_vector(3940, 16),
50453 => conv_std_logic_vector(4137, 16),
50454 => conv_std_logic_vector(4334, 16),
50455 => conv_std_logic_vector(4531, 16),
50456 => conv_std_logic_vector(4728, 16),
50457 => conv_std_logic_vector(4925, 16),
50458 => conv_std_logic_vector(5122, 16),
50459 => conv_std_logic_vector(5319, 16),
50460 => conv_std_logic_vector(5516, 16),
50461 => conv_std_logic_vector(5713, 16),
50462 => conv_std_logic_vector(5910, 16),
50463 => conv_std_logic_vector(6107, 16),
50464 => conv_std_logic_vector(6304, 16),
50465 => conv_std_logic_vector(6501, 16),
50466 => conv_std_logic_vector(6698, 16),
50467 => conv_std_logic_vector(6895, 16),
50468 => conv_std_logic_vector(7092, 16),
50469 => conv_std_logic_vector(7289, 16),
50470 => conv_std_logic_vector(7486, 16),
50471 => conv_std_logic_vector(7683, 16),
50472 => conv_std_logic_vector(7880, 16),
50473 => conv_std_logic_vector(8077, 16),
50474 => conv_std_logic_vector(8274, 16),
50475 => conv_std_logic_vector(8471, 16),
50476 => conv_std_logic_vector(8668, 16),
50477 => conv_std_logic_vector(8865, 16),
50478 => conv_std_logic_vector(9062, 16),
50479 => conv_std_logic_vector(9259, 16),
50480 => conv_std_logic_vector(9456, 16),
50481 => conv_std_logic_vector(9653, 16),
50482 => conv_std_logic_vector(9850, 16),
50483 => conv_std_logic_vector(10047, 16),
50484 => conv_std_logic_vector(10244, 16),
50485 => conv_std_logic_vector(10441, 16),
50486 => conv_std_logic_vector(10638, 16),
50487 => conv_std_logic_vector(10835, 16),
50488 => conv_std_logic_vector(11032, 16),
50489 => conv_std_logic_vector(11229, 16),
50490 => conv_std_logic_vector(11426, 16),
50491 => conv_std_logic_vector(11623, 16),
50492 => conv_std_logic_vector(11820, 16),
50493 => conv_std_logic_vector(12017, 16),
50494 => conv_std_logic_vector(12214, 16),
50495 => conv_std_logic_vector(12411, 16),
50496 => conv_std_logic_vector(12608, 16),
50497 => conv_std_logic_vector(12805, 16),
50498 => conv_std_logic_vector(13002, 16),
50499 => conv_std_logic_vector(13199, 16),
50500 => conv_std_logic_vector(13396, 16),
50501 => conv_std_logic_vector(13593, 16),
50502 => conv_std_logic_vector(13790, 16),
50503 => conv_std_logic_vector(13987, 16),
50504 => conv_std_logic_vector(14184, 16),
50505 => conv_std_logic_vector(14381, 16),
50506 => conv_std_logic_vector(14578, 16),
50507 => conv_std_logic_vector(14775, 16),
50508 => conv_std_logic_vector(14972, 16),
50509 => conv_std_logic_vector(15169, 16),
50510 => conv_std_logic_vector(15366, 16),
50511 => conv_std_logic_vector(15563, 16),
50512 => conv_std_logic_vector(15760, 16),
50513 => conv_std_logic_vector(15957, 16),
50514 => conv_std_logic_vector(16154, 16),
50515 => conv_std_logic_vector(16351, 16),
50516 => conv_std_logic_vector(16548, 16),
50517 => conv_std_logic_vector(16745, 16),
50518 => conv_std_logic_vector(16942, 16),
50519 => conv_std_logic_vector(17139, 16),
50520 => conv_std_logic_vector(17336, 16),
50521 => conv_std_logic_vector(17533, 16),
50522 => conv_std_logic_vector(17730, 16),
50523 => conv_std_logic_vector(17927, 16),
50524 => conv_std_logic_vector(18124, 16),
50525 => conv_std_logic_vector(18321, 16),
50526 => conv_std_logic_vector(18518, 16),
50527 => conv_std_logic_vector(18715, 16),
50528 => conv_std_logic_vector(18912, 16),
50529 => conv_std_logic_vector(19109, 16),
50530 => conv_std_logic_vector(19306, 16),
50531 => conv_std_logic_vector(19503, 16),
50532 => conv_std_logic_vector(19700, 16),
50533 => conv_std_logic_vector(19897, 16),
50534 => conv_std_logic_vector(20094, 16),
50535 => conv_std_logic_vector(20291, 16),
50536 => conv_std_logic_vector(20488, 16),
50537 => conv_std_logic_vector(20685, 16),
50538 => conv_std_logic_vector(20882, 16),
50539 => conv_std_logic_vector(21079, 16),
50540 => conv_std_logic_vector(21276, 16),
50541 => conv_std_logic_vector(21473, 16),
50542 => conv_std_logic_vector(21670, 16),
50543 => conv_std_logic_vector(21867, 16),
50544 => conv_std_logic_vector(22064, 16),
50545 => conv_std_logic_vector(22261, 16),
50546 => conv_std_logic_vector(22458, 16),
50547 => conv_std_logic_vector(22655, 16),
50548 => conv_std_logic_vector(22852, 16),
50549 => conv_std_logic_vector(23049, 16),
50550 => conv_std_logic_vector(23246, 16),
50551 => conv_std_logic_vector(23443, 16),
50552 => conv_std_logic_vector(23640, 16),
50553 => conv_std_logic_vector(23837, 16),
50554 => conv_std_logic_vector(24034, 16),
50555 => conv_std_logic_vector(24231, 16),
50556 => conv_std_logic_vector(24428, 16),
50557 => conv_std_logic_vector(24625, 16),
50558 => conv_std_logic_vector(24822, 16),
50559 => conv_std_logic_vector(25019, 16),
50560 => conv_std_logic_vector(25216, 16),
50561 => conv_std_logic_vector(25413, 16),
50562 => conv_std_logic_vector(25610, 16),
50563 => conv_std_logic_vector(25807, 16),
50564 => conv_std_logic_vector(26004, 16),
50565 => conv_std_logic_vector(26201, 16),
50566 => conv_std_logic_vector(26398, 16),
50567 => conv_std_logic_vector(26595, 16),
50568 => conv_std_logic_vector(26792, 16),
50569 => conv_std_logic_vector(26989, 16),
50570 => conv_std_logic_vector(27186, 16),
50571 => conv_std_logic_vector(27383, 16),
50572 => conv_std_logic_vector(27580, 16),
50573 => conv_std_logic_vector(27777, 16),
50574 => conv_std_logic_vector(27974, 16),
50575 => conv_std_logic_vector(28171, 16),
50576 => conv_std_logic_vector(28368, 16),
50577 => conv_std_logic_vector(28565, 16),
50578 => conv_std_logic_vector(28762, 16),
50579 => conv_std_logic_vector(28959, 16),
50580 => conv_std_logic_vector(29156, 16),
50581 => conv_std_logic_vector(29353, 16),
50582 => conv_std_logic_vector(29550, 16),
50583 => conv_std_logic_vector(29747, 16),
50584 => conv_std_logic_vector(29944, 16),
50585 => conv_std_logic_vector(30141, 16),
50586 => conv_std_logic_vector(30338, 16),
50587 => conv_std_logic_vector(30535, 16),
50588 => conv_std_logic_vector(30732, 16),
50589 => conv_std_logic_vector(30929, 16),
50590 => conv_std_logic_vector(31126, 16),
50591 => conv_std_logic_vector(31323, 16),
50592 => conv_std_logic_vector(31520, 16),
50593 => conv_std_logic_vector(31717, 16),
50594 => conv_std_logic_vector(31914, 16),
50595 => conv_std_logic_vector(32111, 16),
50596 => conv_std_logic_vector(32308, 16),
50597 => conv_std_logic_vector(32505, 16),
50598 => conv_std_logic_vector(32702, 16),
50599 => conv_std_logic_vector(32899, 16),
50600 => conv_std_logic_vector(33096, 16),
50601 => conv_std_logic_vector(33293, 16),
50602 => conv_std_logic_vector(33490, 16),
50603 => conv_std_logic_vector(33687, 16),
50604 => conv_std_logic_vector(33884, 16),
50605 => conv_std_logic_vector(34081, 16),
50606 => conv_std_logic_vector(34278, 16),
50607 => conv_std_logic_vector(34475, 16),
50608 => conv_std_logic_vector(34672, 16),
50609 => conv_std_logic_vector(34869, 16),
50610 => conv_std_logic_vector(35066, 16),
50611 => conv_std_logic_vector(35263, 16),
50612 => conv_std_logic_vector(35460, 16),
50613 => conv_std_logic_vector(35657, 16),
50614 => conv_std_logic_vector(35854, 16),
50615 => conv_std_logic_vector(36051, 16),
50616 => conv_std_logic_vector(36248, 16),
50617 => conv_std_logic_vector(36445, 16),
50618 => conv_std_logic_vector(36642, 16),
50619 => conv_std_logic_vector(36839, 16),
50620 => conv_std_logic_vector(37036, 16),
50621 => conv_std_logic_vector(37233, 16),
50622 => conv_std_logic_vector(37430, 16),
50623 => conv_std_logic_vector(37627, 16),
50624 => conv_std_logic_vector(37824, 16),
50625 => conv_std_logic_vector(38021, 16),
50626 => conv_std_logic_vector(38218, 16),
50627 => conv_std_logic_vector(38415, 16),
50628 => conv_std_logic_vector(38612, 16),
50629 => conv_std_logic_vector(38809, 16),
50630 => conv_std_logic_vector(39006, 16),
50631 => conv_std_logic_vector(39203, 16),
50632 => conv_std_logic_vector(39400, 16),
50633 => conv_std_logic_vector(39597, 16),
50634 => conv_std_logic_vector(39794, 16),
50635 => conv_std_logic_vector(39991, 16),
50636 => conv_std_logic_vector(40188, 16),
50637 => conv_std_logic_vector(40385, 16),
50638 => conv_std_logic_vector(40582, 16),
50639 => conv_std_logic_vector(40779, 16),
50640 => conv_std_logic_vector(40976, 16),
50641 => conv_std_logic_vector(41173, 16),
50642 => conv_std_logic_vector(41370, 16),
50643 => conv_std_logic_vector(41567, 16),
50644 => conv_std_logic_vector(41764, 16),
50645 => conv_std_logic_vector(41961, 16),
50646 => conv_std_logic_vector(42158, 16),
50647 => conv_std_logic_vector(42355, 16),
50648 => conv_std_logic_vector(42552, 16),
50649 => conv_std_logic_vector(42749, 16),
50650 => conv_std_logic_vector(42946, 16),
50651 => conv_std_logic_vector(43143, 16),
50652 => conv_std_logic_vector(43340, 16),
50653 => conv_std_logic_vector(43537, 16),
50654 => conv_std_logic_vector(43734, 16),
50655 => conv_std_logic_vector(43931, 16),
50656 => conv_std_logic_vector(44128, 16),
50657 => conv_std_logic_vector(44325, 16),
50658 => conv_std_logic_vector(44522, 16),
50659 => conv_std_logic_vector(44719, 16),
50660 => conv_std_logic_vector(44916, 16),
50661 => conv_std_logic_vector(45113, 16),
50662 => conv_std_logic_vector(45310, 16),
50663 => conv_std_logic_vector(45507, 16),
50664 => conv_std_logic_vector(45704, 16),
50665 => conv_std_logic_vector(45901, 16),
50666 => conv_std_logic_vector(46098, 16),
50667 => conv_std_logic_vector(46295, 16),
50668 => conv_std_logic_vector(46492, 16),
50669 => conv_std_logic_vector(46689, 16),
50670 => conv_std_logic_vector(46886, 16),
50671 => conv_std_logic_vector(47083, 16),
50672 => conv_std_logic_vector(47280, 16),
50673 => conv_std_logic_vector(47477, 16),
50674 => conv_std_logic_vector(47674, 16),
50675 => conv_std_logic_vector(47871, 16),
50676 => conv_std_logic_vector(48068, 16),
50677 => conv_std_logic_vector(48265, 16),
50678 => conv_std_logic_vector(48462, 16),
50679 => conv_std_logic_vector(48659, 16),
50680 => conv_std_logic_vector(48856, 16),
50681 => conv_std_logic_vector(49053, 16),
50682 => conv_std_logic_vector(49250, 16),
50683 => conv_std_logic_vector(49447, 16),
50684 => conv_std_logic_vector(49644, 16),
50685 => conv_std_logic_vector(49841, 16),
50686 => conv_std_logic_vector(50038, 16),
50687 => conv_std_logic_vector(50235, 16),
50688 => conv_std_logic_vector(0, 16),
50689 => conv_std_logic_vector(198, 16),
50690 => conv_std_logic_vector(396, 16),
50691 => conv_std_logic_vector(594, 16),
50692 => conv_std_logic_vector(792, 16),
50693 => conv_std_logic_vector(990, 16),
50694 => conv_std_logic_vector(1188, 16),
50695 => conv_std_logic_vector(1386, 16),
50696 => conv_std_logic_vector(1584, 16),
50697 => conv_std_logic_vector(1782, 16),
50698 => conv_std_logic_vector(1980, 16),
50699 => conv_std_logic_vector(2178, 16),
50700 => conv_std_logic_vector(2376, 16),
50701 => conv_std_logic_vector(2574, 16),
50702 => conv_std_logic_vector(2772, 16),
50703 => conv_std_logic_vector(2970, 16),
50704 => conv_std_logic_vector(3168, 16),
50705 => conv_std_logic_vector(3366, 16),
50706 => conv_std_logic_vector(3564, 16),
50707 => conv_std_logic_vector(3762, 16),
50708 => conv_std_logic_vector(3960, 16),
50709 => conv_std_logic_vector(4158, 16),
50710 => conv_std_logic_vector(4356, 16),
50711 => conv_std_logic_vector(4554, 16),
50712 => conv_std_logic_vector(4752, 16),
50713 => conv_std_logic_vector(4950, 16),
50714 => conv_std_logic_vector(5148, 16),
50715 => conv_std_logic_vector(5346, 16),
50716 => conv_std_logic_vector(5544, 16),
50717 => conv_std_logic_vector(5742, 16),
50718 => conv_std_logic_vector(5940, 16),
50719 => conv_std_logic_vector(6138, 16),
50720 => conv_std_logic_vector(6336, 16),
50721 => conv_std_logic_vector(6534, 16),
50722 => conv_std_logic_vector(6732, 16),
50723 => conv_std_logic_vector(6930, 16),
50724 => conv_std_logic_vector(7128, 16),
50725 => conv_std_logic_vector(7326, 16),
50726 => conv_std_logic_vector(7524, 16),
50727 => conv_std_logic_vector(7722, 16),
50728 => conv_std_logic_vector(7920, 16),
50729 => conv_std_logic_vector(8118, 16),
50730 => conv_std_logic_vector(8316, 16),
50731 => conv_std_logic_vector(8514, 16),
50732 => conv_std_logic_vector(8712, 16),
50733 => conv_std_logic_vector(8910, 16),
50734 => conv_std_logic_vector(9108, 16),
50735 => conv_std_logic_vector(9306, 16),
50736 => conv_std_logic_vector(9504, 16),
50737 => conv_std_logic_vector(9702, 16),
50738 => conv_std_logic_vector(9900, 16),
50739 => conv_std_logic_vector(10098, 16),
50740 => conv_std_logic_vector(10296, 16),
50741 => conv_std_logic_vector(10494, 16),
50742 => conv_std_logic_vector(10692, 16),
50743 => conv_std_logic_vector(10890, 16),
50744 => conv_std_logic_vector(11088, 16),
50745 => conv_std_logic_vector(11286, 16),
50746 => conv_std_logic_vector(11484, 16),
50747 => conv_std_logic_vector(11682, 16),
50748 => conv_std_logic_vector(11880, 16),
50749 => conv_std_logic_vector(12078, 16),
50750 => conv_std_logic_vector(12276, 16),
50751 => conv_std_logic_vector(12474, 16),
50752 => conv_std_logic_vector(12672, 16),
50753 => conv_std_logic_vector(12870, 16),
50754 => conv_std_logic_vector(13068, 16),
50755 => conv_std_logic_vector(13266, 16),
50756 => conv_std_logic_vector(13464, 16),
50757 => conv_std_logic_vector(13662, 16),
50758 => conv_std_logic_vector(13860, 16),
50759 => conv_std_logic_vector(14058, 16),
50760 => conv_std_logic_vector(14256, 16),
50761 => conv_std_logic_vector(14454, 16),
50762 => conv_std_logic_vector(14652, 16),
50763 => conv_std_logic_vector(14850, 16),
50764 => conv_std_logic_vector(15048, 16),
50765 => conv_std_logic_vector(15246, 16),
50766 => conv_std_logic_vector(15444, 16),
50767 => conv_std_logic_vector(15642, 16),
50768 => conv_std_logic_vector(15840, 16),
50769 => conv_std_logic_vector(16038, 16),
50770 => conv_std_logic_vector(16236, 16),
50771 => conv_std_logic_vector(16434, 16),
50772 => conv_std_logic_vector(16632, 16),
50773 => conv_std_logic_vector(16830, 16),
50774 => conv_std_logic_vector(17028, 16),
50775 => conv_std_logic_vector(17226, 16),
50776 => conv_std_logic_vector(17424, 16),
50777 => conv_std_logic_vector(17622, 16),
50778 => conv_std_logic_vector(17820, 16),
50779 => conv_std_logic_vector(18018, 16),
50780 => conv_std_logic_vector(18216, 16),
50781 => conv_std_logic_vector(18414, 16),
50782 => conv_std_logic_vector(18612, 16),
50783 => conv_std_logic_vector(18810, 16),
50784 => conv_std_logic_vector(19008, 16),
50785 => conv_std_logic_vector(19206, 16),
50786 => conv_std_logic_vector(19404, 16),
50787 => conv_std_logic_vector(19602, 16),
50788 => conv_std_logic_vector(19800, 16),
50789 => conv_std_logic_vector(19998, 16),
50790 => conv_std_logic_vector(20196, 16),
50791 => conv_std_logic_vector(20394, 16),
50792 => conv_std_logic_vector(20592, 16),
50793 => conv_std_logic_vector(20790, 16),
50794 => conv_std_logic_vector(20988, 16),
50795 => conv_std_logic_vector(21186, 16),
50796 => conv_std_logic_vector(21384, 16),
50797 => conv_std_logic_vector(21582, 16),
50798 => conv_std_logic_vector(21780, 16),
50799 => conv_std_logic_vector(21978, 16),
50800 => conv_std_logic_vector(22176, 16),
50801 => conv_std_logic_vector(22374, 16),
50802 => conv_std_logic_vector(22572, 16),
50803 => conv_std_logic_vector(22770, 16),
50804 => conv_std_logic_vector(22968, 16),
50805 => conv_std_logic_vector(23166, 16),
50806 => conv_std_logic_vector(23364, 16),
50807 => conv_std_logic_vector(23562, 16),
50808 => conv_std_logic_vector(23760, 16),
50809 => conv_std_logic_vector(23958, 16),
50810 => conv_std_logic_vector(24156, 16),
50811 => conv_std_logic_vector(24354, 16),
50812 => conv_std_logic_vector(24552, 16),
50813 => conv_std_logic_vector(24750, 16),
50814 => conv_std_logic_vector(24948, 16),
50815 => conv_std_logic_vector(25146, 16),
50816 => conv_std_logic_vector(25344, 16),
50817 => conv_std_logic_vector(25542, 16),
50818 => conv_std_logic_vector(25740, 16),
50819 => conv_std_logic_vector(25938, 16),
50820 => conv_std_logic_vector(26136, 16),
50821 => conv_std_logic_vector(26334, 16),
50822 => conv_std_logic_vector(26532, 16),
50823 => conv_std_logic_vector(26730, 16),
50824 => conv_std_logic_vector(26928, 16),
50825 => conv_std_logic_vector(27126, 16),
50826 => conv_std_logic_vector(27324, 16),
50827 => conv_std_logic_vector(27522, 16),
50828 => conv_std_logic_vector(27720, 16),
50829 => conv_std_logic_vector(27918, 16),
50830 => conv_std_logic_vector(28116, 16),
50831 => conv_std_logic_vector(28314, 16),
50832 => conv_std_logic_vector(28512, 16),
50833 => conv_std_logic_vector(28710, 16),
50834 => conv_std_logic_vector(28908, 16),
50835 => conv_std_logic_vector(29106, 16),
50836 => conv_std_logic_vector(29304, 16),
50837 => conv_std_logic_vector(29502, 16),
50838 => conv_std_logic_vector(29700, 16),
50839 => conv_std_logic_vector(29898, 16),
50840 => conv_std_logic_vector(30096, 16),
50841 => conv_std_logic_vector(30294, 16),
50842 => conv_std_logic_vector(30492, 16),
50843 => conv_std_logic_vector(30690, 16),
50844 => conv_std_logic_vector(30888, 16),
50845 => conv_std_logic_vector(31086, 16),
50846 => conv_std_logic_vector(31284, 16),
50847 => conv_std_logic_vector(31482, 16),
50848 => conv_std_logic_vector(31680, 16),
50849 => conv_std_logic_vector(31878, 16),
50850 => conv_std_logic_vector(32076, 16),
50851 => conv_std_logic_vector(32274, 16),
50852 => conv_std_logic_vector(32472, 16),
50853 => conv_std_logic_vector(32670, 16),
50854 => conv_std_logic_vector(32868, 16),
50855 => conv_std_logic_vector(33066, 16),
50856 => conv_std_logic_vector(33264, 16),
50857 => conv_std_logic_vector(33462, 16),
50858 => conv_std_logic_vector(33660, 16),
50859 => conv_std_logic_vector(33858, 16),
50860 => conv_std_logic_vector(34056, 16),
50861 => conv_std_logic_vector(34254, 16),
50862 => conv_std_logic_vector(34452, 16),
50863 => conv_std_logic_vector(34650, 16),
50864 => conv_std_logic_vector(34848, 16),
50865 => conv_std_logic_vector(35046, 16),
50866 => conv_std_logic_vector(35244, 16),
50867 => conv_std_logic_vector(35442, 16),
50868 => conv_std_logic_vector(35640, 16),
50869 => conv_std_logic_vector(35838, 16),
50870 => conv_std_logic_vector(36036, 16),
50871 => conv_std_logic_vector(36234, 16),
50872 => conv_std_logic_vector(36432, 16),
50873 => conv_std_logic_vector(36630, 16),
50874 => conv_std_logic_vector(36828, 16),
50875 => conv_std_logic_vector(37026, 16),
50876 => conv_std_logic_vector(37224, 16),
50877 => conv_std_logic_vector(37422, 16),
50878 => conv_std_logic_vector(37620, 16),
50879 => conv_std_logic_vector(37818, 16),
50880 => conv_std_logic_vector(38016, 16),
50881 => conv_std_logic_vector(38214, 16),
50882 => conv_std_logic_vector(38412, 16),
50883 => conv_std_logic_vector(38610, 16),
50884 => conv_std_logic_vector(38808, 16),
50885 => conv_std_logic_vector(39006, 16),
50886 => conv_std_logic_vector(39204, 16),
50887 => conv_std_logic_vector(39402, 16),
50888 => conv_std_logic_vector(39600, 16),
50889 => conv_std_logic_vector(39798, 16),
50890 => conv_std_logic_vector(39996, 16),
50891 => conv_std_logic_vector(40194, 16),
50892 => conv_std_logic_vector(40392, 16),
50893 => conv_std_logic_vector(40590, 16),
50894 => conv_std_logic_vector(40788, 16),
50895 => conv_std_logic_vector(40986, 16),
50896 => conv_std_logic_vector(41184, 16),
50897 => conv_std_logic_vector(41382, 16),
50898 => conv_std_logic_vector(41580, 16),
50899 => conv_std_logic_vector(41778, 16),
50900 => conv_std_logic_vector(41976, 16),
50901 => conv_std_logic_vector(42174, 16),
50902 => conv_std_logic_vector(42372, 16),
50903 => conv_std_logic_vector(42570, 16),
50904 => conv_std_logic_vector(42768, 16),
50905 => conv_std_logic_vector(42966, 16),
50906 => conv_std_logic_vector(43164, 16),
50907 => conv_std_logic_vector(43362, 16),
50908 => conv_std_logic_vector(43560, 16),
50909 => conv_std_logic_vector(43758, 16),
50910 => conv_std_logic_vector(43956, 16),
50911 => conv_std_logic_vector(44154, 16),
50912 => conv_std_logic_vector(44352, 16),
50913 => conv_std_logic_vector(44550, 16),
50914 => conv_std_logic_vector(44748, 16),
50915 => conv_std_logic_vector(44946, 16),
50916 => conv_std_logic_vector(45144, 16),
50917 => conv_std_logic_vector(45342, 16),
50918 => conv_std_logic_vector(45540, 16),
50919 => conv_std_logic_vector(45738, 16),
50920 => conv_std_logic_vector(45936, 16),
50921 => conv_std_logic_vector(46134, 16),
50922 => conv_std_logic_vector(46332, 16),
50923 => conv_std_logic_vector(46530, 16),
50924 => conv_std_logic_vector(46728, 16),
50925 => conv_std_logic_vector(46926, 16),
50926 => conv_std_logic_vector(47124, 16),
50927 => conv_std_logic_vector(47322, 16),
50928 => conv_std_logic_vector(47520, 16),
50929 => conv_std_logic_vector(47718, 16),
50930 => conv_std_logic_vector(47916, 16),
50931 => conv_std_logic_vector(48114, 16),
50932 => conv_std_logic_vector(48312, 16),
50933 => conv_std_logic_vector(48510, 16),
50934 => conv_std_logic_vector(48708, 16),
50935 => conv_std_logic_vector(48906, 16),
50936 => conv_std_logic_vector(49104, 16),
50937 => conv_std_logic_vector(49302, 16),
50938 => conv_std_logic_vector(49500, 16),
50939 => conv_std_logic_vector(49698, 16),
50940 => conv_std_logic_vector(49896, 16),
50941 => conv_std_logic_vector(50094, 16),
50942 => conv_std_logic_vector(50292, 16),
50943 => conv_std_logic_vector(50490, 16),
50944 => conv_std_logic_vector(0, 16),
50945 => conv_std_logic_vector(199, 16),
50946 => conv_std_logic_vector(398, 16),
50947 => conv_std_logic_vector(597, 16),
50948 => conv_std_logic_vector(796, 16),
50949 => conv_std_logic_vector(995, 16),
50950 => conv_std_logic_vector(1194, 16),
50951 => conv_std_logic_vector(1393, 16),
50952 => conv_std_logic_vector(1592, 16),
50953 => conv_std_logic_vector(1791, 16),
50954 => conv_std_logic_vector(1990, 16),
50955 => conv_std_logic_vector(2189, 16),
50956 => conv_std_logic_vector(2388, 16),
50957 => conv_std_logic_vector(2587, 16),
50958 => conv_std_logic_vector(2786, 16),
50959 => conv_std_logic_vector(2985, 16),
50960 => conv_std_logic_vector(3184, 16),
50961 => conv_std_logic_vector(3383, 16),
50962 => conv_std_logic_vector(3582, 16),
50963 => conv_std_logic_vector(3781, 16),
50964 => conv_std_logic_vector(3980, 16),
50965 => conv_std_logic_vector(4179, 16),
50966 => conv_std_logic_vector(4378, 16),
50967 => conv_std_logic_vector(4577, 16),
50968 => conv_std_logic_vector(4776, 16),
50969 => conv_std_logic_vector(4975, 16),
50970 => conv_std_logic_vector(5174, 16),
50971 => conv_std_logic_vector(5373, 16),
50972 => conv_std_logic_vector(5572, 16),
50973 => conv_std_logic_vector(5771, 16),
50974 => conv_std_logic_vector(5970, 16),
50975 => conv_std_logic_vector(6169, 16),
50976 => conv_std_logic_vector(6368, 16),
50977 => conv_std_logic_vector(6567, 16),
50978 => conv_std_logic_vector(6766, 16),
50979 => conv_std_logic_vector(6965, 16),
50980 => conv_std_logic_vector(7164, 16),
50981 => conv_std_logic_vector(7363, 16),
50982 => conv_std_logic_vector(7562, 16),
50983 => conv_std_logic_vector(7761, 16),
50984 => conv_std_logic_vector(7960, 16),
50985 => conv_std_logic_vector(8159, 16),
50986 => conv_std_logic_vector(8358, 16),
50987 => conv_std_logic_vector(8557, 16),
50988 => conv_std_logic_vector(8756, 16),
50989 => conv_std_logic_vector(8955, 16),
50990 => conv_std_logic_vector(9154, 16),
50991 => conv_std_logic_vector(9353, 16),
50992 => conv_std_logic_vector(9552, 16),
50993 => conv_std_logic_vector(9751, 16),
50994 => conv_std_logic_vector(9950, 16),
50995 => conv_std_logic_vector(10149, 16),
50996 => conv_std_logic_vector(10348, 16),
50997 => conv_std_logic_vector(10547, 16),
50998 => conv_std_logic_vector(10746, 16),
50999 => conv_std_logic_vector(10945, 16),
51000 => conv_std_logic_vector(11144, 16),
51001 => conv_std_logic_vector(11343, 16),
51002 => conv_std_logic_vector(11542, 16),
51003 => conv_std_logic_vector(11741, 16),
51004 => conv_std_logic_vector(11940, 16),
51005 => conv_std_logic_vector(12139, 16),
51006 => conv_std_logic_vector(12338, 16),
51007 => conv_std_logic_vector(12537, 16),
51008 => conv_std_logic_vector(12736, 16),
51009 => conv_std_logic_vector(12935, 16),
51010 => conv_std_logic_vector(13134, 16),
51011 => conv_std_logic_vector(13333, 16),
51012 => conv_std_logic_vector(13532, 16),
51013 => conv_std_logic_vector(13731, 16),
51014 => conv_std_logic_vector(13930, 16),
51015 => conv_std_logic_vector(14129, 16),
51016 => conv_std_logic_vector(14328, 16),
51017 => conv_std_logic_vector(14527, 16),
51018 => conv_std_logic_vector(14726, 16),
51019 => conv_std_logic_vector(14925, 16),
51020 => conv_std_logic_vector(15124, 16),
51021 => conv_std_logic_vector(15323, 16),
51022 => conv_std_logic_vector(15522, 16),
51023 => conv_std_logic_vector(15721, 16),
51024 => conv_std_logic_vector(15920, 16),
51025 => conv_std_logic_vector(16119, 16),
51026 => conv_std_logic_vector(16318, 16),
51027 => conv_std_logic_vector(16517, 16),
51028 => conv_std_logic_vector(16716, 16),
51029 => conv_std_logic_vector(16915, 16),
51030 => conv_std_logic_vector(17114, 16),
51031 => conv_std_logic_vector(17313, 16),
51032 => conv_std_logic_vector(17512, 16),
51033 => conv_std_logic_vector(17711, 16),
51034 => conv_std_logic_vector(17910, 16),
51035 => conv_std_logic_vector(18109, 16),
51036 => conv_std_logic_vector(18308, 16),
51037 => conv_std_logic_vector(18507, 16),
51038 => conv_std_logic_vector(18706, 16),
51039 => conv_std_logic_vector(18905, 16),
51040 => conv_std_logic_vector(19104, 16),
51041 => conv_std_logic_vector(19303, 16),
51042 => conv_std_logic_vector(19502, 16),
51043 => conv_std_logic_vector(19701, 16),
51044 => conv_std_logic_vector(19900, 16),
51045 => conv_std_logic_vector(20099, 16),
51046 => conv_std_logic_vector(20298, 16),
51047 => conv_std_logic_vector(20497, 16),
51048 => conv_std_logic_vector(20696, 16),
51049 => conv_std_logic_vector(20895, 16),
51050 => conv_std_logic_vector(21094, 16),
51051 => conv_std_logic_vector(21293, 16),
51052 => conv_std_logic_vector(21492, 16),
51053 => conv_std_logic_vector(21691, 16),
51054 => conv_std_logic_vector(21890, 16),
51055 => conv_std_logic_vector(22089, 16),
51056 => conv_std_logic_vector(22288, 16),
51057 => conv_std_logic_vector(22487, 16),
51058 => conv_std_logic_vector(22686, 16),
51059 => conv_std_logic_vector(22885, 16),
51060 => conv_std_logic_vector(23084, 16),
51061 => conv_std_logic_vector(23283, 16),
51062 => conv_std_logic_vector(23482, 16),
51063 => conv_std_logic_vector(23681, 16),
51064 => conv_std_logic_vector(23880, 16),
51065 => conv_std_logic_vector(24079, 16),
51066 => conv_std_logic_vector(24278, 16),
51067 => conv_std_logic_vector(24477, 16),
51068 => conv_std_logic_vector(24676, 16),
51069 => conv_std_logic_vector(24875, 16),
51070 => conv_std_logic_vector(25074, 16),
51071 => conv_std_logic_vector(25273, 16),
51072 => conv_std_logic_vector(25472, 16),
51073 => conv_std_logic_vector(25671, 16),
51074 => conv_std_logic_vector(25870, 16),
51075 => conv_std_logic_vector(26069, 16),
51076 => conv_std_logic_vector(26268, 16),
51077 => conv_std_logic_vector(26467, 16),
51078 => conv_std_logic_vector(26666, 16),
51079 => conv_std_logic_vector(26865, 16),
51080 => conv_std_logic_vector(27064, 16),
51081 => conv_std_logic_vector(27263, 16),
51082 => conv_std_logic_vector(27462, 16),
51083 => conv_std_logic_vector(27661, 16),
51084 => conv_std_logic_vector(27860, 16),
51085 => conv_std_logic_vector(28059, 16),
51086 => conv_std_logic_vector(28258, 16),
51087 => conv_std_logic_vector(28457, 16),
51088 => conv_std_logic_vector(28656, 16),
51089 => conv_std_logic_vector(28855, 16),
51090 => conv_std_logic_vector(29054, 16),
51091 => conv_std_logic_vector(29253, 16),
51092 => conv_std_logic_vector(29452, 16),
51093 => conv_std_logic_vector(29651, 16),
51094 => conv_std_logic_vector(29850, 16),
51095 => conv_std_logic_vector(30049, 16),
51096 => conv_std_logic_vector(30248, 16),
51097 => conv_std_logic_vector(30447, 16),
51098 => conv_std_logic_vector(30646, 16),
51099 => conv_std_logic_vector(30845, 16),
51100 => conv_std_logic_vector(31044, 16),
51101 => conv_std_logic_vector(31243, 16),
51102 => conv_std_logic_vector(31442, 16),
51103 => conv_std_logic_vector(31641, 16),
51104 => conv_std_logic_vector(31840, 16),
51105 => conv_std_logic_vector(32039, 16),
51106 => conv_std_logic_vector(32238, 16),
51107 => conv_std_logic_vector(32437, 16),
51108 => conv_std_logic_vector(32636, 16),
51109 => conv_std_logic_vector(32835, 16),
51110 => conv_std_logic_vector(33034, 16),
51111 => conv_std_logic_vector(33233, 16),
51112 => conv_std_logic_vector(33432, 16),
51113 => conv_std_logic_vector(33631, 16),
51114 => conv_std_logic_vector(33830, 16),
51115 => conv_std_logic_vector(34029, 16),
51116 => conv_std_logic_vector(34228, 16),
51117 => conv_std_logic_vector(34427, 16),
51118 => conv_std_logic_vector(34626, 16),
51119 => conv_std_logic_vector(34825, 16),
51120 => conv_std_logic_vector(35024, 16),
51121 => conv_std_logic_vector(35223, 16),
51122 => conv_std_logic_vector(35422, 16),
51123 => conv_std_logic_vector(35621, 16),
51124 => conv_std_logic_vector(35820, 16),
51125 => conv_std_logic_vector(36019, 16),
51126 => conv_std_logic_vector(36218, 16),
51127 => conv_std_logic_vector(36417, 16),
51128 => conv_std_logic_vector(36616, 16),
51129 => conv_std_logic_vector(36815, 16),
51130 => conv_std_logic_vector(37014, 16),
51131 => conv_std_logic_vector(37213, 16),
51132 => conv_std_logic_vector(37412, 16),
51133 => conv_std_logic_vector(37611, 16),
51134 => conv_std_logic_vector(37810, 16),
51135 => conv_std_logic_vector(38009, 16),
51136 => conv_std_logic_vector(38208, 16),
51137 => conv_std_logic_vector(38407, 16),
51138 => conv_std_logic_vector(38606, 16),
51139 => conv_std_logic_vector(38805, 16),
51140 => conv_std_logic_vector(39004, 16),
51141 => conv_std_logic_vector(39203, 16),
51142 => conv_std_logic_vector(39402, 16),
51143 => conv_std_logic_vector(39601, 16),
51144 => conv_std_logic_vector(39800, 16),
51145 => conv_std_logic_vector(39999, 16),
51146 => conv_std_logic_vector(40198, 16),
51147 => conv_std_logic_vector(40397, 16),
51148 => conv_std_logic_vector(40596, 16),
51149 => conv_std_logic_vector(40795, 16),
51150 => conv_std_logic_vector(40994, 16),
51151 => conv_std_logic_vector(41193, 16),
51152 => conv_std_logic_vector(41392, 16),
51153 => conv_std_logic_vector(41591, 16),
51154 => conv_std_logic_vector(41790, 16),
51155 => conv_std_logic_vector(41989, 16),
51156 => conv_std_logic_vector(42188, 16),
51157 => conv_std_logic_vector(42387, 16),
51158 => conv_std_logic_vector(42586, 16),
51159 => conv_std_logic_vector(42785, 16),
51160 => conv_std_logic_vector(42984, 16),
51161 => conv_std_logic_vector(43183, 16),
51162 => conv_std_logic_vector(43382, 16),
51163 => conv_std_logic_vector(43581, 16),
51164 => conv_std_logic_vector(43780, 16),
51165 => conv_std_logic_vector(43979, 16),
51166 => conv_std_logic_vector(44178, 16),
51167 => conv_std_logic_vector(44377, 16),
51168 => conv_std_logic_vector(44576, 16),
51169 => conv_std_logic_vector(44775, 16),
51170 => conv_std_logic_vector(44974, 16),
51171 => conv_std_logic_vector(45173, 16),
51172 => conv_std_logic_vector(45372, 16),
51173 => conv_std_logic_vector(45571, 16),
51174 => conv_std_logic_vector(45770, 16),
51175 => conv_std_logic_vector(45969, 16),
51176 => conv_std_logic_vector(46168, 16),
51177 => conv_std_logic_vector(46367, 16),
51178 => conv_std_logic_vector(46566, 16),
51179 => conv_std_logic_vector(46765, 16),
51180 => conv_std_logic_vector(46964, 16),
51181 => conv_std_logic_vector(47163, 16),
51182 => conv_std_logic_vector(47362, 16),
51183 => conv_std_logic_vector(47561, 16),
51184 => conv_std_logic_vector(47760, 16),
51185 => conv_std_logic_vector(47959, 16),
51186 => conv_std_logic_vector(48158, 16),
51187 => conv_std_logic_vector(48357, 16),
51188 => conv_std_logic_vector(48556, 16),
51189 => conv_std_logic_vector(48755, 16),
51190 => conv_std_logic_vector(48954, 16),
51191 => conv_std_logic_vector(49153, 16),
51192 => conv_std_logic_vector(49352, 16),
51193 => conv_std_logic_vector(49551, 16),
51194 => conv_std_logic_vector(49750, 16),
51195 => conv_std_logic_vector(49949, 16),
51196 => conv_std_logic_vector(50148, 16),
51197 => conv_std_logic_vector(50347, 16),
51198 => conv_std_logic_vector(50546, 16),
51199 => conv_std_logic_vector(50745, 16),
51200 => conv_std_logic_vector(0, 16),
51201 => conv_std_logic_vector(200, 16),
51202 => conv_std_logic_vector(400, 16),
51203 => conv_std_logic_vector(600, 16),
51204 => conv_std_logic_vector(800, 16),
51205 => conv_std_logic_vector(1000, 16),
51206 => conv_std_logic_vector(1200, 16),
51207 => conv_std_logic_vector(1400, 16),
51208 => conv_std_logic_vector(1600, 16),
51209 => conv_std_logic_vector(1800, 16),
51210 => conv_std_logic_vector(2000, 16),
51211 => conv_std_logic_vector(2200, 16),
51212 => conv_std_logic_vector(2400, 16),
51213 => conv_std_logic_vector(2600, 16),
51214 => conv_std_logic_vector(2800, 16),
51215 => conv_std_logic_vector(3000, 16),
51216 => conv_std_logic_vector(3200, 16),
51217 => conv_std_logic_vector(3400, 16),
51218 => conv_std_logic_vector(3600, 16),
51219 => conv_std_logic_vector(3800, 16),
51220 => conv_std_logic_vector(4000, 16),
51221 => conv_std_logic_vector(4200, 16),
51222 => conv_std_logic_vector(4400, 16),
51223 => conv_std_logic_vector(4600, 16),
51224 => conv_std_logic_vector(4800, 16),
51225 => conv_std_logic_vector(5000, 16),
51226 => conv_std_logic_vector(5200, 16),
51227 => conv_std_logic_vector(5400, 16),
51228 => conv_std_logic_vector(5600, 16),
51229 => conv_std_logic_vector(5800, 16),
51230 => conv_std_logic_vector(6000, 16),
51231 => conv_std_logic_vector(6200, 16),
51232 => conv_std_logic_vector(6400, 16),
51233 => conv_std_logic_vector(6600, 16),
51234 => conv_std_logic_vector(6800, 16),
51235 => conv_std_logic_vector(7000, 16),
51236 => conv_std_logic_vector(7200, 16),
51237 => conv_std_logic_vector(7400, 16),
51238 => conv_std_logic_vector(7600, 16),
51239 => conv_std_logic_vector(7800, 16),
51240 => conv_std_logic_vector(8000, 16),
51241 => conv_std_logic_vector(8200, 16),
51242 => conv_std_logic_vector(8400, 16),
51243 => conv_std_logic_vector(8600, 16),
51244 => conv_std_logic_vector(8800, 16),
51245 => conv_std_logic_vector(9000, 16),
51246 => conv_std_logic_vector(9200, 16),
51247 => conv_std_logic_vector(9400, 16),
51248 => conv_std_logic_vector(9600, 16),
51249 => conv_std_logic_vector(9800, 16),
51250 => conv_std_logic_vector(10000, 16),
51251 => conv_std_logic_vector(10200, 16),
51252 => conv_std_logic_vector(10400, 16),
51253 => conv_std_logic_vector(10600, 16),
51254 => conv_std_logic_vector(10800, 16),
51255 => conv_std_logic_vector(11000, 16),
51256 => conv_std_logic_vector(11200, 16),
51257 => conv_std_logic_vector(11400, 16),
51258 => conv_std_logic_vector(11600, 16),
51259 => conv_std_logic_vector(11800, 16),
51260 => conv_std_logic_vector(12000, 16),
51261 => conv_std_logic_vector(12200, 16),
51262 => conv_std_logic_vector(12400, 16),
51263 => conv_std_logic_vector(12600, 16),
51264 => conv_std_logic_vector(12800, 16),
51265 => conv_std_logic_vector(13000, 16),
51266 => conv_std_logic_vector(13200, 16),
51267 => conv_std_logic_vector(13400, 16),
51268 => conv_std_logic_vector(13600, 16),
51269 => conv_std_logic_vector(13800, 16),
51270 => conv_std_logic_vector(14000, 16),
51271 => conv_std_logic_vector(14200, 16),
51272 => conv_std_logic_vector(14400, 16),
51273 => conv_std_logic_vector(14600, 16),
51274 => conv_std_logic_vector(14800, 16),
51275 => conv_std_logic_vector(15000, 16),
51276 => conv_std_logic_vector(15200, 16),
51277 => conv_std_logic_vector(15400, 16),
51278 => conv_std_logic_vector(15600, 16),
51279 => conv_std_logic_vector(15800, 16),
51280 => conv_std_logic_vector(16000, 16),
51281 => conv_std_logic_vector(16200, 16),
51282 => conv_std_logic_vector(16400, 16),
51283 => conv_std_logic_vector(16600, 16),
51284 => conv_std_logic_vector(16800, 16),
51285 => conv_std_logic_vector(17000, 16),
51286 => conv_std_logic_vector(17200, 16),
51287 => conv_std_logic_vector(17400, 16),
51288 => conv_std_logic_vector(17600, 16),
51289 => conv_std_logic_vector(17800, 16),
51290 => conv_std_logic_vector(18000, 16),
51291 => conv_std_logic_vector(18200, 16),
51292 => conv_std_logic_vector(18400, 16),
51293 => conv_std_logic_vector(18600, 16),
51294 => conv_std_logic_vector(18800, 16),
51295 => conv_std_logic_vector(19000, 16),
51296 => conv_std_logic_vector(19200, 16),
51297 => conv_std_logic_vector(19400, 16),
51298 => conv_std_logic_vector(19600, 16),
51299 => conv_std_logic_vector(19800, 16),
51300 => conv_std_logic_vector(20000, 16),
51301 => conv_std_logic_vector(20200, 16),
51302 => conv_std_logic_vector(20400, 16),
51303 => conv_std_logic_vector(20600, 16),
51304 => conv_std_logic_vector(20800, 16),
51305 => conv_std_logic_vector(21000, 16),
51306 => conv_std_logic_vector(21200, 16),
51307 => conv_std_logic_vector(21400, 16),
51308 => conv_std_logic_vector(21600, 16),
51309 => conv_std_logic_vector(21800, 16),
51310 => conv_std_logic_vector(22000, 16),
51311 => conv_std_logic_vector(22200, 16),
51312 => conv_std_logic_vector(22400, 16),
51313 => conv_std_logic_vector(22600, 16),
51314 => conv_std_logic_vector(22800, 16),
51315 => conv_std_logic_vector(23000, 16),
51316 => conv_std_logic_vector(23200, 16),
51317 => conv_std_logic_vector(23400, 16),
51318 => conv_std_logic_vector(23600, 16),
51319 => conv_std_logic_vector(23800, 16),
51320 => conv_std_logic_vector(24000, 16),
51321 => conv_std_logic_vector(24200, 16),
51322 => conv_std_logic_vector(24400, 16),
51323 => conv_std_logic_vector(24600, 16),
51324 => conv_std_logic_vector(24800, 16),
51325 => conv_std_logic_vector(25000, 16),
51326 => conv_std_logic_vector(25200, 16),
51327 => conv_std_logic_vector(25400, 16),
51328 => conv_std_logic_vector(25600, 16),
51329 => conv_std_logic_vector(25800, 16),
51330 => conv_std_logic_vector(26000, 16),
51331 => conv_std_logic_vector(26200, 16),
51332 => conv_std_logic_vector(26400, 16),
51333 => conv_std_logic_vector(26600, 16),
51334 => conv_std_logic_vector(26800, 16),
51335 => conv_std_logic_vector(27000, 16),
51336 => conv_std_logic_vector(27200, 16),
51337 => conv_std_logic_vector(27400, 16),
51338 => conv_std_logic_vector(27600, 16),
51339 => conv_std_logic_vector(27800, 16),
51340 => conv_std_logic_vector(28000, 16),
51341 => conv_std_logic_vector(28200, 16),
51342 => conv_std_logic_vector(28400, 16),
51343 => conv_std_logic_vector(28600, 16),
51344 => conv_std_logic_vector(28800, 16),
51345 => conv_std_logic_vector(29000, 16),
51346 => conv_std_logic_vector(29200, 16),
51347 => conv_std_logic_vector(29400, 16),
51348 => conv_std_logic_vector(29600, 16),
51349 => conv_std_logic_vector(29800, 16),
51350 => conv_std_logic_vector(30000, 16),
51351 => conv_std_logic_vector(30200, 16),
51352 => conv_std_logic_vector(30400, 16),
51353 => conv_std_logic_vector(30600, 16),
51354 => conv_std_logic_vector(30800, 16),
51355 => conv_std_logic_vector(31000, 16),
51356 => conv_std_logic_vector(31200, 16),
51357 => conv_std_logic_vector(31400, 16),
51358 => conv_std_logic_vector(31600, 16),
51359 => conv_std_logic_vector(31800, 16),
51360 => conv_std_logic_vector(32000, 16),
51361 => conv_std_logic_vector(32200, 16),
51362 => conv_std_logic_vector(32400, 16),
51363 => conv_std_logic_vector(32600, 16),
51364 => conv_std_logic_vector(32800, 16),
51365 => conv_std_logic_vector(33000, 16),
51366 => conv_std_logic_vector(33200, 16),
51367 => conv_std_logic_vector(33400, 16),
51368 => conv_std_logic_vector(33600, 16),
51369 => conv_std_logic_vector(33800, 16),
51370 => conv_std_logic_vector(34000, 16),
51371 => conv_std_logic_vector(34200, 16),
51372 => conv_std_logic_vector(34400, 16),
51373 => conv_std_logic_vector(34600, 16),
51374 => conv_std_logic_vector(34800, 16),
51375 => conv_std_logic_vector(35000, 16),
51376 => conv_std_logic_vector(35200, 16),
51377 => conv_std_logic_vector(35400, 16),
51378 => conv_std_logic_vector(35600, 16),
51379 => conv_std_logic_vector(35800, 16),
51380 => conv_std_logic_vector(36000, 16),
51381 => conv_std_logic_vector(36200, 16),
51382 => conv_std_logic_vector(36400, 16),
51383 => conv_std_logic_vector(36600, 16),
51384 => conv_std_logic_vector(36800, 16),
51385 => conv_std_logic_vector(37000, 16),
51386 => conv_std_logic_vector(37200, 16),
51387 => conv_std_logic_vector(37400, 16),
51388 => conv_std_logic_vector(37600, 16),
51389 => conv_std_logic_vector(37800, 16),
51390 => conv_std_logic_vector(38000, 16),
51391 => conv_std_logic_vector(38200, 16),
51392 => conv_std_logic_vector(38400, 16),
51393 => conv_std_logic_vector(38600, 16),
51394 => conv_std_logic_vector(38800, 16),
51395 => conv_std_logic_vector(39000, 16),
51396 => conv_std_logic_vector(39200, 16),
51397 => conv_std_logic_vector(39400, 16),
51398 => conv_std_logic_vector(39600, 16),
51399 => conv_std_logic_vector(39800, 16),
51400 => conv_std_logic_vector(40000, 16),
51401 => conv_std_logic_vector(40200, 16),
51402 => conv_std_logic_vector(40400, 16),
51403 => conv_std_logic_vector(40600, 16),
51404 => conv_std_logic_vector(40800, 16),
51405 => conv_std_logic_vector(41000, 16),
51406 => conv_std_logic_vector(41200, 16),
51407 => conv_std_logic_vector(41400, 16),
51408 => conv_std_logic_vector(41600, 16),
51409 => conv_std_logic_vector(41800, 16),
51410 => conv_std_logic_vector(42000, 16),
51411 => conv_std_logic_vector(42200, 16),
51412 => conv_std_logic_vector(42400, 16),
51413 => conv_std_logic_vector(42600, 16),
51414 => conv_std_logic_vector(42800, 16),
51415 => conv_std_logic_vector(43000, 16),
51416 => conv_std_logic_vector(43200, 16),
51417 => conv_std_logic_vector(43400, 16),
51418 => conv_std_logic_vector(43600, 16),
51419 => conv_std_logic_vector(43800, 16),
51420 => conv_std_logic_vector(44000, 16),
51421 => conv_std_logic_vector(44200, 16),
51422 => conv_std_logic_vector(44400, 16),
51423 => conv_std_logic_vector(44600, 16),
51424 => conv_std_logic_vector(44800, 16),
51425 => conv_std_logic_vector(45000, 16),
51426 => conv_std_logic_vector(45200, 16),
51427 => conv_std_logic_vector(45400, 16),
51428 => conv_std_logic_vector(45600, 16),
51429 => conv_std_logic_vector(45800, 16),
51430 => conv_std_logic_vector(46000, 16),
51431 => conv_std_logic_vector(46200, 16),
51432 => conv_std_logic_vector(46400, 16),
51433 => conv_std_logic_vector(46600, 16),
51434 => conv_std_logic_vector(46800, 16),
51435 => conv_std_logic_vector(47000, 16),
51436 => conv_std_logic_vector(47200, 16),
51437 => conv_std_logic_vector(47400, 16),
51438 => conv_std_logic_vector(47600, 16),
51439 => conv_std_logic_vector(47800, 16),
51440 => conv_std_logic_vector(48000, 16),
51441 => conv_std_logic_vector(48200, 16),
51442 => conv_std_logic_vector(48400, 16),
51443 => conv_std_logic_vector(48600, 16),
51444 => conv_std_logic_vector(48800, 16),
51445 => conv_std_logic_vector(49000, 16),
51446 => conv_std_logic_vector(49200, 16),
51447 => conv_std_logic_vector(49400, 16),
51448 => conv_std_logic_vector(49600, 16),
51449 => conv_std_logic_vector(49800, 16),
51450 => conv_std_logic_vector(50000, 16),
51451 => conv_std_logic_vector(50200, 16),
51452 => conv_std_logic_vector(50400, 16),
51453 => conv_std_logic_vector(50600, 16),
51454 => conv_std_logic_vector(50800, 16),
51455 => conv_std_logic_vector(51000, 16),
51456 => conv_std_logic_vector(0, 16),
51457 => conv_std_logic_vector(201, 16),
51458 => conv_std_logic_vector(402, 16),
51459 => conv_std_logic_vector(603, 16),
51460 => conv_std_logic_vector(804, 16),
51461 => conv_std_logic_vector(1005, 16),
51462 => conv_std_logic_vector(1206, 16),
51463 => conv_std_logic_vector(1407, 16),
51464 => conv_std_logic_vector(1608, 16),
51465 => conv_std_logic_vector(1809, 16),
51466 => conv_std_logic_vector(2010, 16),
51467 => conv_std_logic_vector(2211, 16),
51468 => conv_std_logic_vector(2412, 16),
51469 => conv_std_logic_vector(2613, 16),
51470 => conv_std_logic_vector(2814, 16),
51471 => conv_std_logic_vector(3015, 16),
51472 => conv_std_logic_vector(3216, 16),
51473 => conv_std_logic_vector(3417, 16),
51474 => conv_std_logic_vector(3618, 16),
51475 => conv_std_logic_vector(3819, 16),
51476 => conv_std_logic_vector(4020, 16),
51477 => conv_std_logic_vector(4221, 16),
51478 => conv_std_logic_vector(4422, 16),
51479 => conv_std_logic_vector(4623, 16),
51480 => conv_std_logic_vector(4824, 16),
51481 => conv_std_logic_vector(5025, 16),
51482 => conv_std_logic_vector(5226, 16),
51483 => conv_std_logic_vector(5427, 16),
51484 => conv_std_logic_vector(5628, 16),
51485 => conv_std_logic_vector(5829, 16),
51486 => conv_std_logic_vector(6030, 16),
51487 => conv_std_logic_vector(6231, 16),
51488 => conv_std_logic_vector(6432, 16),
51489 => conv_std_logic_vector(6633, 16),
51490 => conv_std_logic_vector(6834, 16),
51491 => conv_std_logic_vector(7035, 16),
51492 => conv_std_logic_vector(7236, 16),
51493 => conv_std_logic_vector(7437, 16),
51494 => conv_std_logic_vector(7638, 16),
51495 => conv_std_logic_vector(7839, 16),
51496 => conv_std_logic_vector(8040, 16),
51497 => conv_std_logic_vector(8241, 16),
51498 => conv_std_logic_vector(8442, 16),
51499 => conv_std_logic_vector(8643, 16),
51500 => conv_std_logic_vector(8844, 16),
51501 => conv_std_logic_vector(9045, 16),
51502 => conv_std_logic_vector(9246, 16),
51503 => conv_std_logic_vector(9447, 16),
51504 => conv_std_logic_vector(9648, 16),
51505 => conv_std_logic_vector(9849, 16),
51506 => conv_std_logic_vector(10050, 16),
51507 => conv_std_logic_vector(10251, 16),
51508 => conv_std_logic_vector(10452, 16),
51509 => conv_std_logic_vector(10653, 16),
51510 => conv_std_logic_vector(10854, 16),
51511 => conv_std_logic_vector(11055, 16),
51512 => conv_std_logic_vector(11256, 16),
51513 => conv_std_logic_vector(11457, 16),
51514 => conv_std_logic_vector(11658, 16),
51515 => conv_std_logic_vector(11859, 16),
51516 => conv_std_logic_vector(12060, 16),
51517 => conv_std_logic_vector(12261, 16),
51518 => conv_std_logic_vector(12462, 16),
51519 => conv_std_logic_vector(12663, 16),
51520 => conv_std_logic_vector(12864, 16),
51521 => conv_std_logic_vector(13065, 16),
51522 => conv_std_logic_vector(13266, 16),
51523 => conv_std_logic_vector(13467, 16),
51524 => conv_std_logic_vector(13668, 16),
51525 => conv_std_logic_vector(13869, 16),
51526 => conv_std_logic_vector(14070, 16),
51527 => conv_std_logic_vector(14271, 16),
51528 => conv_std_logic_vector(14472, 16),
51529 => conv_std_logic_vector(14673, 16),
51530 => conv_std_logic_vector(14874, 16),
51531 => conv_std_logic_vector(15075, 16),
51532 => conv_std_logic_vector(15276, 16),
51533 => conv_std_logic_vector(15477, 16),
51534 => conv_std_logic_vector(15678, 16),
51535 => conv_std_logic_vector(15879, 16),
51536 => conv_std_logic_vector(16080, 16),
51537 => conv_std_logic_vector(16281, 16),
51538 => conv_std_logic_vector(16482, 16),
51539 => conv_std_logic_vector(16683, 16),
51540 => conv_std_logic_vector(16884, 16),
51541 => conv_std_logic_vector(17085, 16),
51542 => conv_std_logic_vector(17286, 16),
51543 => conv_std_logic_vector(17487, 16),
51544 => conv_std_logic_vector(17688, 16),
51545 => conv_std_logic_vector(17889, 16),
51546 => conv_std_logic_vector(18090, 16),
51547 => conv_std_logic_vector(18291, 16),
51548 => conv_std_logic_vector(18492, 16),
51549 => conv_std_logic_vector(18693, 16),
51550 => conv_std_logic_vector(18894, 16),
51551 => conv_std_logic_vector(19095, 16),
51552 => conv_std_logic_vector(19296, 16),
51553 => conv_std_logic_vector(19497, 16),
51554 => conv_std_logic_vector(19698, 16),
51555 => conv_std_logic_vector(19899, 16),
51556 => conv_std_logic_vector(20100, 16),
51557 => conv_std_logic_vector(20301, 16),
51558 => conv_std_logic_vector(20502, 16),
51559 => conv_std_logic_vector(20703, 16),
51560 => conv_std_logic_vector(20904, 16),
51561 => conv_std_logic_vector(21105, 16),
51562 => conv_std_logic_vector(21306, 16),
51563 => conv_std_logic_vector(21507, 16),
51564 => conv_std_logic_vector(21708, 16),
51565 => conv_std_logic_vector(21909, 16),
51566 => conv_std_logic_vector(22110, 16),
51567 => conv_std_logic_vector(22311, 16),
51568 => conv_std_logic_vector(22512, 16),
51569 => conv_std_logic_vector(22713, 16),
51570 => conv_std_logic_vector(22914, 16),
51571 => conv_std_logic_vector(23115, 16),
51572 => conv_std_logic_vector(23316, 16),
51573 => conv_std_logic_vector(23517, 16),
51574 => conv_std_logic_vector(23718, 16),
51575 => conv_std_logic_vector(23919, 16),
51576 => conv_std_logic_vector(24120, 16),
51577 => conv_std_logic_vector(24321, 16),
51578 => conv_std_logic_vector(24522, 16),
51579 => conv_std_logic_vector(24723, 16),
51580 => conv_std_logic_vector(24924, 16),
51581 => conv_std_logic_vector(25125, 16),
51582 => conv_std_logic_vector(25326, 16),
51583 => conv_std_logic_vector(25527, 16),
51584 => conv_std_logic_vector(25728, 16),
51585 => conv_std_logic_vector(25929, 16),
51586 => conv_std_logic_vector(26130, 16),
51587 => conv_std_logic_vector(26331, 16),
51588 => conv_std_logic_vector(26532, 16),
51589 => conv_std_logic_vector(26733, 16),
51590 => conv_std_logic_vector(26934, 16),
51591 => conv_std_logic_vector(27135, 16),
51592 => conv_std_logic_vector(27336, 16),
51593 => conv_std_logic_vector(27537, 16),
51594 => conv_std_logic_vector(27738, 16),
51595 => conv_std_logic_vector(27939, 16),
51596 => conv_std_logic_vector(28140, 16),
51597 => conv_std_logic_vector(28341, 16),
51598 => conv_std_logic_vector(28542, 16),
51599 => conv_std_logic_vector(28743, 16),
51600 => conv_std_logic_vector(28944, 16),
51601 => conv_std_logic_vector(29145, 16),
51602 => conv_std_logic_vector(29346, 16),
51603 => conv_std_logic_vector(29547, 16),
51604 => conv_std_logic_vector(29748, 16),
51605 => conv_std_logic_vector(29949, 16),
51606 => conv_std_logic_vector(30150, 16),
51607 => conv_std_logic_vector(30351, 16),
51608 => conv_std_logic_vector(30552, 16),
51609 => conv_std_logic_vector(30753, 16),
51610 => conv_std_logic_vector(30954, 16),
51611 => conv_std_logic_vector(31155, 16),
51612 => conv_std_logic_vector(31356, 16),
51613 => conv_std_logic_vector(31557, 16),
51614 => conv_std_logic_vector(31758, 16),
51615 => conv_std_logic_vector(31959, 16),
51616 => conv_std_logic_vector(32160, 16),
51617 => conv_std_logic_vector(32361, 16),
51618 => conv_std_logic_vector(32562, 16),
51619 => conv_std_logic_vector(32763, 16),
51620 => conv_std_logic_vector(32964, 16),
51621 => conv_std_logic_vector(33165, 16),
51622 => conv_std_logic_vector(33366, 16),
51623 => conv_std_logic_vector(33567, 16),
51624 => conv_std_logic_vector(33768, 16),
51625 => conv_std_logic_vector(33969, 16),
51626 => conv_std_logic_vector(34170, 16),
51627 => conv_std_logic_vector(34371, 16),
51628 => conv_std_logic_vector(34572, 16),
51629 => conv_std_logic_vector(34773, 16),
51630 => conv_std_logic_vector(34974, 16),
51631 => conv_std_logic_vector(35175, 16),
51632 => conv_std_logic_vector(35376, 16),
51633 => conv_std_logic_vector(35577, 16),
51634 => conv_std_logic_vector(35778, 16),
51635 => conv_std_logic_vector(35979, 16),
51636 => conv_std_logic_vector(36180, 16),
51637 => conv_std_logic_vector(36381, 16),
51638 => conv_std_logic_vector(36582, 16),
51639 => conv_std_logic_vector(36783, 16),
51640 => conv_std_logic_vector(36984, 16),
51641 => conv_std_logic_vector(37185, 16),
51642 => conv_std_logic_vector(37386, 16),
51643 => conv_std_logic_vector(37587, 16),
51644 => conv_std_logic_vector(37788, 16),
51645 => conv_std_logic_vector(37989, 16),
51646 => conv_std_logic_vector(38190, 16),
51647 => conv_std_logic_vector(38391, 16),
51648 => conv_std_logic_vector(38592, 16),
51649 => conv_std_logic_vector(38793, 16),
51650 => conv_std_logic_vector(38994, 16),
51651 => conv_std_logic_vector(39195, 16),
51652 => conv_std_logic_vector(39396, 16),
51653 => conv_std_logic_vector(39597, 16),
51654 => conv_std_logic_vector(39798, 16),
51655 => conv_std_logic_vector(39999, 16),
51656 => conv_std_logic_vector(40200, 16),
51657 => conv_std_logic_vector(40401, 16),
51658 => conv_std_logic_vector(40602, 16),
51659 => conv_std_logic_vector(40803, 16),
51660 => conv_std_logic_vector(41004, 16),
51661 => conv_std_logic_vector(41205, 16),
51662 => conv_std_logic_vector(41406, 16),
51663 => conv_std_logic_vector(41607, 16),
51664 => conv_std_logic_vector(41808, 16),
51665 => conv_std_logic_vector(42009, 16),
51666 => conv_std_logic_vector(42210, 16),
51667 => conv_std_logic_vector(42411, 16),
51668 => conv_std_logic_vector(42612, 16),
51669 => conv_std_logic_vector(42813, 16),
51670 => conv_std_logic_vector(43014, 16),
51671 => conv_std_logic_vector(43215, 16),
51672 => conv_std_logic_vector(43416, 16),
51673 => conv_std_logic_vector(43617, 16),
51674 => conv_std_logic_vector(43818, 16),
51675 => conv_std_logic_vector(44019, 16),
51676 => conv_std_logic_vector(44220, 16),
51677 => conv_std_logic_vector(44421, 16),
51678 => conv_std_logic_vector(44622, 16),
51679 => conv_std_logic_vector(44823, 16),
51680 => conv_std_logic_vector(45024, 16),
51681 => conv_std_logic_vector(45225, 16),
51682 => conv_std_logic_vector(45426, 16),
51683 => conv_std_logic_vector(45627, 16),
51684 => conv_std_logic_vector(45828, 16),
51685 => conv_std_logic_vector(46029, 16),
51686 => conv_std_logic_vector(46230, 16),
51687 => conv_std_logic_vector(46431, 16),
51688 => conv_std_logic_vector(46632, 16),
51689 => conv_std_logic_vector(46833, 16),
51690 => conv_std_logic_vector(47034, 16),
51691 => conv_std_logic_vector(47235, 16),
51692 => conv_std_logic_vector(47436, 16),
51693 => conv_std_logic_vector(47637, 16),
51694 => conv_std_logic_vector(47838, 16),
51695 => conv_std_logic_vector(48039, 16),
51696 => conv_std_logic_vector(48240, 16),
51697 => conv_std_logic_vector(48441, 16),
51698 => conv_std_logic_vector(48642, 16),
51699 => conv_std_logic_vector(48843, 16),
51700 => conv_std_logic_vector(49044, 16),
51701 => conv_std_logic_vector(49245, 16),
51702 => conv_std_logic_vector(49446, 16),
51703 => conv_std_logic_vector(49647, 16),
51704 => conv_std_logic_vector(49848, 16),
51705 => conv_std_logic_vector(50049, 16),
51706 => conv_std_logic_vector(50250, 16),
51707 => conv_std_logic_vector(50451, 16),
51708 => conv_std_logic_vector(50652, 16),
51709 => conv_std_logic_vector(50853, 16),
51710 => conv_std_logic_vector(51054, 16),
51711 => conv_std_logic_vector(51255, 16),
51712 => conv_std_logic_vector(0, 16),
51713 => conv_std_logic_vector(202, 16),
51714 => conv_std_logic_vector(404, 16),
51715 => conv_std_logic_vector(606, 16),
51716 => conv_std_logic_vector(808, 16),
51717 => conv_std_logic_vector(1010, 16),
51718 => conv_std_logic_vector(1212, 16),
51719 => conv_std_logic_vector(1414, 16),
51720 => conv_std_logic_vector(1616, 16),
51721 => conv_std_logic_vector(1818, 16),
51722 => conv_std_logic_vector(2020, 16),
51723 => conv_std_logic_vector(2222, 16),
51724 => conv_std_logic_vector(2424, 16),
51725 => conv_std_logic_vector(2626, 16),
51726 => conv_std_logic_vector(2828, 16),
51727 => conv_std_logic_vector(3030, 16),
51728 => conv_std_logic_vector(3232, 16),
51729 => conv_std_logic_vector(3434, 16),
51730 => conv_std_logic_vector(3636, 16),
51731 => conv_std_logic_vector(3838, 16),
51732 => conv_std_logic_vector(4040, 16),
51733 => conv_std_logic_vector(4242, 16),
51734 => conv_std_logic_vector(4444, 16),
51735 => conv_std_logic_vector(4646, 16),
51736 => conv_std_logic_vector(4848, 16),
51737 => conv_std_logic_vector(5050, 16),
51738 => conv_std_logic_vector(5252, 16),
51739 => conv_std_logic_vector(5454, 16),
51740 => conv_std_logic_vector(5656, 16),
51741 => conv_std_logic_vector(5858, 16),
51742 => conv_std_logic_vector(6060, 16),
51743 => conv_std_logic_vector(6262, 16),
51744 => conv_std_logic_vector(6464, 16),
51745 => conv_std_logic_vector(6666, 16),
51746 => conv_std_logic_vector(6868, 16),
51747 => conv_std_logic_vector(7070, 16),
51748 => conv_std_logic_vector(7272, 16),
51749 => conv_std_logic_vector(7474, 16),
51750 => conv_std_logic_vector(7676, 16),
51751 => conv_std_logic_vector(7878, 16),
51752 => conv_std_logic_vector(8080, 16),
51753 => conv_std_logic_vector(8282, 16),
51754 => conv_std_logic_vector(8484, 16),
51755 => conv_std_logic_vector(8686, 16),
51756 => conv_std_logic_vector(8888, 16),
51757 => conv_std_logic_vector(9090, 16),
51758 => conv_std_logic_vector(9292, 16),
51759 => conv_std_logic_vector(9494, 16),
51760 => conv_std_logic_vector(9696, 16),
51761 => conv_std_logic_vector(9898, 16),
51762 => conv_std_logic_vector(10100, 16),
51763 => conv_std_logic_vector(10302, 16),
51764 => conv_std_logic_vector(10504, 16),
51765 => conv_std_logic_vector(10706, 16),
51766 => conv_std_logic_vector(10908, 16),
51767 => conv_std_logic_vector(11110, 16),
51768 => conv_std_logic_vector(11312, 16),
51769 => conv_std_logic_vector(11514, 16),
51770 => conv_std_logic_vector(11716, 16),
51771 => conv_std_logic_vector(11918, 16),
51772 => conv_std_logic_vector(12120, 16),
51773 => conv_std_logic_vector(12322, 16),
51774 => conv_std_logic_vector(12524, 16),
51775 => conv_std_logic_vector(12726, 16),
51776 => conv_std_logic_vector(12928, 16),
51777 => conv_std_logic_vector(13130, 16),
51778 => conv_std_logic_vector(13332, 16),
51779 => conv_std_logic_vector(13534, 16),
51780 => conv_std_logic_vector(13736, 16),
51781 => conv_std_logic_vector(13938, 16),
51782 => conv_std_logic_vector(14140, 16),
51783 => conv_std_logic_vector(14342, 16),
51784 => conv_std_logic_vector(14544, 16),
51785 => conv_std_logic_vector(14746, 16),
51786 => conv_std_logic_vector(14948, 16),
51787 => conv_std_logic_vector(15150, 16),
51788 => conv_std_logic_vector(15352, 16),
51789 => conv_std_logic_vector(15554, 16),
51790 => conv_std_logic_vector(15756, 16),
51791 => conv_std_logic_vector(15958, 16),
51792 => conv_std_logic_vector(16160, 16),
51793 => conv_std_logic_vector(16362, 16),
51794 => conv_std_logic_vector(16564, 16),
51795 => conv_std_logic_vector(16766, 16),
51796 => conv_std_logic_vector(16968, 16),
51797 => conv_std_logic_vector(17170, 16),
51798 => conv_std_logic_vector(17372, 16),
51799 => conv_std_logic_vector(17574, 16),
51800 => conv_std_logic_vector(17776, 16),
51801 => conv_std_logic_vector(17978, 16),
51802 => conv_std_logic_vector(18180, 16),
51803 => conv_std_logic_vector(18382, 16),
51804 => conv_std_logic_vector(18584, 16),
51805 => conv_std_logic_vector(18786, 16),
51806 => conv_std_logic_vector(18988, 16),
51807 => conv_std_logic_vector(19190, 16),
51808 => conv_std_logic_vector(19392, 16),
51809 => conv_std_logic_vector(19594, 16),
51810 => conv_std_logic_vector(19796, 16),
51811 => conv_std_logic_vector(19998, 16),
51812 => conv_std_logic_vector(20200, 16),
51813 => conv_std_logic_vector(20402, 16),
51814 => conv_std_logic_vector(20604, 16),
51815 => conv_std_logic_vector(20806, 16),
51816 => conv_std_logic_vector(21008, 16),
51817 => conv_std_logic_vector(21210, 16),
51818 => conv_std_logic_vector(21412, 16),
51819 => conv_std_logic_vector(21614, 16),
51820 => conv_std_logic_vector(21816, 16),
51821 => conv_std_logic_vector(22018, 16),
51822 => conv_std_logic_vector(22220, 16),
51823 => conv_std_logic_vector(22422, 16),
51824 => conv_std_logic_vector(22624, 16),
51825 => conv_std_logic_vector(22826, 16),
51826 => conv_std_logic_vector(23028, 16),
51827 => conv_std_logic_vector(23230, 16),
51828 => conv_std_logic_vector(23432, 16),
51829 => conv_std_logic_vector(23634, 16),
51830 => conv_std_logic_vector(23836, 16),
51831 => conv_std_logic_vector(24038, 16),
51832 => conv_std_logic_vector(24240, 16),
51833 => conv_std_logic_vector(24442, 16),
51834 => conv_std_logic_vector(24644, 16),
51835 => conv_std_logic_vector(24846, 16),
51836 => conv_std_logic_vector(25048, 16),
51837 => conv_std_logic_vector(25250, 16),
51838 => conv_std_logic_vector(25452, 16),
51839 => conv_std_logic_vector(25654, 16),
51840 => conv_std_logic_vector(25856, 16),
51841 => conv_std_logic_vector(26058, 16),
51842 => conv_std_logic_vector(26260, 16),
51843 => conv_std_logic_vector(26462, 16),
51844 => conv_std_logic_vector(26664, 16),
51845 => conv_std_logic_vector(26866, 16),
51846 => conv_std_logic_vector(27068, 16),
51847 => conv_std_logic_vector(27270, 16),
51848 => conv_std_logic_vector(27472, 16),
51849 => conv_std_logic_vector(27674, 16),
51850 => conv_std_logic_vector(27876, 16),
51851 => conv_std_logic_vector(28078, 16),
51852 => conv_std_logic_vector(28280, 16),
51853 => conv_std_logic_vector(28482, 16),
51854 => conv_std_logic_vector(28684, 16),
51855 => conv_std_logic_vector(28886, 16),
51856 => conv_std_logic_vector(29088, 16),
51857 => conv_std_logic_vector(29290, 16),
51858 => conv_std_logic_vector(29492, 16),
51859 => conv_std_logic_vector(29694, 16),
51860 => conv_std_logic_vector(29896, 16),
51861 => conv_std_logic_vector(30098, 16),
51862 => conv_std_logic_vector(30300, 16),
51863 => conv_std_logic_vector(30502, 16),
51864 => conv_std_logic_vector(30704, 16),
51865 => conv_std_logic_vector(30906, 16),
51866 => conv_std_logic_vector(31108, 16),
51867 => conv_std_logic_vector(31310, 16),
51868 => conv_std_logic_vector(31512, 16),
51869 => conv_std_logic_vector(31714, 16),
51870 => conv_std_logic_vector(31916, 16),
51871 => conv_std_logic_vector(32118, 16),
51872 => conv_std_logic_vector(32320, 16),
51873 => conv_std_logic_vector(32522, 16),
51874 => conv_std_logic_vector(32724, 16),
51875 => conv_std_logic_vector(32926, 16),
51876 => conv_std_logic_vector(33128, 16),
51877 => conv_std_logic_vector(33330, 16),
51878 => conv_std_logic_vector(33532, 16),
51879 => conv_std_logic_vector(33734, 16),
51880 => conv_std_logic_vector(33936, 16),
51881 => conv_std_logic_vector(34138, 16),
51882 => conv_std_logic_vector(34340, 16),
51883 => conv_std_logic_vector(34542, 16),
51884 => conv_std_logic_vector(34744, 16),
51885 => conv_std_logic_vector(34946, 16),
51886 => conv_std_logic_vector(35148, 16),
51887 => conv_std_logic_vector(35350, 16),
51888 => conv_std_logic_vector(35552, 16),
51889 => conv_std_logic_vector(35754, 16),
51890 => conv_std_logic_vector(35956, 16),
51891 => conv_std_logic_vector(36158, 16),
51892 => conv_std_logic_vector(36360, 16),
51893 => conv_std_logic_vector(36562, 16),
51894 => conv_std_logic_vector(36764, 16),
51895 => conv_std_logic_vector(36966, 16),
51896 => conv_std_logic_vector(37168, 16),
51897 => conv_std_logic_vector(37370, 16),
51898 => conv_std_logic_vector(37572, 16),
51899 => conv_std_logic_vector(37774, 16),
51900 => conv_std_logic_vector(37976, 16),
51901 => conv_std_logic_vector(38178, 16),
51902 => conv_std_logic_vector(38380, 16),
51903 => conv_std_logic_vector(38582, 16),
51904 => conv_std_logic_vector(38784, 16),
51905 => conv_std_logic_vector(38986, 16),
51906 => conv_std_logic_vector(39188, 16),
51907 => conv_std_logic_vector(39390, 16),
51908 => conv_std_logic_vector(39592, 16),
51909 => conv_std_logic_vector(39794, 16),
51910 => conv_std_logic_vector(39996, 16),
51911 => conv_std_logic_vector(40198, 16),
51912 => conv_std_logic_vector(40400, 16),
51913 => conv_std_logic_vector(40602, 16),
51914 => conv_std_logic_vector(40804, 16),
51915 => conv_std_logic_vector(41006, 16),
51916 => conv_std_logic_vector(41208, 16),
51917 => conv_std_logic_vector(41410, 16),
51918 => conv_std_logic_vector(41612, 16),
51919 => conv_std_logic_vector(41814, 16),
51920 => conv_std_logic_vector(42016, 16),
51921 => conv_std_logic_vector(42218, 16),
51922 => conv_std_logic_vector(42420, 16),
51923 => conv_std_logic_vector(42622, 16),
51924 => conv_std_logic_vector(42824, 16),
51925 => conv_std_logic_vector(43026, 16),
51926 => conv_std_logic_vector(43228, 16),
51927 => conv_std_logic_vector(43430, 16),
51928 => conv_std_logic_vector(43632, 16),
51929 => conv_std_logic_vector(43834, 16),
51930 => conv_std_logic_vector(44036, 16),
51931 => conv_std_logic_vector(44238, 16),
51932 => conv_std_logic_vector(44440, 16),
51933 => conv_std_logic_vector(44642, 16),
51934 => conv_std_logic_vector(44844, 16),
51935 => conv_std_logic_vector(45046, 16),
51936 => conv_std_logic_vector(45248, 16),
51937 => conv_std_logic_vector(45450, 16),
51938 => conv_std_logic_vector(45652, 16),
51939 => conv_std_logic_vector(45854, 16),
51940 => conv_std_logic_vector(46056, 16),
51941 => conv_std_logic_vector(46258, 16),
51942 => conv_std_logic_vector(46460, 16),
51943 => conv_std_logic_vector(46662, 16),
51944 => conv_std_logic_vector(46864, 16),
51945 => conv_std_logic_vector(47066, 16),
51946 => conv_std_logic_vector(47268, 16),
51947 => conv_std_logic_vector(47470, 16),
51948 => conv_std_logic_vector(47672, 16),
51949 => conv_std_logic_vector(47874, 16),
51950 => conv_std_logic_vector(48076, 16),
51951 => conv_std_logic_vector(48278, 16),
51952 => conv_std_logic_vector(48480, 16),
51953 => conv_std_logic_vector(48682, 16),
51954 => conv_std_logic_vector(48884, 16),
51955 => conv_std_logic_vector(49086, 16),
51956 => conv_std_logic_vector(49288, 16),
51957 => conv_std_logic_vector(49490, 16),
51958 => conv_std_logic_vector(49692, 16),
51959 => conv_std_logic_vector(49894, 16),
51960 => conv_std_logic_vector(50096, 16),
51961 => conv_std_logic_vector(50298, 16),
51962 => conv_std_logic_vector(50500, 16),
51963 => conv_std_logic_vector(50702, 16),
51964 => conv_std_logic_vector(50904, 16),
51965 => conv_std_logic_vector(51106, 16),
51966 => conv_std_logic_vector(51308, 16),
51967 => conv_std_logic_vector(51510, 16),
51968 => conv_std_logic_vector(0, 16),
51969 => conv_std_logic_vector(203, 16),
51970 => conv_std_logic_vector(406, 16),
51971 => conv_std_logic_vector(609, 16),
51972 => conv_std_logic_vector(812, 16),
51973 => conv_std_logic_vector(1015, 16),
51974 => conv_std_logic_vector(1218, 16),
51975 => conv_std_logic_vector(1421, 16),
51976 => conv_std_logic_vector(1624, 16),
51977 => conv_std_logic_vector(1827, 16),
51978 => conv_std_logic_vector(2030, 16),
51979 => conv_std_logic_vector(2233, 16),
51980 => conv_std_logic_vector(2436, 16),
51981 => conv_std_logic_vector(2639, 16),
51982 => conv_std_logic_vector(2842, 16),
51983 => conv_std_logic_vector(3045, 16),
51984 => conv_std_logic_vector(3248, 16),
51985 => conv_std_logic_vector(3451, 16),
51986 => conv_std_logic_vector(3654, 16),
51987 => conv_std_logic_vector(3857, 16),
51988 => conv_std_logic_vector(4060, 16),
51989 => conv_std_logic_vector(4263, 16),
51990 => conv_std_logic_vector(4466, 16),
51991 => conv_std_logic_vector(4669, 16),
51992 => conv_std_logic_vector(4872, 16),
51993 => conv_std_logic_vector(5075, 16),
51994 => conv_std_logic_vector(5278, 16),
51995 => conv_std_logic_vector(5481, 16),
51996 => conv_std_logic_vector(5684, 16),
51997 => conv_std_logic_vector(5887, 16),
51998 => conv_std_logic_vector(6090, 16),
51999 => conv_std_logic_vector(6293, 16),
52000 => conv_std_logic_vector(6496, 16),
52001 => conv_std_logic_vector(6699, 16),
52002 => conv_std_logic_vector(6902, 16),
52003 => conv_std_logic_vector(7105, 16),
52004 => conv_std_logic_vector(7308, 16),
52005 => conv_std_logic_vector(7511, 16),
52006 => conv_std_logic_vector(7714, 16),
52007 => conv_std_logic_vector(7917, 16),
52008 => conv_std_logic_vector(8120, 16),
52009 => conv_std_logic_vector(8323, 16),
52010 => conv_std_logic_vector(8526, 16),
52011 => conv_std_logic_vector(8729, 16),
52012 => conv_std_logic_vector(8932, 16),
52013 => conv_std_logic_vector(9135, 16),
52014 => conv_std_logic_vector(9338, 16),
52015 => conv_std_logic_vector(9541, 16),
52016 => conv_std_logic_vector(9744, 16),
52017 => conv_std_logic_vector(9947, 16),
52018 => conv_std_logic_vector(10150, 16),
52019 => conv_std_logic_vector(10353, 16),
52020 => conv_std_logic_vector(10556, 16),
52021 => conv_std_logic_vector(10759, 16),
52022 => conv_std_logic_vector(10962, 16),
52023 => conv_std_logic_vector(11165, 16),
52024 => conv_std_logic_vector(11368, 16),
52025 => conv_std_logic_vector(11571, 16),
52026 => conv_std_logic_vector(11774, 16),
52027 => conv_std_logic_vector(11977, 16),
52028 => conv_std_logic_vector(12180, 16),
52029 => conv_std_logic_vector(12383, 16),
52030 => conv_std_logic_vector(12586, 16),
52031 => conv_std_logic_vector(12789, 16),
52032 => conv_std_logic_vector(12992, 16),
52033 => conv_std_logic_vector(13195, 16),
52034 => conv_std_logic_vector(13398, 16),
52035 => conv_std_logic_vector(13601, 16),
52036 => conv_std_logic_vector(13804, 16),
52037 => conv_std_logic_vector(14007, 16),
52038 => conv_std_logic_vector(14210, 16),
52039 => conv_std_logic_vector(14413, 16),
52040 => conv_std_logic_vector(14616, 16),
52041 => conv_std_logic_vector(14819, 16),
52042 => conv_std_logic_vector(15022, 16),
52043 => conv_std_logic_vector(15225, 16),
52044 => conv_std_logic_vector(15428, 16),
52045 => conv_std_logic_vector(15631, 16),
52046 => conv_std_logic_vector(15834, 16),
52047 => conv_std_logic_vector(16037, 16),
52048 => conv_std_logic_vector(16240, 16),
52049 => conv_std_logic_vector(16443, 16),
52050 => conv_std_logic_vector(16646, 16),
52051 => conv_std_logic_vector(16849, 16),
52052 => conv_std_logic_vector(17052, 16),
52053 => conv_std_logic_vector(17255, 16),
52054 => conv_std_logic_vector(17458, 16),
52055 => conv_std_logic_vector(17661, 16),
52056 => conv_std_logic_vector(17864, 16),
52057 => conv_std_logic_vector(18067, 16),
52058 => conv_std_logic_vector(18270, 16),
52059 => conv_std_logic_vector(18473, 16),
52060 => conv_std_logic_vector(18676, 16),
52061 => conv_std_logic_vector(18879, 16),
52062 => conv_std_logic_vector(19082, 16),
52063 => conv_std_logic_vector(19285, 16),
52064 => conv_std_logic_vector(19488, 16),
52065 => conv_std_logic_vector(19691, 16),
52066 => conv_std_logic_vector(19894, 16),
52067 => conv_std_logic_vector(20097, 16),
52068 => conv_std_logic_vector(20300, 16),
52069 => conv_std_logic_vector(20503, 16),
52070 => conv_std_logic_vector(20706, 16),
52071 => conv_std_logic_vector(20909, 16),
52072 => conv_std_logic_vector(21112, 16),
52073 => conv_std_logic_vector(21315, 16),
52074 => conv_std_logic_vector(21518, 16),
52075 => conv_std_logic_vector(21721, 16),
52076 => conv_std_logic_vector(21924, 16),
52077 => conv_std_logic_vector(22127, 16),
52078 => conv_std_logic_vector(22330, 16),
52079 => conv_std_logic_vector(22533, 16),
52080 => conv_std_logic_vector(22736, 16),
52081 => conv_std_logic_vector(22939, 16),
52082 => conv_std_logic_vector(23142, 16),
52083 => conv_std_logic_vector(23345, 16),
52084 => conv_std_logic_vector(23548, 16),
52085 => conv_std_logic_vector(23751, 16),
52086 => conv_std_logic_vector(23954, 16),
52087 => conv_std_logic_vector(24157, 16),
52088 => conv_std_logic_vector(24360, 16),
52089 => conv_std_logic_vector(24563, 16),
52090 => conv_std_logic_vector(24766, 16),
52091 => conv_std_logic_vector(24969, 16),
52092 => conv_std_logic_vector(25172, 16),
52093 => conv_std_logic_vector(25375, 16),
52094 => conv_std_logic_vector(25578, 16),
52095 => conv_std_logic_vector(25781, 16),
52096 => conv_std_logic_vector(25984, 16),
52097 => conv_std_logic_vector(26187, 16),
52098 => conv_std_logic_vector(26390, 16),
52099 => conv_std_logic_vector(26593, 16),
52100 => conv_std_logic_vector(26796, 16),
52101 => conv_std_logic_vector(26999, 16),
52102 => conv_std_logic_vector(27202, 16),
52103 => conv_std_logic_vector(27405, 16),
52104 => conv_std_logic_vector(27608, 16),
52105 => conv_std_logic_vector(27811, 16),
52106 => conv_std_logic_vector(28014, 16),
52107 => conv_std_logic_vector(28217, 16),
52108 => conv_std_logic_vector(28420, 16),
52109 => conv_std_logic_vector(28623, 16),
52110 => conv_std_logic_vector(28826, 16),
52111 => conv_std_logic_vector(29029, 16),
52112 => conv_std_logic_vector(29232, 16),
52113 => conv_std_logic_vector(29435, 16),
52114 => conv_std_logic_vector(29638, 16),
52115 => conv_std_logic_vector(29841, 16),
52116 => conv_std_logic_vector(30044, 16),
52117 => conv_std_logic_vector(30247, 16),
52118 => conv_std_logic_vector(30450, 16),
52119 => conv_std_logic_vector(30653, 16),
52120 => conv_std_logic_vector(30856, 16),
52121 => conv_std_logic_vector(31059, 16),
52122 => conv_std_logic_vector(31262, 16),
52123 => conv_std_logic_vector(31465, 16),
52124 => conv_std_logic_vector(31668, 16),
52125 => conv_std_logic_vector(31871, 16),
52126 => conv_std_logic_vector(32074, 16),
52127 => conv_std_logic_vector(32277, 16),
52128 => conv_std_logic_vector(32480, 16),
52129 => conv_std_logic_vector(32683, 16),
52130 => conv_std_logic_vector(32886, 16),
52131 => conv_std_logic_vector(33089, 16),
52132 => conv_std_logic_vector(33292, 16),
52133 => conv_std_logic_vector(33495, 16),
52134 => conv_std_logic_vector(33698, 16),
52135 => conv_std_logic_vector(33901, 16),
52136 => conv_std_logic_vector(34104, 16),
52137 => conv_std_logic_vector(34307, 16),
52138 => conv_std_logic_vector(34510, 16),
52139 => conv_std_logic_vector(34713, 16),
52140 => conv_std_logic_vector(34916, 16),
52141 => conv_std_logic_vector(35119, 16),
52142 => conv_std_logic_vector(35322, 16),
52143 => conv_std_logic_vector(35525, 16),
52144 => conv_std_logic_vector(35728, 16),
52145 => conv_std_logic_vector(35931, 16),
52146 => conv_std_logic_vector(36134, 16),
52147 => conv_std_logic_vector(36337, 16),
52148 => conv_std_logic_vector(36540, 16),
52149 => conv_std_logic_vector(36743, 16),
52150 => conv_std_logic_vector(36946, 16),
52151 => conv_std_logic_vector(37149, 16),
52152 => conv_std_logic_vector(37352, 16),
52153 => conv_std_logic_vector(37555, 16),
52154 => conv_std_logic_vector(37758, 16),
52155 => conv_std_logic_vector(37961, 16),
52156 => conv_std_logic_vector(38164, 16),
52157 => conv_std_logic_vector(38367, 16),
52158 => conv_std_logic_vector(38570, 16),
52159 => conv_std_logic_vector(38773, 16),
52160 => conv_std_logic_vector(38976, 16),
52161 => conv_std_logic_vector(39179, 16),
52162 => conv_std_logic_vector(39382, 16),
52163 => conv_std_logic_vector(39585, 16),
52164 => conv_std_logic_vector(39788, 16),
52165 => conv_std_logic_vector(39991, 16),
52166 => conv_std_logic_vector(40194, 16),
52167 => conv_std_logic_vector(40397, 16),
52168 => conv_std_logic_vector(40600, 16),
52169 => conv_std_logic_vector(40803, 16),
52170 => conv_std_logic_vector(41006, 16),
52171 => conv_std_logic_vector(41209, 16),
52172 => conv_std_logic_vector(41412, 16),
52173 => conv_std_logic_vector(41615, 16),
52174 => conv_std_logic_vector(41818, 16),
52175 => conv_std_logic_vector(42021, 16),
52176 => conv_std_logic_vector(42224, 16),
52177 => conv_std_logic_vector(42427, 16),
52178 => conv_std_logic_vector(42630, 16),
52179 => conv_std_logic_vector(42833, 16),
52180 => conv_std_logic_vector(43036, 16),
52181 => conv_std_logic_vector(43239, 16),
52182 => conv_std_logic_vector(43442, 16),
52183 => conv_std_logic_vector(43645, 16),
52184 => conv_std_logic_vector(43848, 16),
52185 => conv_std_logic_vector(44051, 16),
52186 => conv_std_logic_vector(44254, 16),
52187 => conv_std_logic_vector(44457, 16),
52188 => conv_std_logic_vector(44660, 16),
52189 => conv_std_logic_vector(44863, 16),
52190 => conv_std_logic_vector(45066, 16),
52191 => conv_std_logic_vector(45269, 16),
52192 => conv_std_logic_vector(45472, 16),
52193 => conv_std_logic_vector(45675, 16),
52194 => conv_std_logic_vector(45878, 16),
52195 => conv_std_logic_vector(46081, 16),
52196 => conv_std_logic_vector(46284, 16),
52197 => conv_std_logic_vector(46487, 16),
52198 => conv_std_logic_vector(46690, 16),
52199 => conv_std_logic_vector(46893, 16),
52200 => conv_std_logic_vector(47096, 16),
52201 => conv_std_logic_vector(47299, 16),
52202 => conv_std_logic_vector(47502, 16),
52203 => conv_std_logic_vector(47705, 16),
52204 => conv_std_logic_vector(47908, 16),
52205 => conv_std_logic_vector(48111, 16),
52206 => conv_std_logic_vector(48314, 16),
52207 => conv_std_logic_vector(48517, 16),
52208 => conv_std_logic_vector(48720, 16),
52209 => conv_std_logic_vector(48923, 16),
52210 => conv_std_logic_vector(49126, 16),
52211 => conv_std_logic_vector(49329, 16),
52212 => conv_std_logic_vector(49532, 16),
52213 => conv_std_logic_vector(49735, 16),
52214 => conv_std_logic_vector(49938, 16),
52215 => conv_std_logic_vector(50141, 16),
52216 => conv_std_logic_vector(50344, 16),
52217 => conv_std_logic_vector(50547, 16),
52218 => conv_std_logic_vector(50750, 16),
52219 => conv_std_logic_vector(50953, 16),
52220 => conv_std_logic_vector(51156, 16),
52221 => conv_std_logic_vector(51359, 16),
52222 => conv_std_logic_vector(51562, 16),
52223 => conv_std_logic_vector(51765, 16),
52224 => conv_std_logic_vector(0, 16),
52225 => conv_std_logic_vector(204, 16),
52226 => conv_std_logic_vector(408, 16),
52227 => conv_std_logic_vector(612, 16),
52228 => conv_std_logic_vector(816, 16),
52229 => conv_std_logic_vector(1020, 16),
52230 => conv_std_logic_vector(1224, 16),
52231 => conv_std_logic_vector(1428, 16),
52232 => conv_std_logic_vector(1632, 16),
52233 => conv_std_logic_vector(1836, 16),
52234 => conv_std_logic_vector(2040, 16),
52235 => conv_std_logic_vector(2244, 16),
52236 => conv_std_logic_vector(2448, 16),
52237 => conv_std_logic_vector(2652, 16),
52238 => conv_std_logic_vector(2856, 16),
52239 => conv_std_logic_vector(3060, 16),
52240 => conv_std_logic_vector(3264, 16),
52241 => conv_std_logic_vector(3468, 16),
52242 => conv_std_logic_vector(3672, 16),
52243 => conv_std_logic_vector(3876, 16),
52244 => conv_std_logic_vector(4080, 16),
52245 => conv_std_logic_vector(4284, 16),
52246 => conv_std_logic_vector(4488, 16),
52247 => conv_std_logic_vector(4692, 16),
52248 => conv_std_logic_vector(4896, 16),
52249 => conv_std_logic_vector(5100, 16),
52250 => conv_std_logic_vector(5304, 16),
52251 => conv_std_logic_vector(5508, 16),
52252 => conv_std_logic_vector(5712, 16),
52253 => conv_std_logic_vector(5916, 16),
52254 => conv_std_logic_vector(6120, 16),
52255 => conv_std_logic_vector(6324, 16),
52256 => conv_std_logic_vector(6528, 16),
52257 => conv_std_logic_vector(6732, 16),
52258 => conv_std_logic_vector(6936, 16),
52259 => conv_std_logic_vector(7140, 16),
52260 => conv_std_logic_vector(7344, 16),
52261 => conv_std_logic_vector(7548, 16),
52262 => conv_std_logic_vector(7752, 16),
52263 => conv_std_logic_vector(7956, 16),
52264 => conv_std_logic_vector(8160, 16),
52265 => conv_std_logic_vector(8364, 16),
52266 => conv_std_logic_vector(8568, 16),
52267 => conv_std_logic_vector(8772, 16),
52268 => conv_std_logic_vector(8976, 16),
52269 => conv_std_logic_vector(9180, 16),
52270 => conv_std_logic_vector(9384, 16),
52271 => conv_std_logic_vector(9588, 16),
52272 => conv_std_logic_vector(9792, 16),
52273 => conv_std_logic_vector(9996, 16),
52274 => conv_std_logic_vector(10200, 16),
52275 => conv_std_logic_vector(10404, 16),
52276 => conv_std_logic_vector(10608, 16),
52277 => conv_std_logic_vector(10812, 16),
52278 => conv_std_logic_vector(11016, 16),
52279 => conv_std_logic_vector(11220, 16),
52280 => conv_std_logic_vector(11424, 16),
52281 => conv_std_logic_vector(11628, 16),
52282 => conv_std_logic_vector(11832, 16),
52283 => conv_std_logic_vector(12036, 16),
52284 => conv_std_logic_vector(12240, 16),
52285 => conv_std_logic_vector(12444, 16),
52286 => conv_std_logic_vector(12648, 16),
52287 => conv_std_logic_vector(12852, 16),
52288 => conv_std_logic_vector(13056, 16),
52289 => conv_std_logic_vector(13260, 16),
52290 => conv_std_logic_vector(13464, 16),
52291 => conv_std_logic_vector(13668, 16),
52292 => conv_std_logic_vector(13872, 16),
52293 => conv_std_logic_vector(14076, 16),
52294 => conv_std_logic_vector(14280, 16),
52295 => conv_std_logic_vector(14484, 16),
52296 => conv_std_logic_vector(14688, 16),
52297 => conv_std_logic_vector(14892, 16),
52298 => conv_std_logic_vector(15096, 16),
52299 => conv_std_logic_vector(15300, 16),
52300 => conv_std_logic_vector(15504, 16),
52301 => conv_std_logic_vector(15708, 16),
52302 => conv_std_logic_vector(15912, 16),
52303 => conv_std_logic_vector(16116, 16),
52304 => conv_std_logic_vector(16320, 16),
52305 => conv_std_logic_vector(16524, 16),
52306 => conv_std_logic_vector(16728, 16),
52307 => conv_std_logic_vector(16932, 16),
52308 => conv_std_logic_vector(17136, 16),
52309 => conv_std_logic_vector(17340, 16),
52310 => conv_std_logic_vector(17544, 16),
52311 => conv_std_logic_vector(17748, 16),
52312 => conv_std_logic_vector(17952, 16),
52313 => conv_std_logic_vector(18156, 16),
52314 => conv_std_logic_vector(18360, 16),
52315 => conv_std_logic_vector(18564, 16),
52316 => conv_std_logic_vector(18768, 16),
52317 => conv_std_logic_vector(18972, 16),
52318 => conv_std_logic_vector(19176, 16),
52319 => conv_std_logic_vector(19380, 16),
52320 => conv_std_logic_vector(19584, 16),
52321 => conv_std_logic_vector(19788, 16),
52322 => conv_std_logic_vector(19992, 16),
52323 => conv_std_logic_vector(20196, 16),
52324 => conv_std_logic_vector(20400, 16),
52325 => conv_std_logic_vector(20604, 16),
52326 => conv_std_logic_vector(20808, 16),
52327 => conv_std_logic_vector(21012, 16),
52328 => conv_std_logic_vector(21216, 16),
52329 => conv_std_logic_vector(21420, 16),
52330 => conv_std_logic_vector(21624, 16),
52331 => conv_std_logic_vector(21828, 16),
52332 => conv_std_logic_vector(22032, 16),
52333 => conv_std_logic_vector(22236, 16),
52334 => conv_std_logic_vector(22440, 16),
52335 => conv_std_logic_vector(22644, 16),
52336 => conv_std_logic_vector(22848, 16),
52337 => conv_std_logic_vector(23052, 16),
52338 => conv_std_logic_vector(23256, 16),
52339 => conv_std_logic_vector(23460, 16),
52340 => conv_std_logic_vector(23664, 16),
52341 => conv_std_logic_vector(23868, 16),
52342 => conv_std_logic_vector(24072, 16),
52343 => conv_std_logic_vector(24276, 16),
52344 => conv_std_logic_vector(24480, 16),
52345 => conv_std_logic_vector(24684, 16),
52346 => conv_std_logic_vector(24888, 16),
52347 => conv_std_logic_vector(25092, 16),
52348 => conv_std_logic_vector(25296, 16),
52349 => conv_std_logic_vector(25500, 16),
52350 => conv_std_logic_vector(25704, 16),
52351 => conv_std_logic_vector(25908, 16),
52352 => conv_std_logic_vector(26112, 16),
52353 => conv_std_logic_vector(26316, 16),
52354 => conv_std_logic_vector(26520, 16),
52355 => conv_std_logic_vector(26724, 16),
52356 => conv_std_logic_vector(26928, 16),
52357 => conv_std_logic_vector(27132, 16),
52358 => conv_std_logic_vector(27336, 16),
52359 => conv_std_logic_vector(27540, 16),
52360 => conv_std_logic_vector(27744, 16),
52361 => conv_std_logic_vector(27948, 16),
52362 => conv_std_logic_vector(28152, 16),
52363 => conv_std_logic_vector(28356, 16),
52364 => conv_std_logic_vector(28560, 16),
52365 => conv_std_logic_vector(28764, 16),
52366 => conv_std_logic_vector(28968, 16),
52367 => conv_std_logic_vector(29172, 16),
52368 => conv_std_logic_vector(29376, 16),
52369 => conv_std_logic_vector(29580, 16),
52370 => conv_std_logic_vector(29784, 16),
52371 => conv_std_logic_vector(29988, 16),
52372 => conv_std_logic_vector(30192, 16),
52373 => conv_std_logic_vector(30396, 16),
52374 => conv_std_logic_vector(30600, 16),
52375 => conv_std_logic_vector(30804, 16),
52376 => conv_std_logic_vector(31008, 16),
52377 => conv_std_logic_vector(31212, 16),
52378 => conv_std_logic_vector(31416, 16),
52379 => conv_std_logic_vector(31620, 16),
52380 => conv_std_logic_vector(31824, 16),
52381 => conv_std_logic_vector(32028, 16),
52382 => conv_std_logic_vector(32232, 16),
52383 => conv_std_logic_vector(32436, 16),
52384 => conv_std_logic_vector(32640, 16),
52385 => conv_std_logic_vector(32844, 16),
52386 => conv_std_logic_vector(33048, 16),
52387 => conv_std_logic_vector(33252, 16),
52388 => conv_std_logic_vector(33456, 16),
52389 => conv_std_logic_vector(33660, 16),
52390 => conv_std_logic_vector(33864, 16),
52391 => conv_std_logic_vector(34068, 16),
52392 => conv_std_logic_vector(34272, 16),
52393 => conv_std_logic_vector(34476, 16),
52394 => conv_std_logic_vector(34680, 16),
52395 => conv_std_logic_vector(34884, 16),
52396 => conv_std_logic_vector(35088, 16),
52397 => conv_std_logic_vector(35292, 16),
52398 => conv_std_logic_vector(35496, 16),
52399 => conv_std_logic_vector(35700, 16),
52400 => conv_std_logic_vector(35904, 16),
52401 => conv_std_logic_vector(36108, 16),
52402 => conv_std_logic_vector(36312, 16),
52403 => conv_std_logic_vector(36516, 16),
52404 => conv_std_logic_vector(36720, 16),
52405 => conv_std_logic_vector(36924, 16),
52406 => conv_std_logic_vector(37128, 16),
52407 => conv_std_logic_vector(37332, 16),
52408 => conv_std_logic_vector(37536, 16),
52409 => conv_std_logic_vector(37740, 16),
52410 => conv_std_logic_vector(37944, 16),
52411 => conv_std_logic_vector(38148, 16),
52412 => conv_std_logic_vector(38352, 16),
52413 => conv_std_logic_vector(38556, 16),
52414 => conv_std_logic_vector(38760, 16),
52415 => conv_std_logic_vector(38964, 16),
52416 => conv_std_logic_vector(39168, 16),
52417 => conv_std_logic_vector(39372, 16),
52418 => conv_std_logic_vector(39576, 16),
52419 => conv_std_logic_vector(39780, 16),
52420 => conv_std_logic_vector(39984, 16),
52421 => conv_std_logic_vector(40188, 16),
52422 => conv_std_logic_vector(40392, 16),
52423 => conv_std_logic_vector(40596, 16),
52424 => conv_std_logic_vector(40800, 16),
52425 => conv_std_logic_vector(41004, 16),
52426 => conv_std_logic_vector(41208, 16),
52427 => conv_std_logic_vector(41412, 16),
52428 => conv_std_logic_vector(41616, 16),
52429 => conv_std_logic_vector(41820, 16),
52430 => conv_std_logic_vector(42024, 16),
52431 => conv_std_logic_vector(42228, 16),
52432 => conv_std_logic_vector(42432, 16),
52433 => conv_std_logic_vector(42636, 16),
52434 => conv_std_logic_vector(42840, 16),
52435 => conv_std_logic_vector(43044, 16),
52436 => conv_std_logic_vector(43248, 16),
52437 => conv_std_logic_vector(43452, 16),
52438 => conv_std_logic_vector(43656, 16),
52439 => conv_std_logic_vector(43860, 16),
52440 => conv_std_logic_vector(44064, 16),
52441 => conv_std_logic_vector(44268, 16),
52442 => conv_std_logic_vector(44472, 16),
52443 => conv_std_logic_vector(44676, 16),
52444 => conv_std_logic_vector(44880, 16),
52445 => conv_std_logic_vector(45084, 16),
52446 => conv_std_logic_vector(45288, 16),
52447 => conv_std_logic_vector(45492, 16),
52448 => conv_std_logic_vector(45696, 16),
52449 => conv_std_logic_vector(45900, 16),
52450 => conv_std_logic_vector(46104, 16),
52451 => conv_std_logic_vector(46308, 16),
52452 => conv_std_logic_vector(46512, 16),
52453 => conv_std_logic_vector(46716, 16),
52454 => conv_std_logic_vector(46920, 16),
52455 => conv_std_logic_vector(47124, 16),
52456 => conv_std_logic_vector(47328, 16),
52457 => conv_std_logic_vector(47532, 16),
52458 => conv_std_logic_vector(47736, 16),
52459 => conv_std_logic_vector(47940, 16),
52460 => conv_std_logic_vector(48144, 16),
52461 => conv_std_logic_vector(48348, 16),
52462 => conv_std_logic_vector(48552, 16),
52463 => conv_std_logic_vector(48756, 16),
52464 => conv_std_logic_vector(48960, 16),
52465 => conv_std_logic_vector(49164, 16),
52466 => conv_std_logic_vector(49368, 16),
52467 => conv_std_logic_vector(49572, 16),
52468 => conv_std_logic_vector(49776, 16),
52469 => conv_std_logic_vector(49980, 16),
52470 => conv_std_logic_vector(50184, 16),
52471 => conv_std_logic_vector(50388, 16),
52472 => conv_std_logic_vector(50592, 16),
52473 => conv_std_logic_vector(50796, 16),
52474 => conv_std_logic_vector(51000, 16),
52475 => conv_std_logic_vector(51204, 16),
52476 => conv_std_logic_vector(51408, 16),
52477 => conv_std_logic_vector(51612, 16),
52478 => conv_std_logic_vector(51816, 16),
52479 => conv_std_logic_vector(52020, 16),
52480 => conv_std_logic_vector(0, 16),
52481 => conv_std_logic_vector(205, 16),
52482 => conv_std_logic_vector(410, 16),
52483 => conv_std_logic_vector(615, 16),
52484 => conv_std_logic_vector(820, 16),
52485 => conv_std_logic_vector(1025, 16),
52486 => conv_std_logic_vector(1230, 16),
52487 => conv_std_logic_vector(1435, 16),
52488 => conv_std_logic_vector(1640, 16),
52489 => conv_std_logic_vector(1845, 16),
52490 => conv_std_logic_vector(2050, 16),
52491 => conv_std_logic_vector(2255, 16),
52492 => conv_std_logic_vector(2460, 16),
52493 => conv_std_logic_vector(2665, 16),
52494 => conv_std_logic_vector(2870, 16),
52495 => conv_std_logic_vector(3075, 16),
52496 => conv_std_logic_vector(3280, 16),
52497 => conv_std_logic_vector(3485, 16),
52498 => conv_std_logic_vector(3690, 16),
52499 => conv_std_logic_vector(3895, 16),
52500 => conv_std_logic_vector(4100, 16),
52501 => conv_std_logic_vector(4305, 16),
52502 => conv_std_logic_vector(4510, 16),
52503 => conv_std_logic_vector(4715, 16),
52504 => conv_std_logic_vector(4920, 16),
52505 => conv_std_logic_vector(5125, 16),
52506 => conv_std_logic_vector(5330, 16),
52507 => conv_std_logic_vector(5535, 16),
52508 => conv_std_logic_vector(5740, 16),
52509 => conv_std_logic_vector(5945, 16),
52510 => conv_std_logic_vector(6150, 16),
52511 => conv_std_logic_vector(6355, 16),
52512 => conv_std_logic_vector(6560, 16),
52513 => conv_std_logic_vector(6765, 16),
52514 => conv_std_logic_vector(6970, 16),
52515 => conv_std_logic_vector(7175, 16),
52516 => conv_std_logic_vector(7380, 16),
52517 => conv_std_logic_vector(7585, 16),
52518 => conv_std_logic_vector(7790, 16),
52519 => conv_std_logic_vector(7995, 16),
52520 => conv_std_logic_vector(8200, 16),
52521 => conv_std_logic_vector(8405, 16),
52522 => conv_std_logic_vector(8610, 16),
52523 => conv_std_logic_vector(8815, 16),
52524 => conv_std_logic_vector(9020, 16),
52525 => conv_std_logic_vector(9225, 16),
52526 => conv_std_logic_vector(9430, 16),
52527 => conv_std_logic_vector(9635, 16),
52528 => conv_std_logic_vector(9840, 16),
52529 => conv_std_logic_vector(10045, 16),
52530 => conv_std_logic_vector(10250, 16),
52531 => conv_std_logic_vector(10455, 16),
52532 => conv_std_logic_vector(10660, 16),
52533 => conv_std_logic_vector(10865, 16),
52534 => conv_std_logic_vector(11070, 16),
52535 => conv_std_logic_vector(11275, 16),
52536 => conv_std_logic_vector(11480, 16),
52537 => conv_std_logic_vector(11685, 16),
52538 => conv_std_logic_vector(11890, 16),
52539 => conv_std_logic_vector(12095, 16),
52540 => conv_std_logic_vector(12300, 16),
52541 => conv_std_logic_vector(12505, 16),
52542 => conv_std_logic_vector(12710, 16),
52543 => conv_std_logic_vector(12915, 16),
52544 => conv_std_logic_vector(13120, 16),
52545 => conv_std_logic_vector(13325, 16),
52546 => conv_std_logic_vector(13530, 16),
52547 => conv_std_logic_vector(13735, 16),
52548 => conv_std_logic_vector(13940, 16),
52549 => conv_std_logic_vector(14145, 16),
52550 => conv_std_logic_vector(14350, 16),
52551 => conv_std_logic_vector(14555, 16),
52552 => conv_std_logic_vector(14760, 16),
52553 => conv_std_logic_vector(14965, 16),
52554 => conv_std_logic_vector(15170, 16),
52555 => conv_std_logic_vector(15375, 16),
52556 => conv_std_logic_vector(15580, 16),
52557 => conv_std_logic_vector(15785, 16),
52558 => conv_std_logic_vector(15990, 16),
52559 => conv_std_logic_vector(16195, 16),
52560 => conv_std_logic_vector(16400, 16),
52561 => conv_std_logic_vector(16605, 16),
52562 => conv_std_logic_vector(16810, 16),
52563 => conv_std_logic_vector(17015, 16),
52564 => conv_std_logic_vector(17220, 16),
52565 => conv_std_logic_vector(17425, 16),
52566 => conv_std_logic_vector(17630, 16),
52567 => conv_std_logic_vector(17835, 16),
52568 => conv_std_logic_vector(18040, 16),
52569 => conv_std_logic_vector(18245, 16),
52570 => conv_std_logic_vector(18450, 16),
52571 => conv_std_logic_vector(18655, 16),
52572 => conv_std_logic_vector(18860, 16),
52573 => conv_std_logic_vector(19065, 16),
52574 => conv_std_logic_vector(19270, 16),
52575 => conv_std_logic_vector(19475, 16),
52576 => conv_std_logic_vector(19680, 16),
52577 => conv_std_logic_vector(19885, 16),
52578 => conv_std_logic_vector(20090, 16),
52579 => conv_std_logic_vector(20295, 16),
52580 => conv_std_logic_vector(20500, 16),
52581 => conv_std_logic_vector(20705, 16),
52582 => conv_std_logic_vector(20910, 16),
52583 => conv_std_logic_vector(21115, 16),
52584 => conv_std_logic_vector(21320, 16),
52585 => conv_std_logic_vector(21525, 16),
52586 => conv_std_logic_vector(21730, 16),
52587 => conv_std_logic_vector(21935, 16),
52588 => conv_std_logic_vector(22140, 16),
52589 => conv_std_logic_vector(22345, 16),
52590 => conv_std_logic_vector(22550, 16),
52591 => conv_std_logic_vector(22755, 16),
52592 => conv_std_logic_vector(22960, 16),
52593 => conv_std_logic_vector(23165, 16),
52594 => conv_std_logic_vector(23370, 16),
52595 => conv_std_logic_vector(23575, 16),
52596 => conv_std_logic_vector(23780, 16),
52597 => conv_std_logic_vector(23985, 16),
52598 => conv_std_logic_vector(24190, 16),
52599 => conv_std_logic_vector(24395, 16),
52600 => conv_std_logic_vector(24600, 16),
52601 => conv_std_logic_vector(24805, 16),
52602 => conv_std_logic_vector(25010, 16),
52603 => conv_std_logic_vector(25215, 16),
52604 => conv_std_logic_vector(25420, 16),
52605 => conv_std_logic_vector(25625, 16),
52606 => conv_std_logic_vector(25830, 16),
52607 => conv_std_logic_vector(26035, 16),
52608 => conv_std_logic_vector(26240, 16),
52609 => conv_std_logic_vector(26445, 16),
52610 => conv_std_logic_vector(26650, 16),
52611 => conv_std_logic_vector(26855, 16),
52612 => conv_std_logic_vector(27060, 16),
52613 => conv_std_logic_vector(27265, 16),
52614 => conv_std_logic_vector(27470, 16),
52615 => conv_std_logic_vector(27675, 16),
52616 => conv_std_logic_vector(27880, 16),
52617 => conv_std_logic_vector(28085, 16),
52618 => conv_std_logic_vector(28290, 16),
52619 => conv_std_logic_vector(28495, 16),
52620 => conv_std_logic_vector(28700, 16),
52621 => conv_std_logic_vector(28905, 16),
52622 => conv_std_logic_vector(29110, 16),
52623 => conv_std_logic_vector(29315, 16),
52624 => conv_std_logic_vector(29520, 16),
52625 => conv_std_logic_vector(29725, 16),
52626 => conv_std_logic_vector(29930, 16),
52627 => conv_std_logic_vector(30135, 16),
52628 => conv_std_logic_vector(30340, 16),
52629 => conv_std_logic_vector(30545, 16),
52630 => conv_std_logic_vector(30750, 16),
52631 => conv_std_logic_vector(30955, 16),
52632 => conv_std_logic_vector(31160, 16),
52633 => conv_std_logic_vector(31365, 16),
52634 => conv_std_logic_vector(31570, 16),
52635 => conv_std_logic_vector(31775, 16),
52636 => conv_std_logic_vector(31980, 16),
52637 => conv_std_logic_vector(32185, 16),
52638 => conv_std_logic_vector(32390, 16),
52639 => conv_std_logic_vector(32595, 16),
52640 => conv_std_logic_vector(32800, 16),
52641 => conv_std_logic_vector(33005, 16),
52642 => conv_std_logic_vector(33210, 16),
52643 => conv_std_logic_vector(33415, 16),
52644 => conv_std_logic_vector(33620, 16),
52645 => conv_std_logic_vector(33825, 16),
52646 => conv_std_logic_vector(34030, 16),
52647 => conv_std_logic_vector(34235, 16),
52648 => conv_std_logic_vector(34440, 16),
52649 => conv_std_logic_vector(34645, 16),
52650 => conv_std_logic_vector(34850, 16),
52651 => conv_std_logic_vector(35055, 16),
52652 => conv_std_logic_vector(35260, 16),
52653 => conv_std_logic_vector(35465, 16),
52654 => conv_std_logic_vector(35670, 16),
52655 => conv_std_logic_vector(35875, 16),
52656 => conv_std_logic_vector(36080, 16),
52657 => conv_std_logic_vector(36285, 16),
52658 => conv_std_logic_vector(36490, 16),
52659 => conv_std_logic_vector(36695, 16),
52660 => conv_std_logic_vector(36900, 16),
52661 => conv_std_logic_vector(37105, 16),
52662 => conv_std_logic_vector(37310, 16),
52663 => conv_std_logic_vector(37515, 16),
52664 => conv_std_logic_vector(37720, 16),
52665 => conv_std_logic_vector(37925, 16),
52666 => conv_std_logic_vector(38130, 16),
52667 => conv_std_logic_vector(38335, 16),
52668 => conv_std_logic_vector(38540, 16),
52669 => conv_std_logic_vector(38745, 16),
52670 => conv_std_logic_vector(38950, 16),
52671 => conv_std_logic_vector(39155, 16),
52672 => conv_std_logic_vector(39360, 16),
52673 => conv_std_logic_vector(39565, 16),
52674 => conv_std_logic_vector(39770, 16),
52675 => conv_std_logic_vector(39975, 16),
52676 => conv_std_logic_vector(40180, 16),
52677 => conv_std_logic_vector(40385, 16),
52678 => conv_std_logic_vector(40590, 16),
52679 => conv_std_logic_vector(40795, 16),
52680 => conv_std_logic_vector(41000, 16),
52681 => conv_std_logic_vector(41205, 16),
52682 => conv_std_logic_vector(41410, 16),
52683 => conv_std_logic_vector(41615, 16),
52684 => conv_std_logic_vector(41820, 16),
52685 => conv_std_logic_vector(42025, 16),
52686 => conv_std_logic_vector(42230, 16),
52687 => conv_std_logic_vector(42435, 16),
52688 => conv_std_logic_vector(42640, 16),
52689 => conv_std_logic_vector(42845, 16),
52690 => conv_std_logic_vector(43050, 16),
52691 => conv_std_logic_vector(43255, 16),
52692 => conv_std_logic_vector(43460, 16),
52693 => conv_std_logic_vector(43665, 16),
52694 => conv_std_logic_vector(43870, 16),
52695 => conv_std_logic_vector(44075, 16),
52696 => conv_std_logic_vector(44280, 16),
52697 => conv_std_logic_vector(44485, 16),
52698 => conv_std_logic_vector(44690, 16),
52699 => conv_std_logic_vector(44895, 16),
52700 => conv_std_logic_vector(45100, 16),
52701 => conv_std_logic_vector(45305, 16),
52702 => conv_std_logic_vector(45510, 16),
52703 => conv_std_logic_vector(45715, 16),
52704 => conv_std_logic_vector(45920, 16),
52705 => conv_std_logic_vector(46125, 16),
52706 => conv_std_logic_vector(46330, 16),
52707 => conv_std_logic_vector(46535, 16),
52708 => conv_std_logic_vector(46740, 16),
52709 => conv_std_logic_vector(46945, 16),
52710 => conv_std_logic_vector(47150, 16),
52711 => conv_std_logic_vector(47355, 16),
52712 => conv_std_logic_vector(47560, 16),
52713 => conv_std_logic_vector(47765, 16),
52714 => conv_std_logic_vector(47970, 16),
52715 => conv_std_logic_vector(48175, 16),
52716 => conv_std_logic_vector(48380, 16),
52717 => conv_std_logic_vector(48585, 16),
52718 => conv_std_logic_vector(48790, 16),
52719 => conv_std_logic_vector(48995, 16),
52720 => conv_std_logic_vector(49200, 16),
52721 => conv_std_logic_vector(49405, 16),
52722 => conv_std_logic_vector(49610, 16),
52723 => conv_std_logic_vector(49815, 16),
52724 => conv_std_logic_vector(50020, 16),
52725 => conv_std_logic_vector(50225, 16),
52726 => conv_std_logic_vector(50430, 16),
52727 => conv_std_logic_vector(50635, 16),
52728 => conv_std_logic_vector(50840, 16),
52729 => conv_std_logic_vector(51045, 16),
52730 => conv_std_logic_vector(51250, 16),
52731 => conv_std_logic_vector(51455, 16),
52732 => conv_std_logic_vector(51660, 16),
52733 => conv_std_logic_vector(51865, 16),
52734 => conv_std_logic_vector(52070, 16),
52735 => conv_std_logic_vector(52275, 16),
52736 => conv_std_logic_vector(0, 16),
52737 => conv_std_logic_vector(206, 16),
52738 => conv_std_logic_vector(412, 16),
52739 => conv_std_logic_vector(618, 16),
52740 => conv_std_logic_vector(824, 16),
52741 => conv_std_logic_vector(1030, 16),
52742 => conv_std_logic_vector(1236, 16),
52743 => conv_std_logic_vector(1442, 16),
52744 => conv_std_logic_vector(1648, 16),
52745 => conv_std_logic_vector(1854, 16),
52746 => conv_std_logic_vector(2060, 16),
52747 => conv_std_logic_vector(2266, 16),
52748 => conv_std_logic_vector(2472, 16),
52749 => conv_std_logic_vector(2678, 16),
52750 => conv_std_logic_vector(2884, 16),
52751 => conv_std_logic_vector(3090, 16),
52752 => conv_std_logic_vector(3296, 16),
52753 => conv_std_logic_vector(3502, 16),
52754 => conv_std_logic_vector(3708, 16),
52755 => conv_std_logic_vector(3914, 16),
52756 => conv_std_logic_vector(4120, 16),
52757 => conv_std_logic_vector(4326, 16),
52758 => conv_std_logic_vector(4532, 16),
52759 => conv_std_logic_vector(4738, 16),
52760 => conv_std_logic_vector(4944, 16),
52761 => conv_std_logic_vector(5150, 16),
52762 => conv_std_logic_vector(5356, 16),
52763 => conv_std_logic_vector(5562, 16),
52764 => conv_std_logic_vector(5768, 16),
52765 => conv_std_logic_vector(5974, 16),
52766 => conv_std_logic_vector(6180, 16),
52767 => conv_std_logic_vector(6386, 16),
52768 => conv_std_logic_vector(6592, 16),
52769 => conv_std_logic_vector(6798, 16),
52770 => conv_std_logic_vector(7004, 16),
52771 => conv_std_logic_vector(7210, 16),
52772 => conv_std_logic_vector(7416, 16),
52773 => conv_std_logic_vector(7622, 16),
52774 => conv_std_logic_vector(7828, 16),
52775 => conv_std_logic_vector(8034, 16),
52776 => conv_std_logic_vector(8240, 16),
52777 => conv_std_logic_vector(8446, 16),
52778 => conv_std_logic_vector(8652, 16),
52779 => conv_std_logic_vector(8858, 16),
52780 => conv_std_logic_vector(9064, 16),
52781 => conv_std_logic_vector(9270, 16),
52782 => conv_std_logic_vector(9476, 16),
52783 => conv_std_logic_vector(9682, 16),
52784 => conv_std_logic_vector(9888, 16),
52785 => conv_std_logic_vector(10094, 16),
52786 => conv_std_logic_vector(10300, 16),
52787 => conv_std_logic_vector(10506, 16),
52788 => conv_std_logic_vector(10712, 16),
52789 => conv_std_logic_vector(10918, 16),
52790 => conv_std_logic_vector(11124, 16),
52791 => conv_std_logic_vector(11330, 16),
52792 => conv_std_logic_vector(11536, 16),
52793 => conv_std_logic_vector(11742, 16),
52794 => conv_std_logic_vector(11948, 16),
52795 => conv_std_logic_vector(12154, 16),
52796 => conv_std_logic_vector(12360, 16),
52797 => conv_std_logic_vector(12566, 16),
52798 => conv_std_logic_vector(12772, 16),
52799 => conv_std_logic_vector(12978, 16),
52800 => conv_std_logic_vector(13184, 16),
52801 => conv_std_logic_vector(13390, 16),
52802 => conv_std_logic_vector(13596, 16),
52803 => conv_std_logic_vector(13802, 16),
52804 => conv_std_logic_vector(14008, 16),
52805 => conv_std_logic_vector(14214, 16),
52806 => conv_std_logic_vector(14420, 16),
52807 => conv_std_logic_vector(14626, 16),
52808 => conv_std_logic_vector(14832, 16),
52809 => conv_std_logic_vector(15038, 16),
52810 => conv_std_logic_vector(15244, 16),
52811 => conv_std_logic_vector(15450, 16),
52812 => conv_std_logic_vector(15656, 16),
52813 => conv_std_logic_vector(15862, 16),
52814 => conv_std_logic_vector(16068, 16),
52815 => conv_std_logic_vector(16274, 16),
52816 => conv_std_logic_vector(16480, 16),
52817 => conv_std_logic_vector(16686, 16),
52818 => conv_std_logic_vector(16892, 16),
52819 => conv_std_logic_vector(17098, 16),
52820 => conv_std_logic_vector(17304, 16),
52821 => conv_std_logic_vector(17510, 16),
52822 => conv_std_logic_vector(17716, 16),
52823 => conv_std_logic_vector(17922, 16),
52824 => conv_std_logic_vector(18128, 16),
52825 => conv_std_logic_vector(18334, 16),
52826 => conv_std_logic_vector(18540, 16),
52827 => conv_std_logic_vector(18746, 16),
52828 => conv_std_logic_vector(18952, 16),
52829 => conv_std_logic_vector(19158, 16),
52830 => conv_std_logic_vector(19364, 16),
52831 => conv_std_logic_vector(19570, 16),
52832 => conv_std_logic_vector(19776, 16),
52833 => conv_std_logic_vector(19982, 16),
52834 => conv_std_logic_vector(20188, 16),
52835 => conv_std_logic_vector(20394, 16),
52836 => conv_std_logic_vector(20600, 16),
52837 => conv_std_logic_vector(20806, 16),
52838 => conv_std_logic_vector(21012, 16),
52839 => conv_std_logic_vector(21218, 16),
52840 => conv_std_logic_vector(21424, 16),
52841 => conv_std_logic_vector(21630, 16),
52842 => conv_std_logic_vector(21836, 16),
52843 => conv_std_logic_vector(22042, 16),
52844 => conv_std_logic_vector(22248, 16),
52845 => conv_std_logic_vector(22454, 16),
52846 => conv_std_logic_vector(22660, 16),
52847 => conv_std_logic_vector(22866, 16),
52848 => conv_std_logic_vector(23072, 16),
52849 => conv_std_logic_vector(23278, 16),
52850 => conv_std_logic_vector(23484, 16),
52851 => conv_std_logic_vector(23690, 16),
52852 => conv_std_logic_vector(23896, 16),
52853 => conv_std_logic_vector(24102, 16),
52854 => conv_std_logic_vector(24308, 16),
52855 => conv_std_logic_vector(24514, 16),
52856 => conv_std_logic_vector(24720, 16),
52857 => conv_std_logic_vector(24926, 16),
52858 => conv_std_logic_vector(25132, 16),
52859 => conv_std_logic_vector(25338, 16),
52860 => conv_std_logic_vector(25544, 16),
52861 => conv_std_logic_vector(25750, 16),
52862 => conv_std_logic_vector(25956, 16),
52863 => conv_std_logic_vector(26162, 16),
52864 => conv_std_logic_vector(26368, 16),
52865 => conv_std_logic_vector(26574, 16),
52866 => conv_std_logic_vector(26780, 16),
52867 => conv_std_logic_vector(26986, 16),
52868 => conv_std_logic_vector(27192, 16),
52869 => conv_std_logic_vector(27398, 16),
52870 => conv_std_logic_vector(27604, 16),
52871 => conv_std_logic_vector(27810, 16),
52872 => conv_std_logic_vector(28016, 16),
52873 => conv_std_logic_vector(28222, 16),
52874 => conv_std_logic_vector(28428, 16),
52875 => conv_std_logic_vector(28634, 16),
52876 => conv_std_logic_vector(28840, 16),
52877 => conv_std_logic_vector(29046, 16),
52878 => conv_std_logic_vector(29252, 16),
52879 => conv_std_logic_vector(29458, 16),
52880 => conv_std_logic_vector(29664, 16),
52881 => conv_std_logic_vector(29870, 16),
52882 => conv_std_logic_vector(30076, 16),
52883 => conv_std_logic_vector(30282, 16),
52884 => conv_std_logic_vector(30488, 16),
52885 => conv_std_logic_vector(30694, 16),
52886 => conv_std_logic_vector(30900, 16),
52887 => conv_std_logic_vector(31106, 16),
52888 => conv_std_logic_vector(31312, 16),
52889 => conv_std_logic_vector(31518, 16),
52890 => conv_std_logic_vector(31724, 16),
52891 => conv_std_logic_vector(31930, 16),
52892 => conv_std_logic_vector(32136, 16),
52893 => conv_std_logic_vector(32342, 16),
52894 => conv_std_logic_vector(32548, 16),
52895 => conv_std_logic_vector(32754, 16),
52896 => conv_std_logic_vector(32960, 16),
52897 => conv_std_logic_vector(33166, 16),
52898 => conv_std_logic_vector(33372, 16),
52899 => conv_std_logic_vector(33578, 16),
52900 => conv_std_logic_vector(33784, 16),
52901 => conv_std_logic_vector(33990, 16),
52902 => conv_std_logic_vector(34196, 16),
52903 => conv_std_logic_vector(34402, 16),
52904 => conv_std_logic_vector(34608, 16),
52905 => conv_std_logic_vector(34814, 16),
52906 => conv_std_logic_vector(35020, 16),
52907 => conv_std_logic_vector(35226, 16),
52908 => conv_std_logic_vector(35432, 16),
52909 => conv_std_logic_vector(35638, 16),
52910 => conv_std_logic_vector(35844, 16),
52911 => conv_std_logic_vector(36050, 16),
52912 => conv_std_logic_vector(36256, 16),
52913 => conv_std_logic_vector(36462, 16),
52914 => conv_std_logic_vector(36668, 16),
52915 => conv_std_logic_vector(36874, 16),
52916 => conv_std_logic_vector(37080, 16),
52917 => conv_std_logic_vector(37286, 16),
52918 => conv_std_logic_vector(37492, 16),
52919 => conv_std_logic_vector(37698, 16),
52920 => conv_std_logic_vector(37904, 16),
52921 => conv_std_logic_vector(38110, 16),
52922 => conv_std_logic_vector(38316, 16),
52923 => conv_std_logic_vector(38522, 16),
52924 => conv_std_logic_vector(38728, 16),
52925 => conv_std_logic_vector(38934, 16),
52926 => conv_std_logic_vector(39140, 16),
52927 => conv_std_logic_vector(39346, 16),
52928 => conv_std_logic_vector(39552, 16),
52929 => conv_std_logic_vector(39758, 16),
52930 => conv_std_logic_vector(39964, 16),
52931 => conv_std_logic_vector(40170, 16),
52932 => conv_std_logic_vector(40376, 16),
52933 => conv_std_logic_vector(40582, 16),
52934 => conv_std_logic_vector(40788, 16),
52935 => conv_std_logic_vector(40994, 16),
52936 => conv_std_logic_vector(41200, 16),
52937 => conv_std_logic_vector(41406, 16),
52938 => conv_std_logic_vector(41612, 16),
52939 => conv_std_logic_vector(41818, 16),
52940 => conv_std_logic_vector(42024, 16),
52941 => conv_std_logic_vector(42230, 16),
52942 => conv_std_logic_vector(42436, 16),
52943 => conv_std_logic_vector(42642, 16),
52944 => conv_std_logic_vector(42848, 16),
52945 => conv_std_logic_vector(43054, 16),
52946 => conv_std_logic_vector(43260, 16),
52947 => conv_std_logic_vector(43466, 16),
52948 => conv_std_logic_vector(43672, 16),
52949 => conv_std_logic_vector(43878, 16),
52950 => conv_std_logic_vector(44084, 16),
52951 => conv_std_logic_vector(44290, 16),
52952 => conv_std_logic_vector(44496, 16),
52953 => conv_std_logic_vector(44702, 16),
52954 => conv_std_logic_vector(44908, 16),
52955 => conv_std_logic_vector(45114, 16),
52956 => conv_std_logic_vector(45320, 16),
52957 => conv_std_logic_vector(45526, 16),
52958 => conv_std_logic_vector(45732, 16),
52959 => conv_std_logic_vector(45938, 16),
52960 => conv_std_logic_vector(46144, 16),
52961 => conv_std_logic_vector(46350, 16),
52962 => conv_std_logic_vector(46556, 16),
52963 => conv_std_logic_vector(46762, 16),
52964 => conv_std_logic_vector(46968, 16),
52965 => conv_std_logic_vector(47174, 16),
52966 => conv_std_logic_vector(47380, 16),
52967 => conv_std_logic_vector(47586, 16),
52968 => conv_std_logic_vector(47792, 16),
52969 => conv_std_logic_vector(47998, 16),
52970 => conv_std_logic_vector(48204, 16),
52971 => conv_std_logic_vector(48410, 16),
52972 => conv_std_logic_vector(48616, 16),
52973 => conv_std_logic_vector(48822, 16),
52974 => conv_std_logic_vector(49028, 16),
52975 => conv_std_logic_vector(49234, 16),
52976 => conv_std_logic_vector(49440, 16),
52977 => conv_std_logic_vector(49646, 16),
52978 => conv_std_logic_vector(49852, 16),
52979 => conv_std_logic_vector(50058, 16),
52980 => conv_std_logic_vector(50264, 16),
52981 => conv_std_logic_vector(50470, 16),
52982 => conv_std_logic_vector(50676, 16),
52983 => conv_std_logic_vector(50882, 16),
52984 => conv_std_logic_vector(51088, 16),
52985 => conv_std_logic_vector(51294, 16),
52986 => conv_std_logic_vector(51500, 16),
52987 => conv_std_logic_vector(51706, 16),
52988 => conv_std_logic_vector(51912, 16),
52989 => conv_std_logic_vector(52118, 16),
52990 => conv_std_logic_vector(52324, 16),
52991 => conv_std_logic_vector(52530, 16),
52992 => conv_std_logic_vector(0, 16),
52993 => conv_std_logic_vector(207, 16),
52994 => conv_std_logic_vector(414, 16),
52995 => conv_std_logic_vector(621, 16),
52996 => conv_std_logic_vector(828, 16),
52997 => conv_std_logic_vector(1035, 16),
52998 => conv_std_logic_vector(1242, 16),
52999 => conv_std_logic_vector(1449, 16),
53000 => conv_std_logic_vector(1656, 16),
53001 => conv_std_logic_vector(1863, 16),
53002 => conv_std_logic_vector(2070, 16),
53003 => conv_std_logic_vector(2277, 16),
53004 => conv_std_logic_vector(2484, 16),
53005 => conv_std_logic_vector(2691, 16),
53006 => conv_std_logic_vector(2898, 16),
53007 => conv_std_logic_vector(3105, 16),
53008 => conv_std_logic_vector(3312, 16),
53009 => conv_std_logic_vector(3519, 16),
53010 => conv_std_logic_vector(3726, 16),
53011 => conv_std_logic_vector(3933, 16),
53012 => conv_std_logic_vector(4140, 16),
53013 => conv_std_logic_vector(4347, 16),
53014 => conv_std_logic_vector(4554, 16),
53015 => conv_std_logic_vector(4761, 16),
53016 => conv_std_logic_vector(4968, 16),
53017 => conv_std_logic_vector(5175, 16),
53018 => conv_std_logic_vector(5382, 16),
53019 => conv_std_logic_vector(5589, 16),
53020 => conv_std_logic_vector(5796, 16),
53021 => conv_std_logic_vector(6003, 16),
53022 => conv_std_logic_vector(6210, 16),
53023 => conv_std_logic_vector(6417, 16),
53024 => conv_std_logic_vector(6624, 16),
53025 => conv_std_logic_vector(6831, 16),
53026 => conv_std_logic_vector(7038, 16),
53027 => conv_std_logic_vector(7245, 16),
53028 => conv_std_logic_vector(7452, 16),
53029 => conv_std_logic_vector(7659, 16),
53030 => conv_std_logic_vector(7866, 16),
53031 => conv_std_logic_vector(8073, 16),
53032 => conv_std_logic_vector(8280, 16),
53033 => conv_std_logic_vector(8487, 16),
53034 => conv_std_logic_vector(8694, 16),
53035 => conv_std_logic_vector(8901, 16),
53036 => conv_std_logic_vector(9108, 16),
53037 => conv_std_logic_vector(9315, 16),
53038 => conv_std_logic_vector(9522, 16),
53039 => conv_std_logic_vector(9729, 16),
53040 => conv_std_logic_vector(9936, 16),
53041 => conv_std_logic_vector(10143, 16),
53042 => conv_std_logic_vector(10350, 16),
53043 => conv_std_logic_vector(10557, 16),
53044 => conv_std_logic_vector(10764, 16),
53045 => conv_std_logic_vector(10971, 16),
53046 => conv_std_logic_vector(11178, 16),
53047 => conv_std_logic_vector(11385, 16),
53048 => conv_std_logic_vector(11592, 16),
53049 => conv_std_logic_vector(11799, 16),
53050 => conv_std_logic_vector(12006, 16),
53051 => conv_std_logic_vector(12213, 16),
53052 => conv_std_logic_vector(12420, 16),
53053 => conv_std_logic_vector(12627, 16),
53054 => conv_std_logic_vector(12834, 16),
53055 => conv_std_logic_vector(13041, 16),
53056 => conv_std_logic_vector(13248, 16),
53057 => conv_std_logic_vector(13455, 16),
53058 => conv_std_logic_vector(13662, 16),
53059 => conv_std_logic_vector(13869, 16),
53060 => conv_std_logic_vector(14076, 16),
53061 => conv_std_logic_vector(14283, 16),
53062 => conv_std_logic_vector(14490, 16),
53063 => conv_std_logic_vector(14697, 16),
53064 => conv_std_logic_vector(14904, 16),
53065 => conv_std_logic_vector(15111, 16),
53066 => conv_std_logic_vector(15318, 16),
53067 => conv_std_logic_vector(15525, 16),
53068 => conv_std_logic_vector(15732, 16),
53069 => conv_std_logic_vector(15939, 16),
53070 => conv_std_logic_vector(16146, 16),
53071 => conv_std_logic_vector(16353, 16),
53072 => conv_std_logic_vector(16560, 16),
53073 => conv_std_logic_vector(16767, 16),
53074 => conv_std_logic_vector(16974, 16),
53075 => conv_std_logic_vector(17181, 16),
53076 => conv_std_logic_vector(17388, 16),
53077 => conv_std_logic_vector(17595, 16),
53078 => conv_std_logic_vector(17802, 16),
53079 => conv_std_logic_vector(18009, 16),
53080 => conv_std_logic_vector(18216, 16),
53081 => conv_std_logic_vector(18423, 16),
53082 => conv_std_logic_vector(18630, 16),
53083 => conv_std_logic_vector(18837, 16),
53084 => conv_std_logic_vector(19044, 16),
53085 => conv_std_logic_vector(19251, 16),
53086 => conv_std_logic_vector(19458, 16),
53087 => conv_std_logic_vector(19665, 16),
53088 => conv_std_logic_vector(19872, 16),
53089 => conv_std_logic_vector(20079, 16),
53090 => conv_std_logic_vector(20286, 16),
53091 => conv_std_logic_vector(20493, 16),
53092 => conv_std_logic_vector(20700, 16),
53093 => conv_std_logic_vector(20907, 16),
53094 => conv_std_logic_vector(21114, 16),
53095 => conv_std_logic_vector(21321, 16),
53096 => conv_std_logic_vector(21528, 16),
53097 => conv_std_logic_vector(21735, 16),
53098 => conv_std_logic_vector(21942, 16),
53099 => conv_std_logic_vector(22149, 16),
53100 => conv_std_logic_vector(22356, 16),
53101 => conv_std_logic_vector(22563, 16),
53102 => conv_std_logic_vector(22770, 16),
53103 => conv_std_logic_vector(22977, 16),
53104 => conv_std_logic_vector(23184, 16),
53105 => conv_std_logic_vector(23391, 16),
53106 => conv_std_logic_vector(23598, 16),
53107 => conv_std_logic_vector(23805, 16),
53108 => conv_std_logic_vector(24012, 16),
53109 => conv_std_logic_vector(24219, 16),
53110 => conv_std_logic_vector(24426, 16),
53111 => conv_std_logic_vector(24633, 16),
53112 => conv_std_logic_vector(24840, 16),
53113 => conv_std_logic_vector(25047, 16),
53114 => conv_std_logic_vector(25254, 16),
53115 => conv_std_logic_vector(25461, 16),
53116 => conv_std_logic_vector(25668, 16),
53117 => conv_std_logic_vector(25875, 16),
53118 => conv_std_logic_vector(26082, 16),
53119 => conv_std_logic_vector(26289, 16),
53120 => conv_std_logic_vector(26496, 16),
53121 => conv_std_logic_vector(26703, 16),
53122 => conv_std_logic_vector(26910, 16),
53123 => conv_std_logic_vector(27117, 16),
53124 => conv_std_logic_vector(27324, 16),
53125 => conv_std_logic_vector(27531, 16),
53126 => conv_std_logic_vector(27738, 16),
53127 => conv_std_logic_vector(27945, 16),
53128 => conv_std_logic_vector(28152, 16),
53129 => conv_std_logic_vector(28359, 16),
53130 => conv_std_logic_vector(28566, 16),
53131 => conv_std_logic_vector(28773, 16),
53132 => conv_std_logic_vector(28980, 16),
53133 => conv_std_logic_vector(29187, 16),
53134 => conv_std_logic_vector(29394, 16),
53135 => conv_std_logic_vector(29601, 16),
53136 => conv_std_logic_vector(29808, 16),
53137 => conv_std_logic_vector(30015, 16),
53138 => conv_std_logic_vector(30222, 16),
53139 => conv_std_logic_vector(30429, 16),
53140 => conv_std_logic_vector(30636, 16),
53141 => conv_std_logic_vector(30843, 16),
53142 => conv_std_logic_vector(31050, 16),
53143 => conv_std_logic_vector(31257, 16),
53144 => conv_std_logic_vector(31464, 16),
53145 => conv_std_logic_vector(31671, 16),
53146 => conv_std_logic_vector(31878, 16),
53147 => conv_std_logic_vector(32085, 16),
53148 => conv_std_logic_vector(32292, 16),
53149 => conv_std_logic_vector(32499, 16),
53150 => conv_std_logic_vector(32706, 16),
53151 => conv_std_logic_vector(32913, 16),
53152 => conv_std_logic_vector(33120, 16),
53153 => conv_std_logic_vector(33327, 16),
53154 => conv_std_logic_vector(33534, 16),
53155 => conv_std_logic_vector(33741, 16),
53156 => conv_std_logic_vector(33948, 16),
53157 => conv_std_logic_vector(34155, 16),
53158 => conv_std_logic_vector(34362, 16),
53159 => conv_std_logic_vector(34569, 16),
53160 => conv_std_logic_vector(34776, 16),
53161 => conv_std_logic_vector(34983, 16),
53162 => conv_std_logic_vector(35190, 16),
53163 => conv_std_logic_vector(35397, 16),
53164 => conv_std_logic_vector(35604, 16),
53165 => conv_std_logic_vector(35811, 16),
53166 => conv_std_logic_vector(36018, 16),
53167 => conv_std_logic_vector(36225, 16),
53168 => conv_std_logic_vector(36432, 16),
53169 => conv_std_logic_vector(36639, 16),
53170 => conv_std_logic_vector(36846, 16),
53171 => conv_std_logic_vector(37053, 16),
53172 => conv_std_logic_vector(37260, 16),
53173 => conv_std_logic_vector(37467, 16),
53174 => conv_std_logic_vector(37674, 16),
53175 => conv_std_logic_vector(37881, 16),
53176 => conv_std_logic_vector(38088, 16),
53177 => conv_std_logic_vector(38295, 16),
53178 => conv_std_logic_vector(38502, 16),
53179 => conv_std_logic_vector(38709, 16),
53180 => conv_std_logic_vector(38916, 16),
53181 => conv_std_logic_vector(39123, 16),
53182 => conv_std_logic_vector(39330, 16),
53183 => conv_std_logic_vector(39537, 16),
53184 => conv_std_logic_vector(39744, 16),
53185 => conv_std_logic_vector(39951, 16),
53186 => conv_std_logic_vector(40158, 16),
53187 => conv_std_logic_vector(40365, 16),
53188 => conv_std_logic_vector(40572, 16),
53189 => conv_std_logic_vector(40779, 16),
53190 => conv_std_logic_vector(40986, 16),
53191 => conv_std_logic_vector(41193, 16),
53192 => conv_std_logic_vector(41400, 16),
53193 => conv_std_logic_vector(41607, 16),
53194 => conv_std_logic_vector(41814, 16),
53195 => conv_std_logic_vector(42021, 16),
53196 => conv_std_logic_vector(42228, 16),
53197 => conv_std_logic_vector(42435, 16),
53198 => conv_std_logic_vector(42642, 16),
53199 => conv_std_logic_vector(42849, 16),
53200 => conv_std_logic_vector(43056, 16),
53201 => conv_std_logic_vector(43263, 16),
53202 => conv_std_logic_vector(43470, 16),
53203 => conv_std_logic_vector(43677, 16),
53204 => conv_std_logic_vector(43884, 16),
53205 => conv_std_logic_vector(44091, 16),
53206 => conv_std_logic_vector(44298, 16),
53207 => conv_std_logic_vector(44505, 16),
53208 => conv_std_logic_vector(44712, 16),
53209 => conv_std_logic_vector(44919, 16),
53210 => conv_std_logic_vector(45126, 16),
53211 => conv_std_logic_vector(45333, 16),
53212 => conv_std_logic_vector(45540, 16),
53213 => conv_std_logic_vector(45747, 16),
53214 => conv_std_logic_vector(45954, 16),
53215 => conv_std_logic_vector(46161, 16),
53216 => conv_std_logic_vector(46368, 16),
53217 => conv_std_logic_vector(46575, 16),
53218 => conv_std_logic_vector(46782, 16),
53219 => conv_std_logic_vector(46989, 16),
53220 => conv_std_logic_vector(47196, 16),
53221 => conv_std_logic_vector(47403, 16),
53222 => conv_std_logic_vector(47610, 16),
53223 => conv_std_logic_vector(47817, 16),
53224 => conv_std_logic_vector(48024, 16),
53225 => conv_std_logic_vector(48231, 16),
53226 => conv_std_logic_vector(48438, 16),
53227 => conv_std_logic_vector(48645, 16),
53228 => conv_std_logic_vector(48852, 16),
53229 => conv_std_logic_vector(49059, 16),
53230 => conv_std_logic_vector(49266, 16),
53231 => conv_std_logic_vector(49473, 16),
53232 => conv_std_logic_vector(49680, 16),
53233 => conv_std_logic_vector(49887, 16),
53234 => conv_std_logic_vector(50094, 16),
53235 => conv_std_logic_vector(50301, 16),
53236 => conv_std_logic_vector(50508, 16),
53237 => conv_std_logic_vector(50715, 16),
53238 => conv_std_logic_vector(50922, 16),
53239 => conv_std_logic_vector(51129, 16),
53240 => conv_std_logic_vector(51336, 16),
53241 => conv_std_logic_vector(51543, 16),
53242 => conv_std_logic_vector(51750, 16),
53243 => conv_std_logic_vector(51957, 16),
53244 => conv_std_logic_vector(52164, 16),
53245 => conv_std_logic_vector(52371, 16),
53246 => conv_std_logic_vector(52578, 16),
53247 => conv_std_logic_vector(52785, 16),
53248 => conv_std_logic_vector(0, 16),
53249 => conv_std_logic_vector(208, 16),
53250 => conv_std_logic_vector(416, 16),
53251 => conv_std_logic_vector(624, 16),
53252 => conv_std_logic_vector(832, 16),
53253 => conv_std_logic_vector(1040, 16),
53254 => conv_std_logic_vector(1248, 16),
53255 => conv_std_logic_vector(1456, 16),
53256 => conv_std_logic_vector(1664, 16),
53257 => conv_std_logic_vector(1872, 16),
53258 => conv_std_logic_vector(2080, 16),
53259 => conv_std_logic_vector(2288, 16),
53260 => conv_std_logic_vector(2496, 16),
53261 => conv_std_logic_vector(2704, 16),
53262 => conv_std_logic_vector(2912, 16),
53263 => conv_std_logic_vector(3120, 16),
53264 => conv_std_logic_vector(3328, 16),
53265 => conv_std_logic_vector(3536, 16),
53266 => conv_std_logic_vector(3744, 16),
53267 => conv_std_logic_vector(3952, 16),
53268 => conv_std_logic_vector(4160, 16),
53269 => conv_std_logic_vector(4368, 16),
53270 => conv_std_logic_vector(4576, 16),
53271 => conv_std_logic_vector(4784, 16),
53272 => conv_std_logic_vector(4992, 16),
53273 => conv_std_logic_vector(5200, 16),
53274 => conv_std_logic_vector(5408, 16),
53275 => conv_std_logic_vector(5616, 16),
53276 => conv_std_logic_vector(5824, 16),
53277 => conv_std_logic_vector(6032, 16),
53278 => conv_std_logic_vector(6240, 16),
53279 => conv_std_logic_vector(6448, 16),
53280 => conv_std_logic_vector(6656, 16),
53281 => conv_std_logic_vector(6864, 16),
53282 => conv_std_logic_vector(7072, 16),
53283 => conv_std_logic_vector(7280, 16),
53284 => conv_std_logic_vector(7488, 16),
53285 => conv_std_logic_vector(7696, 16),
53286 => conv_std_logic_vector(7904, 16),
53287 => conv_std_logic_vector(8112, 16),
53288 => conv_std_logic_vector(8320, 16),
53289 => conv_std_logic_vector(8528, 16),
53290 => conv_std_logic_vector(8736, 16),
53291 => conv_std_logic_vector(8944, 16),
53292 => conv_std_logic_vector(9152, 16),
53293 => conv_std_logic_vector(9360, 16),
53294 => conv_std_logic_vector(9568, 16),
53295 => conv_std_logic_vector(9776, 16),
53296 => conv_std_logic_vector(9984, 16),
53297 => conv_std_logic_vector(10192, 16),
53298 => conv_std_logic_vector(10400, 16),
53299 => conv_std_logic_vector(10608, 16),
53300 => conv_std_logic_vector(10816, 16),
53301 => conv_std_logic_vector(11024, 16),
53302 => conv_std_logic_vector(11232, 16),
53303 => conv_std_logic_vector(11440, 16),
53304 => conv_std_logic_vector(11648, 16),
53305 => conv_std_logic_vector(11856, 16),
53306 => conv_std_logic_vector(12064, 16),
53307 => conv_std_logic_vector(12272, 16),
53308 => conv_std_logic_vector(12480, 16),
53309 => conv_std_logic_vector(12688, 16),
53310 => conv_std_logic_vector(12896, 16),
53311 => conv_std_logic_vector(13104, 16),
53312 => conv_std_logic_vector(13312, 16),
53313 => conv_std_logic_vector(13520, 16),
53314 => conv_std_logic_vector(13728, 16),
53315 => conv_std_logic_vector(13936, 16),
53316 => conv_std_logic_vector(14144, 16),
53317 => conv_std_logic_vector(14352, 16),
53318 => conv_std_logic_vector(14560, 16),
53319 => conv_std_logic_vector(14768, 16),
53320 => conv_std_logic_vector(14976, 16),
53321 => conv_std_logic_vector(15184, 16),
53322 => conv_std_logic_vector(15392, 16),
53323 => conv_std_logic_vector(15600, 16),
53324 => conv_std_logic_vector(15808, 16),
53325 => conv_std_logic_vector(16016, 16),
53326 => conv_std_logic_vector(16224, 16),
53327 => conv_std_logic_vector(16432, 16),
53328 => conv_std_logic_vector(16640, 16),
53329 => conv_std_logic_vector(16848, 16),
53330 => conv_std_logic_vector(17056, 16),
53331 => conv_std_logic_vector(17264, 16),
53332 => conv_std_logic_vector(17472, 16),
53333 => conv_std_logic_vector(17680, 16),
53334 => conv_std_logic_vector(17888, 16),
53335 => conv_std_logic_vector(18096, 16),
53336 => conv_std_logic_vector(18304, 16),
53337 => conv_std_logic_vector(18512, 16),
53338 => conv_std_logic_vector(18720, 16),
53339 => conv_std_logic_vector(18928, 16),
53340 => conv_std_logic_vector(19136, 16),
53341 => conv_std_logic_vector(19344, 16),
53342 => conv_std_logic_vector(19552, 16),
53343 => conv_std_logic_vector(19760, 16),
53344 => conv_std_logic_vector(19968, 16),
53345 => conv_std_logic_vector(20176, 16),
53346 => conv_std_logic_vector(20384, 16),
53347 => conv_std_logic_vector(20592, 16),
53348 => conv_std_logic_vector(20800, 16),
53349 => conv_std_logic_vector(21008, 16),
53350 => conv_std_logic_vector(21216, 16),
53351 => conv_std_logic_vector(21424, 16),
53352 => conv_std_logic_vector(21632, 16),
53353 => conv_std_logic_vector(21840, 16),
53354 => conv_std_logic_vector(22048, 16),
53355 => conv_std_logic_vector(22256, 16),
53356 => conv_std_logic_vector(22464, 16),
53357 => conv_std_logic_vector(22672, 16),
53358 => conv_std_logic_vector(22880, 16),
53359 => conv_std_logic_vector(23088, 16),
53360 => conv_std_logic_vector(23296, 16),
53361 => conv_std_logic_vector(23504, 16),
53362 => conv_std_logic_vector(23712, 16),
53363 => conv_std_logic_vector(23920, 16),
53364 => conv_std_logic_vector(24128, 16),
53365 => conv_std_logic_vector(24336, 16),
53366 => conv_std_logic_vector(24544, 16),
53367 => conv_std_logic_vector(24752, 16),
53368 => conv_std_logic_vector(24960, 16),
53369 => conv_std_logic_vector(25168, 16),
53370 => conv_std_logic_vector(25376, 16),
53371 => conv_std_logic_vector(25584, 16),
53372 => conv_std_logic_vector(25792, 16),
53373 => conv_std_logic_vector(26000, 16),
53374 => conv_std_logic_vector(26208, 16),
53375 => conv_std_logic_vector(26416, 16),
53376 => conv_std_logic_vector(26624, 16),
53377 => conv_std_logic_vector(26832, 16),
53378 => conv_std_logic_vector(27040, 16),
53379 => conv_std_logic_vector(27248, 16),
53380 => conv_std_logic_vector(27456, 16),
53381 => conv_std_logic_vector(27664, 16),
53382 => conv_std_logic_vector(27872, 16),
53383 => conv_std_logic_vector(28080, 16),
53384 => conv_std_logic_vector(28288, 16),
53385 => conv_std_logic_vector(28496, 16),
53386 => conv_std_logic_vector(28704, 16),
53387 => conv_std_logic_vector(28912, 16),
53388 => conv_std_logic_vector(29120, 16),
53389 => conv_std_logic_vector(29328, 16),
53390 => conv_std_logic_vector(29536, 16),
53391 => conv_std_logic_vector(29744, 16),
53392 => conv_std_logic_vector(29952, 16),
53393 => conv_std_logic_vector(30160, 16),
53394 => conv_std_logic_vector(30368, 16),
53395 => conv_std_logic_vector(30576, 16),
53396 => conv_std_logic_vector(30784, 16),
53397 => conv_std_logic_vector(30992, 16),
53398 => conv_std_logic_vector(31200, 16),
53399 => conv_std_logic_vector(31408, 16),
53400 => conv_std_logic_vector(31616, 16),
53401 => conv_std_logic_vector(31824, 16),
53402 => conv_std_logic_vector(32032, 16),
53403 => conv_std_logic_vector(32240, 16),
53404 => conv_std_logic_vector(32448, 16),
53405 => conv_std_logic_vector(32656, 16),
53406 => conv_std_logic_vector(32864, 16),
53407 => conv_std_logic_vector(33072, 16),
53408 => conv_std_logic_vector(33280, 16),
53409 => conv_std_logic_vector(33488, 16),
53410 => conv_std_logic_vector(33696, 16),
53411 => conv_std_logic_vector(33904, 16),
53412 => conv_std_logic_vector(34112, 16),
53413 => conv_std_logic_vector(34320, 16),
53414 => conv_std_logic_vector(34528, 16),
53415 => conv_std_logic_vector(34736, 16),
53416 => conv_std_logic_vector(34944, 16),
53417 => conv_std_logic_vector(35152, 16),
53418 => conv_std_logic_vector(35360, 16),
53419 => conv_std_logic_vector(35568, 16),
53420 => conv_std_logic_vector(35776, 16),
53421 => conv_std_logic_vector(35984, 16),
53422 => conv_std_logic_vector(36192, 16),
53423 => conv_std_logic_vector(36400, 16),
53424 => conv_std_logic_vector(36608, 16),
53425 => conv_std_logic_vector(36816, 16),
53426 => conv_std_logic_vector(37024, 16),
53427 => conv_std_logic_vector(37232, 16),
53428 => conv_std_logic_vector(37440, 16),
53429 => conv_std_logic_vector(37648, 16),
53430 => conv_std_logic_vector(37856, 16),
53431 => conv_std_logic_vector(38064, 16),
53432 => conv_std_logic_vector(38272, 16),
53433 => conv_std_logic_vector(38480, 16),
53434 => conv_std_logic_vector(38688, 16),
53435 => conv_std_logic_vector(38896, 16),
53436 => conv_std_logic_vector(39104, 16),
53437 => conv_std_logic_vector(39312, 16),
53438 => conv_std_logic_vector(39520, 16),
53439 => conv_std_logic_vector(39728, 16),
53440 => conv_std_logic_vector(39936, 16),
53441 => conv_std_logic_vector(40144, 16),
53442 => conv_std_logic_vector(40352, 16),
53443 => conv_std_logic_vector(40560, 16),
53444 => conv_std_logic_vector(40768, 16),
53445 => conv_std_logic_vector(40976, 16),
53446 => conv_std_logic_vector(41184, 16),
53447 => conv_std_logic_vector(41392, 16),
53448 => conv_std_logic_vector(41600, 16),
53449 => conv_std_logic_vector(41808, 16),
53450 => conv_std_logic_vector(42016, 16),
53451 => conv_std_logic_vector(42224, 16),
53452 => conv_std_logic_vector(42432, 16),
53453 => conv_std_logic_vector(42640, 16),
53454 => conv_std_logic_vector(42848, 16),
53455 => conv_std_logic_vector(43056, 16),
53456 => conv_std_logic_vector(43264, 16),
53457 => conv_std_logic_vector(43472, 16),
53458 => conv_std_logic_vector(43680, 16),
53459 => conv_std_logic_vector(43888, 16),
53460 => conv_std_logic_vector(44096, 16),
53461 => conv_std_logic_vector(44304, 16),
53462 => conv_std_logic_vector(44512, 16),
53463 => conv_std_logic_vector(44720, 16),
53464 => conv_std_logic_vector(44928, 16),
53465 => conv_std_logic_vector(45136, 16),
53466 => conv_std_logic_vector(45344, 16),
53467 => conv_std_logic_vector(45552, 16),
53468 => conv_std_logic_vector(45760, 16),
53469 => conv_std_logic_vector(45968, 16),
53470 => conv_std_logic_vector(46176, 16),
53471 => conv_std_logic_vector(46384, 16),
53472 => conv_std_logic_vector(46592, 16),
53473 => conv_std_logic_vector(46800, 16),
53474 => conv_std_logic_vector(47008, 16),
53475 => conv_std_logic_vector(47216, 16),
53476 => conv_std_logic_vector(47424, 16),
53477 => conv_std_logic_vector(47632, 16),
53478 => conv_std_logic_vector(47840, 16),
53479 => conv_std_logic_vector(48048, 16),
53480 => conv_std_logic_vector(48256, 16),
53481 => conv_std_logic_vector(48464, 16),
53482 => conv_std_logic_vector(48672, 16),
53483 => conv_std_logic_vector(48880, 16),
53484 => conv_std_logic_vector(49088, 16),
53485 => conv_std_logic_vector(49296, 16),
53486 => conv_std_logic_vector(49504, 16),
53487 => conv_std_logic_vector(49712, 16),
53488 => conv_std_logic_vector(49920, 16),
53489 => conv_std_logic_vector(50128, 16),
53490 => conv_std_logic_vector(50336, 16),
53491 => conv_std_logic_vector(50544, 16),
53492 => conv_std_logic_vector(50752, 16),
53493 => conv_std_logic_vector(50960, 16),
53494 => conv_std_logic_vector(51168, 16),
53495 => conv_std_logic_vector(51376, 16),
53496 => conv_std_logic_vector(51584, 16),
53497 => conv_std_logic_vector(51792, 16),
53498 => conv_std_logic_vector(52000, 16),
53499 => conv_std_logic_vector(52208, 16),
53500 => conv_std_logic_vector(52416, 16),
53501 => conv_std_logic_vector(52624, 16),
53502 => conv_std_logic_vector(52832, 16),
53503 => conv_std_logic_vector(53040, 16),
53504 => conv_std_logic_vector(0, 16),
53505 => conv_std_logic_vector(209, 16),
53506 => conv_std_logic_vector(418, 16),
53507 => conv_std_logic_vector(627, 16),
53508 => conv_std_logic_vector(836, 16),
53509 => conv_std_logic_vector(1045, 16),
53510 => conv_std_logic_vector(1254, 16),
53511 => conv_std_logic_vector(1463, 16),
53512 => conv_std_logic_vector(1672, 16),
53513 => conv_std_logic_vector(1881, 16),
53514 => conv_std_logic_vector(2090, 16),
53515 => conv_std_logic_vector(2299, 16),
53516 => conv_std_logic_vector(2508, 16),
53517 => conv_std_logic_vector(2717, 16),
53518 => conv_std_logic_vector(2926, 16),
53519 => conv_std_logic_vector(3135, 16),
53520 => conv_std_logic_vector(3344, 16),
53521 => conv_std_logic_vector(3553, 16),
53522 => conv_std_logic_vector(3762, 16),
53523 => conv_std_logic_vector(3971, 16),
53524 => conv_std_logic_vector(4180, 16),
53525 => conv_std_logic_vector(4389, 16),
53526 => conv_std_logic_vector(4598, 16),
53527 => conv_std_logic_vector(4807, 16),
53528 => conv_std_logic_vector(5016, 16),
53529 => conv_std_logic_vector(5225, 16),
53530 => conv_std_logic_vector(5434, 16),
53531 => conv_std_logic_vector(5643, 16),
53532 => conv_std_logic_vector(5852, 16),
53533 => conv_std_logic_vector(6061, 16),
53534 => conv_std_logic_vector(6270, 16),
53535 => conv_std_logic_vector(6479, 16),
53536 => conv_std_logic_vector(6688, 16),
53537 => conv_std_logic_vector(6897, 16),
53538 => conv_std_logic_vector(7106, 16),
53539 => conv_std_logic_vector(7315, 16),
53540 => conv_std_logic_vector(7524, 16),
53541 => conv_std_logic_vector(7733, 16),
53542 => conv_std_logic_vector(7942, 16),
53543 => conv_std_logic_vector(8151, 16),
53544 => conv_std_logic_vector(8360, 16),
53545 => conv_std_logic_vector(8569, 16),
53546 => conv_std_logic_vector(8778, 16),
53547 => conv_std_logic_vector(8987, 16),
53548 => conv_std_logic_vector(9196, 16),
53549 => conv_std_logic_vector(9405, 16),
53550 => conv_std_logic_vector(9614, 16),
53551 => conv_std_logic_vector(9823, 16),
53552 => conv_std_logic_vector(10032, 16),
53553 => conv_std_logic_vector(10241, 16),
53554 => conv_std_logic_vector(10450, 16),
53555 => conv_std_logic_vector(10659, 16),
53556 => conv_std_logic_vector(10868, 16),
53557 => conv_std_logic_vector(11077, 16),
53558 => conv_std_logic_vector(11286, 16),
53559 => conv_std_logic_vector(11495, 16),
53560 => conv_std_logic_vector(11704, 16),
53561 => conv_std_logic_vector(11913, 16),
53562 => conv_std_logic_vector(12122, 16),
53563 => conv_std_logic_vector(12331, 16),
53564 => conv_std_logic_vector(12540, 16),
53565 => conv_std_logic_vector(12749, 16),
53566 => conv_std_logic_vector(12958, 16),
53567 => conv_std_logic_vector(13167, 16),
53568 => conv_std_logic_vector(13376, 16),
53569 => conv_std_logic_vector(13585, 16),
53570 => conv_std_logic_vector(13794, 16),
53571 => conv_std_logic_vector(14003, 16),
53572 => conv_std_logic_vector(14212, 16),
53573 => conv_std_logic_vector(14421, 16),
53574 => conv_std_logic_vector(14630, 16),
53575 => conv_std_logic_vector(14839, 16),
53576 => conv_std_logic_vector(15048, 16),
53577 => conv_std_logic_vector(15257, 16),
53578 => conv_std_logic_vector(15466, 16),
53579 => conv_std_logic_vector(15675, 16),
53580 => conv_std_logic_vector(15884, 16),
53581 => conv_std_logic_vector(16093, 16),
53582 => conv_std_logic_vector(16302, 16),
53583 => conv_std_logic_vector(16511, 16),
53584 => conv_std_logic_vector(16720, 16),
53585 => conv_std_logic_vector(16929, 16),
53586 => conv_std_logic_vector(17138, 16),
53587 => conv_std_logic_vector(17347, 16),
53588 => conv_std_logic_vector(17556, 16),
53589 => conv_std_logic_vector(17765, 16),
53590 => conv_std_logic_vector(17974, 16),
53591 => conv_std_logic_vector(18183, 16),
53592 => conv_std_logic_vector(18392, 16),
53593 => conv_std_logic_vector(18601, 16),
53594 => conv_std_logic_vector(18810, 16),
53595 => conv_std_logic_vector(19019, 16),
53596 => conv_std_logic_vector(19228, 16),
53597 => conv_std_logic_vector(19437, 16),
53598 => conv_std_logic_vector(19646, 16),
53599 => conv_std_logic_vector(19855, 16),
53600 => conv_std_logic_vector(20064, 16),
53601 => conv_std_logic_vector(20273, 16),
53602 => conv_std_logic_vector(20482, 16),
53603 => conv_std_logic_vector(20691, 16),
53604 => conv_std_logic_vector(20900, 16),
53605 => conv_std_logic_vector(21109, 16),
53606 => conv_std_logic_vector(21318, 16),
53607 => conv_std_logic_vector(21527, 16),
53608 => conv_std_logic_vector(21736, 16),
53609 => conv_std_logic_vector(21945, 16),
53610 => conv_std_logic_vector(22154, 16),
53611 => conv_std_logic_vector(22363, 16),
53612 => conv_std_logic_vector(22572, 16),
53613 => conv_std_logic_vector(22781, 16),
53614 => conv_std_logic_vector(22990, 16),
53615 => conv_std_logic_vector(23199, 16),
53616 => conv_std_logic_vector(23408, 16),
53617 => conv_std_logic_vector(23617, 16),
53618 => conv_std_logic_vector(23826, 16),
53619 => conv_std_logic_vector(24035, 16),
53620 => conv_std_logic_vector(24244, 16),
53621 => conv_std_logic_vector(24453, 16),
53622 => conv_std_logic_vector(24662, 16),
53623 => conv_std_logic_vector(24871, 16),
53624 => conv_std_logic_vector(25080, 16),
53625 => conv_std_logic_vector(25289, 16),
53626 => conv_std_logic_vector(25498, 16),
53627 => conv_std_logic_vector(25707, 16),
53628 => conv_std_logic_vector(25916, 16),
53629 => conv_std_logic_vector(26125, 16),
53630 => conv_std_logic_vector(26334, 16),
53631 => conv_std_logic_vector(26543, 16),
53632 => conv_std_logic_vector(26752, 16),
53633 => conv_std_logic_vector(26961, 16),
53634 => conv_std_logic_vector(27170, 16),
53635 => conv_std_logic_vector(27379, 16),
53636 => conv_std_logic_vector(27588, 16),
53637 => conv_std_logic_vector(27797, 16),
53638 => conv_std_logic_vector(28006, 16),
53639 => conv_std_logic_vector(28215, 16),
53640 => conv_std_logic_vector(28424, 16),
53641 => conv_std_logic_vector(28633, 16),
53642 => conv_std_logic_vector(28842, 16),
53643 => conv_std_logic_vector(29051, 16),
53644 => conv_std_logic_vector(29260, 16),
53645 => conv_std_logic_vector(29469, 16),
53646 => conv_std_logic_vector(29678, 16),
53647 => conv_std_logic_vector(29887, 16),
53648 => conv_std_logic_vector(30096, 16),
53649 => conv_std_logic_vector(30305, 16),
53650 => conv_std_logic_vector(30514, 16),
53651 => conv_std_logic_vector(30723, 16),
53652 => conv_std_logic_vector(30932, 16),
53653 => conv_std_logic_vector(31141, 16),
53654 => conv_std_logic_vector(31350, 16),
53655 => conv_std_logic_vector(31559, 16),
53656 => conv_std_logic_vector(31768, 16),
53657 => conv_std_logic_vector(31977, 16),
53658 => conv_std_logic_vector(32186, 16),
53659 => conv_std_logic_vector(32395, 16),
53660 => conv_std_logic_vector(32604, 16),
53661 => conv_std_logic_vector(32813, 16),
53662 => conv_std_logic_vector(33022, 16),
53663 => conv_std_logic_vector(33231, 16),
53664 => conv_std_logic_vector(33440, 16),
53665 => conv_std_logic_vector(33649, 16),
53666 => conv_std_logic_vector(33858, 16),
53667 => conv_std_logic_vector(34067, 16),
53668 => conv_std_logic_vector(34276, 16),
53669 => conv_std_logic_vector(34485, 16),
53670 => conv_std_logic_vector(34694, 16),
53671 => conv_std_logic_vector(34903, 16),
53672 => conv_std_logic_vector(35112, 16),
53673 => conv_std_logic_vector(35321, 16),
53674 => conv_std_logic_vector(35530, 16),
53675 => conv_std_logic_vector(35739, 16),
53676 => conv_std_logic_vector(35948, 16),
53677 => conv_std_logic_vector(36157, 16),
53678 => conv_std_logic_vector(36366, 16),
53679 => conv_std_logic_vector(36575, 16),
53680 => conv_std_logic_vector(36784, 16),
53681 => conv_std_logic_vector(36993, 16),
53682 => conv_std_logic_vector(37202, 16),
53683 => conv_std_logic_vector(37411, 16),
53684 => conv_std_logic_vector(37620, 16),
53685 => conv_std_logic_vector(37829, 16),
53686 => conv_std_logic_vector(38038, 16),
53687 => conv_std_logic_vector(38247, 16),
53688 => conv_std_logic_vector(38456, 16),
53689 => conv_std_logic_vector(38665, 16),
53690 => conv_std_logic_vector(38874, 16),
53691 => conv_std_logic_vector(39083, 16),
53692 => conv_std_logic_vector(39292, 16),
53693 => conv_std_logic_vector(39501, 16),
53694 => conv_std_logic_vector(39710, 16),
53695 => conv_std_logic_vector(39919, 16),
53696 => conv_std_logic_vector(40128, 16),
53697 => conv_std_logic_vector(40337, 16),
53698 => conv_std_logic_vector(40546, 16),
53699 => conv_std_logic_vector(40755, 16),
53700 => conv_std_logic_vector(40964, 16),
53701 => conv_std_logic_vector(41173, 16),
53702 => conv_std_logic_vector(41382, 16),
53703 => conv_std_logic_vector(41591, 16),
53704 => conv_std_logic_vector(41800, 16),
53705 => conv_std_logic_vector(42009, 16),
53706 => conv_std_logic_vector(42218, 16),
53707 => conv_std_logic_vector(42427, 16),
53708 => conv_std_logic_vector(42636, 16),
53709 => conv_std_logic_vector(42845, 16),
53710 => conv_std_logic_vector(43054, 16),
53711 => conv_std_logic_vector(43263, 16),
53712 => conv_std_logic_vector(43472, 16),
53713 => conv_std_logic_vector(43681, 16),
53714 => conv_std_logic_vector(43890, 16),
53715 => conv_std_logic_vector(44099, 16),
53716 => conv_std_logic_vector(44308, 16),
53717 => conv_std_logic_vector(44517, 16),
53718 => conv_std_logic_vector(44726, 16),
53719 => conv_std_logic_vector(44935, 16),
53720 => conv_std_logic_vector(45144, 16),
53721 => conv_std_logic_vector(45353, 16),
53722 => conv_std_logic_vector(45562, 16),
53723 => conv_std_logic_vector(45771, 16),
53724 => conv_std_logic_vector(45980, 16),
53725 => conv_std_logic_vector(46189, 16),
53726 => conv_std_logic_vector(46398, 16),
53727 => conv_std_logic_vector(46607, 16),
53728 => conv_std_logic_vector(46816, 16),
53729 => conv_std_logic_vector(47025, 16),
53730 => conv_std_logic_vector(47234, 16),
53731 => conv_std_logic_vector(47443, 16),
53732 => conv_std_logic_vector(47652, 16),
53733 => conv_std_logic_vector(47861, 16),
53734 => conv_std_logic_vector(48070, 16),
53735 => conv_std_logic_vector(48279, 16),
53736 => conv_std_logic_vector(48488, 16),
53737 => conv_std_logic_vector(48697, 16),
53738 => conv_std_logic_vector(48906, 16),
53739 => conv_std_logic_vector(49115, 16),
53740 => conv_std_logic_vector(49324, 16),
53741 => conv_std_logic_vector(49533, 16),
53742 => conv_std_logic_vector(49742, 16),
53743 => conv_std_logic_vector(49951, 16),
53744 => conv_std_logic_vector(50160, 16),
53745 => conv_std_logic_vector(50369, 16),
53746 => conv_std_logic_vector(50578, 16),
53747 => conv_std_logic_vector(50787, 16),
53748 => conv_std_logic_vector(50996, 16),
53749 => conv_std_logic_vector(51205, 16),
53750 => conv_std_logic_vector(51414, 16),
53751 => conv_std_logic_vector(51623, 16),
53752 => conv_std_logic_vector(51832, 16),
53753 => conv_std_logic_vector(52041, 16),
53754 => conv_std_logic_vector(52250, 16),
53755 => conv_std_logic_vector(52459, 16),
53756 => conv_std_logic_vector(52668, 16),
53757 => conv_std_logic_vector(52877, 16),
53758 => conv_std_logic_vector(53086, 16),
53759 => conv_std_logic_vector(53295, 16),
53760 => conv_std_logic_vector(0, 16),
53761 => conv_std_logic_vector(210, 16),
53762 => conv_std_logic_vector(420, 16),
53763 => conv_std_logic_vector(630, 16),
53764 => conv_std_logic_vector(840, 16),
53765 => conv_std_logic_vector(1050, 16),
53766 => conv_std_logic_vector(1260, 16),
53767 => conv_std_logic_vector(1470, 16),
53768 => conv_std_logic_vector(1680, 16),
53769 => conv_std_logic_vector(1890, 16),
53770 => conv_std_logic_vector(2100, 16),
53771 => conv_std_logic_vector(2310, 16),
53772 => conv_std_logic_vector(2520, 16),
53773 => conv_std_logic_vector(2730, 16),
53774 => conv_std_logic_vector(2940, 16),
53775 => conv_std_logic_vector(3150, 16),
53776 => conv_std_logic_vector(3360, 16),
53777 => conv_std_logic_vector(3570, 16),
53778 => conv_std_logic_vector(3780, 16),
53779 => conv_std_logic_vector(3990, 16),
53780 => conv_std_logic_vector(4200, 16),
53781 => conv_std_logic_vector(4410, 16),
53782 => conv_std_logic_vector(4620, 16),
53783 => conv_std_logic_vector(4830, 16),
53784 => conv_std_logic_vector(5040, 16),
53785 => conv_std_logic_vector(5250, 16),
53786 => conv_std_logic_vector(5460, 16),
53787 => conv_std_logic_vector(5670, 16),
53788 => conv_std_logic_vector(5880, 16),
53789 => conv_std_logic_vector(6090, 16),
53790 => conv_std_logic_vector(6300, 16),
53791 => conv_std_logic_vector(6510, 16),
53792 => conv_std_logic_vector(6720, 16),
53793 => conv_std_logic_vector(6930, 16),
53794 => conv_std_logic_vector(7140, 16),
53795 => conv_std_logic_vector(7350, 16),
53796 => conv_std_logic_vector(7560, 16),
53797 => conv_std_logic_vector(7770, 16),
53798 => conv_std_logic_vector(7980, 16),
53799 => conv_std_logic_vector(8190, 16),
53800 => conv_std_logic_vector(8400, 16),
53801 => conv_std_logic_vector(8610, 16),
53802 => conv_std_logic_vector(8820, 16),
53803 => conv_std_logic_vector(9030, 16),
53804 => conv_std_logic_vector(9240, 16),
53805 => conv_std_logic_vector(9450, 16),
53806 => conv_std_logic_vector(9660, 16),
53807 => conv_std_logic_vector(9870, 16),
53808 => conv_std_logic_vector(10080, 16),
53809 => conv_std_logic_vector(10290, 16),
53810 => conv_std_logic_vector(10500, 16),
53811 => conv_std_logic_vector(10710, 16),
53812 => conv_std_logic_vector(10920, 16),
53813 => conv_std_logic_vector(11130, 16),
53814 => conv_std_logic_vector(11340, 16),
53815 => conv_std_logic_vector(11550, 16),
53816 => conv_std_logic_vector(11760, 16),
53817 => conv_std_logic_vector(11970, 16),
53818 => conv_std_logic_vector(12180, 16),
53819 => conv_std_logic_vector(12390, 16),
53820 => conv_std_logic_vector(12600, 16),
53821 => conv_std_logic_vector(12810, 16),
53822 => conv_std_logic_vector(13020, 16),
53823 => conv_std_logic_vector(13230, 16),
53824 => conv_std_logic_vector(13440, 16),
53825 => conv_std_logic_vector(13650, 16),
53826 => conv_std_logic_vector(13860, 16),
53827 => conv_std_logic_vector(14070, 16),
53828 => conv_std_logic_vector(14280, 16),
53829 => conv_std_logic_vector(14490, 16),
53830 => conv_std_logic_vector(14700, 16),
53831 => conv_std_logic_vector(14910, 16),
53832 => conv_std_logic_vector(15120, 16),
53833 => conv_std_logic_vector(15330, 16),
53834 => conv_std_logic_vector(15540, 16),
53835 => conv_std_logic_vector(15750, 16),
53836 => conv_std_logic_vector(15960, 16),
53837 => conv_std_logic_vector(16170, 16),
53838 => conv_std_logic_vector(16380, 16),
53839 => conv_std_logic_vector(16590, 16),
53840 => conv_std_logic_vector(16800, 16),
53841 => conv_std_logic_vector(17010, 16),
53842 => conv_std_logic_vector(17220, 16),
53843 => conv_std_logic_vector(17430, 16),
53844 => conv_std_logic_vector(17640, 16),
53845 => conv_std_logic_vector(17850, 16),
53846 => conv_std_logic_vector(18060, 16),
53847 => conv_std_logic_vector(18270, 16),
53848 => conv_std_logic_vector(18480, 16),
53849 => conv_std_logic_vector(18690, 16),
53850 => conv_std_logic_vector(18900, 16),
53851 => conv_std_logic_vector(19110, 16),
53852 => conv_std_logic_vector(19320, 16),
53853 => conv_std_logic_vector(19530, 16),
53854 => conv_std_logic_vector(19740, 16),
53855 => conv_std_logic_vector(19950, 16),
53856 => conv_std_logic_vector(20160, 16),
53857 => conv_std_logic_vector(20370, 16),
53858 => conv_std_logic_vector(20580, 16),
53859 => conv_std_logic_vector(20790, 16),
53860 => conv_std_logic_vector(21000, 16),
53861 => conv_std_logic_vector(21210, 16),
53862 => conv_std_logic_vector(21420, 16),
53863 => conv_std_logic_vector(21630, 16),
53864 => conv_std_logic_vector(21840, 16),
53865 => conv_std_logic_vector(22050, 16),
53866 => conv_std_logic_vector(22260, 16),
53867 => conv_std_logic_vector(22470, 16),
53868 => conv_std_logic_vector(22680, 16),
53869 => conv_std_logic_vector(22890, 16),
53870 => conv_std_logic_vector(23100, 16),
53871 => conv_std_logic_vector(23310, 16),
53872 => conv_std_logic_vector(23520, 16),
53873 => conv_std_logic_vector(23730, 16),
53874 => conv_std_logic_vector(23940, 16),
53875 => conv_std_logic_vector(24150, 16),
53876 => conv_std_logic_vector(24360, 16),
53877 => conv_std_logic_vector(24570, 16),
53878 => conv_std_logic_vector(24780, 16),
53879 => conv_std_logic_vector(24990, 16),
53880 => conv_std_logic_vector(25200, 16),
53881 => conv_std_logic_vector(25410, 16),
53882 => conv_std_logic_vector(25620, 16),
53883 => conv_std_logic_vector(25830, 16),
53884 => conv_std_logic_vector(26040, 16),
53885 => conv_std_logic_vector(26250, 16),
53886 => conv_std_logic_vector(26460, 16),
53887 => conv_std_logic_vector(26670, 16),
53888 => conv_std_logic_vector(26880, 16),
53889 => conv_std_logic_vector(27090, 16),
53890 => conv_std_logic_vector(27300, 16),
53891 => conv_std_logic_vector(27510, 16),
53892 => conv_std_logic_vector(27720, 16),
53893 => conv_std_logic_vector(27930, 16),
53894 => conv_std_logic_vector(28140, 16),
53895 => conv_std_logic_vector(28350, 16),
53896 => conv_std_logic_vector(28560, 16),
53897 => conv_std_logic_vector(28770, 16),
53898 => conv_std_logic_vector(28980, 16),
53899 => conv_std_logic_vector(29190, 16),
53900 => conv_std_logic_vector(29400, 16),
53901 => conv_std_logic_vector(29610, 16),
53902 => conv_std_logic_vector(29820, 16),
53903 => conv_std_logic_vector(30030, 16),
53904 => conv_std_logic_vector(30240, 16),
53905 => conv_std_logic_vector(30450, 16),
53906 => conv_std_logic_vector(30660, 16),
53907 => conv_std_logic_vector(30870, 16),
53908 => conv_std_logic_vector(31080, 16),
53909 => conv_std_logic_vector(31290, 16),
53910 => conv_std_logic_vector(31500, 16),
53911 => conv_std_logic_vector(31710, 16),
53912 => conv_std_logic_vector(31920, 16),
53913 => conv_std_logic_vector(32130, 16),
53914 => conv_std_logic_vector(32340, 16),
53915 => conv_std_logic_vector(32550, 16),
53916 => conv_std_logic_vector(32760, 16),
53917 => conv_std_logic_vector(32970, 16),
53918 => conv_std_logic_vector(33180, 16),
53919 => conv_std_logic_vector(33390, 16),
53920 => conv_std_logic_vector(33600, 16),
53921 => conv_std_logic_vector(33810, 16),
53922 => conv_std_logic_vector(34020, 16),
53923 => conv_std_logic_vector(34230, 16),
53924 => conv_std_logic_vector(34440, 16),
53925 => conv_std_logic_vector(34650, 16),
53926 => conv_std_logic_vector(34860, 16),
53927 => conv_std_logic_vector(35070, 16),
53928 => conv_std_logic_vector(35280, 16),
53929 => conv_std_logic_vector(35490, 16),
53930 => conv_std_logic_vector(35700, 16),
53931 => conv_std_logic_vector(35910, 16),
53932 => conv_std_logic_vector(36120, 16),
53933 => conv_std_logic_vector(36330, 16),
53934 => conv_std_logic_vector(36540, 16),
53935 => conv_std_logic_vector(36750, 16),
53936 => conv_std_logic_vector(36960, 16),
53937 => conv_std_logic_vector(37170, 16),
53938 => conv_std_logic_vector(37380, 16),
53939 => conv_std_logic_vector(37590, 16),
53940 => conv_std_logic_vector(37800, 16),
53941 => conv_std_logic_vector(38010, 16),
53942 => conv_std_logic_vector(38220, 16),
53943 => conv_std_logic_vector(38430, 16),
53944 => conv_std_logic_vector(38640, 16),
53945 => conv_std_logic_vector(38850, 16),
53946 => conv_std_logic_vector(39060, 16),
53947 => conv_std_logic_vector(39270, 16),
53948 => conv_std_logic_vector(39480, 16),
53949 => conv_std_logic_vector(39690, 16),
53950 => conv_std_logic_vector(39900, 16),
53951 => conv_std_logic_vector(40110, 16),
53952 => conv_std_logic_vector(40320, 16),
53953 => conv_std_logic_vector(40530, 16),
53954 => conv_std_logic_vector(40740, 16),
53955 => conv_std_logic_vector(40950, 16),
53956 => conv_std_logic_vector(41160, 16),
53957 => conv_std_logic_vector(41370, 16),
53958 => conv_std_logic_vector(41580, 16),
53959 => conv_std_logic_vector(41790, 16),
53960 => conv_std_logic_vector(42000, 16),
53961 => conv_std_logic_vector(42210, 16),
53962 => conv_std_logic_vector(42420, 16),
53963 => conv_std_logic_vector(42630, 16),
53964 => conv_std_logic_vector(42840, 16),
53965 => conv_std_logic_vector(43050, 16),
53966 => conv_std_logic_vector(43260, 16),
53967 => conv_std_logic_vector(43470, 16),
53968 => conv_std_logic_vector(43680, 16),
53969 => conv_std_logic_vector(43890, 16),
53970 => conv_std_logic_vector(44100, 16),
53971 => conv_std_logic_vector(44310, 16),
53972 => conv_std_logic_vector(44520, 16),
53973 => conv_std_logic_vector(44730, 16),
53974 => conv_std_logic_vector(44940, 16),
53975 => conv_std_logic_vector(45150, 16),
53976 => conv_std_logic_vector(45360, 16),
53977 => conv_std_logic_vector(45570, 16),
53978 => conv_std_logic_vector(45780, 16),
53979 => conv_std_logic_vector(45990, 16),
53980 => conv_std_logic_vector(46200, 16),
53981 => conv_std_logic_vector(46410, 16),
53982 => conv_std_logic_vector(46620, 16),
53983 => conv_std_logic_vector(46830, 16),
53984 => conv_std_logic_vector(47040, 16),
53985 => conv_std_logic_vector(47250, 16),
53986 => conv_std_logic_vector(47460, 16),
53987 => conv_std_logic_vector(47670, 16),
53988 => conv_std_logic_vector(47880, 16),
53989 => conv_std_logic_vector(48090, 16),
53990 => conv_std_logic_vector(48300, 16),
53991 => conv_std_logic_vector(48510, 16),
53992 => conv_std_logic_vector(48720, 16),
53993 => conv_std_logic_vector(48930, 16),
53994 => conv_std_logic_vector(49140, 16),
53995 => conv_std_logic_vector(49350, 16),
53996 => conv_std_logic_vector(49560, 16),
53997 => conv_std_logic_vector(49770, 16),
53998 => conv_std_logic_vector(49980, 16),
53999 => conv_std_logic_vector(50190, 16),
54000 => conv_std_logic_vector(50400, 16),
54001 => conv_std_logic_vector(50610, 16),
54002 => conv_std_logic_vector(50820, 16),
54003 => conv_std_logic_vector(51030, 16),
54004 => conv_std_logic_vector(51240, 16),
54005 => conv_std_logic_vector(51450, 16),
54006 => conv_std_logic_vector(51660, 16),
54007 => conv_std_logic_vector(51870, 16),
54008 => conv_std_logic_vector(52080, 16),
54009 => conv_std_logic_vector(52290, 16),
54010 => conv_std_logic_vector(52500, 16),
54011 => conv_std_logic_vector(52710, 16),
54012 => conv_std_logic_vector(52920, 16),
54013 => conv_std_logic_vector(53130, 16),
54014 => conv_std_logic_vector(53340, 16),
54015 => conv_std_logic_vector(53550, 16),
54016 => conv_std_logic_vector(0, 16),
54017 => conv_std_logic_vector(211, 16),
54018 => conv_std_logic_vector(422, 16),
54019 => conv_std_logic_vector(633, 16),
54020 => conv_std_logic_vector(844, 16),
54021 => conv_std_logic_vector(1055, 16),
54022 => conv_std_logic_vector(1266, 16),
54023 => conv_std_logic_vector(1477, 16),
54024 => conv_std_logic_vector(1688, 16),
54025 => conv_std_logic_vector(1899, 16),
54026 => conv_std_logic_vector(2110, 16),
54027 => conv_std_logic_vector(2321, 16),
54028 => conv_std_logic_vector(2532, 16),
54029 => conv_std_logic_vector(2743, 16),
54030 => conv_std_logic_vector(2954, 16),
54031 => conv_std_logic_vector(3165, 16),
54032 => conv_std_logic_vector(3376, 16),
54033 => conv_std_logic_vector(3587, 16),
54034 => conv_std_logic_vector(3798, 16),
54035 => conv_std_logic_vector(4009, 16),
54036 => conv_std_logic_vector(4220, 16),
54037 => conv_std_logic_vector(4431, 16),
54038 => conv_std_logic_vector(4642, 16),
54039 => conv_std_logic_vector(4853, 16),
54040 => conv_std_logic_vector(5064, 16),
54041 => conv_std_logic_vector(5275, 16),
54042 => conv_std_logic_vector(5486, 16),
54043 => conv_std_logic_vector(5697, 16),
54044 => conv_std_logic_vector(5908, 16),
54045 => conv_std_logic_vector(6119, 16),
54046 => conv_std_logic_vector(6330, 16),
54047 => conv_std_logic_vector(6541, 16),
54048 => conv_std_logic_vector(6752, 16),
54049 => conv_std_logic_vector(6963, 16),
54050 => conv_std_logic_vector(7174, 16),
54051 => conv_std_logic_vector(7385, 16),
54052 => conv_std_logic_vector(7596, 16),
54053 => conv_std_logic_vector(7807, 16),
54054 => conv_std_logic_vector(8018, 16),
54055 => conv_std_logic_vector(8229, 16),
54056 => conv_std_logic_vector(8440, 16),
54057 => conv_std_logic_vector(8651, 16),
54058 => conv_std_logic_vector(8862, 16),
54059 => conv_std_logic_vector(9073, 16),
54060 => conv_std_logic_vector(9284, 16),
54061 => conv_std_logic_vector(9495, 16),
54062 => conv_std_logic_vector(9706, 16),
54063 => conv_std_logic_vector(9917, 16),
54064 => conv_std_logic_vector(10128, 16),
54065 => conv_std_logic_vector(10339, 16),
54066 => conv_std_logic_vector(10550, 16),
54067 => conv_std_logic_vector(10761, 16),
54068 => conv_std_logic_vector(10972, 16),
54069 => conv_std_logic_vector(11183, 16),
54070 => conv_std_logic_vector(11394, 16),
54071 => conv_std_logic_vector(11605, 16),
54072 => conv_std_logic_vector(11816, 16),
54073 => conv_std_logic_vector(12027, 16),
54074 => conv_std_logic_vector(12238, 16),
54075 => conv_std_logic_vector(12449, 16),
54076 => conv_std_logic_vector(12660, 16),
54077 => conv_std_logic_vector(12871, 16),
54078 => conv_std_logic_vector(13082, 16),
54079 => conv_std_logic_vector(13293, 16),
54080 => conv_std_logic_vector(13504, 16),
54081 => conv_std_logic_vector(13715, 16),
54082 => conv_std_logic_vector(13926, 16),
54083 => conv_std_logic_vector(14137, 16),
54084 => conv_std_logic_vector(14348, 16),
54085 => conv_std_logic_vector(14559, 16),
54086 => conv_std_logic_vector(14770, 16),
54087 => conv_std_logic_vector(14981, 16),
54088 => conv_std_logic_vector(15192, 16),
54089 => conv_std_logic_vector(15403, 16),
54090 => conv_std_logic_vector(15614, 16),
54091 => conv_std_logic_vector(15825, 16),
54092 => conv_std_logic_vector(16036, 16),
54093 => conv_std_logic_vector(16247, 16),
54094 => conv_std_logic_vector(16458, 16),
54095 => conv_std_logic_vector(16669, 16),
54096 => conv_std_logic_vector(16880, 16),
54097 => conv_std_logic_vector(17091, 16),
54098 => conv_std_logic_vector(17302, 16),
54099 => conv_std_logic_vector(17513, 16),
54100 => conv_std_logic_vector(17724, 16),
54101 => conv_std_logic_vector(17935, 16),
54102 => conv_std_logic_vector(18146, 16),
54103 => conv_std_logic_vector(18357, 16),
54104 => conv_std_logic_vector(18568, 16),
54105 => conv_std_logic_vector(18779, 16),
54106 => conv_std_logic_vector(18990, 16),
54107 => conv_std_logic_vector(19201, 16),
54108 => conv_std_logic_vector(19412, 16),
54109 => conv_std_logic_vector(19623, 16),
54110 => conv_std_logic_vector(19834, 16),
54111 => conv_std_logic_vector(20045, 16),
54112 => conv_std_logic_vector(20256, 16),
54113 => conv_std_logic_vector(20467, 16),
54114 => conv_std_logic_vector(20678, 16),
54115 => conv_std_logic_vector(20889, 16),
54116 => conv_std_logic_vector(21100, 16),
54117 => conv_std_logic_vector(21311, 16),
54118 => conv_std_logic_vector(21522, 16),
54119 => conv_std_logic_vector(21733, 16),
54120 => conv_std_logic_vector(21944, 16),
54121 => conv_std_logic_vector(22155, 16),
54122 => conv_std_logic_vector(22366, 16),
54123 => conv_std_logic_vector(22577, 16),
54124 => conv_std_logic_vector(22788, 16),
54125 => conv_std_logic_vector(22999, 16),
54126 => conv_std_logic_vector(23210, 16),
54127 => conv_std_logic_vector(23421, 16),
54128 => conv_std_logic_vector(23632, 16),
54129 => conv_std_logic_vector(23843, 16),
54130 => conv_std_logic_vector(24054, 16),
54131 => conv_std_logic_vector(24265, 16),
54132 => conv_std_logic_vector(24476, 16),
54133 => conv_std_logic_vector(24687, 16),
54134 => conv_std_logic_vector(24898, 16),
54135 => conv_std_logic_vector(25109, 16),
54136 => conv_std_logic_vector(25320, 16),
54137 => conv_std_logic_vector(25531, 16),
54138 => conv_std_logic_vector(25742, 16),
54139 => conv_std_logic_vector(25953, 16),
54140 => conv_std_logic_vector(26164, 16),
54141 => conv_std_logic_vector(26375, 16),
54142 => conv_std_logic_vector(26586, 16),
54143 => conv_std_logic_vector(26797, 16),
54144 => conv_std_logic_vector(27008, 16),
54145 => conv_std_logic_vector(27219, 16),
54146 => conv_std_logic_vector(27430, 16),
54147 => conv_std_logic_vector(27641, 16),
54148 => conv_std_logic_vector(27852, 16),
54149 => conv_std_logic_vector(28063, 16),
54150 => conv_std_logic_vector(28274, 16),
54151 => conv_std_logic_vector(28485, 16),
54152 => conv_std_logic_vector(28696, 16),
54153 => conv_std_logic_vector(28907, 16),
54154 => conv_std_logic_vector(29118, 16),
54155 => conv_std_logic_vector(29329, 16),
54156 => conv_std_logic_vector(29540, 16),
54157 => conv_std_logic_vector(29751, 16),
54158 => conv_std_logic_vector(29962, 16),
54159 => conv_std_logic_vector(30173, 16),
54160 => conv_std_logic_vector(30384, 16),
54161 => conv_std_logic_vector(30595, 16),
54162 => conv_std_logic_vector(30806, 16),
54163 => conv_std_logic_vector(31017, 16),
54164 => conv_std_logic_vector(31228, 16),
54165 => conv_std_logic_vector(31439, 16),
54166 => conv_std_logic_vector(31650, 16),
54167 => conv_std_logic_vector(31861, 16),
54168 => conv_std_logic_vector(32072, 16),
54169 => conv_std_logic_vector(32283, 16),
54170 => conv_std_logic_vector(32494, 16),
54171 => conv_std_logic_vector(32705, 16),
54172 => conv_std_logic_vector(32916, 16),
54173 => conv_std_logic_vector(33127, 16),
54174 => conv_std_logic_vector(33338, 16),
54175 => conv_std_logic_vector(33549, 16),
54176 => conv_std_logic_vector(33760, 16),
54177 => conv_std_logic_vector(33971, 16),
54178 => conv_std_logic_vector(34182, 16),
54179 => conv_std_logic_vector(34393, 16),
54180 => conv_std_logic_vector(34604, 16),
54181 => conv_std_logic_vector(34815, 16),
54182 => conv_std_logic_vector(35026, 16),
54183 => conv_std_logic_vector(35237, 16),
54184 => conv_std_logic_vector(35448, 16),
54185 => conv_std_logic_vector(35659, 16),
54186 => conv_std_logic_vector(35870, 16),
54187 => conv_std_logic_vector(36081, 16),
54188 => conv_std_logic_vector(36292, 16),
54189 => conv_std_logic_vector(36503, 16),
54190 => conv_std_logic_vector(36714, 16),
54191 => conv_std_logic_vector(36925, 16),
54192 => conv_std_logic_vector(37136, 16),
54193 => conv_std_logic_vector(37347, 16),
54194 => conv_std_logic_vector(37558, 16),
54195 => conv_std_logic_vector(37769, 16),
54196 => conv_std_logic_vector(37980, 16),
54197 => conv_std_logic_vector(38191, 16),
54198 => conv_std_logic_vector(38402, 16),
54199 => conv_std_logic_vector(38613, 16),
54200 => conv_std_logic_vector(38824, 16),
54201 => conv_std_logic_vector(39035, 16),
54202 => conv_std_logic_vector(39246, 16),
54203 => conv_std_logic_vector(39457, 16),
54204 => conv_std_logic_vector(39668, 16),
54205 => conv_std_logic_vector(39879, 16),
54206 => conv_std_logic_vector(40090, 16),
54207 => conv_std_logic_vector(40301, 16),
54208 => conv_std_logic_vector(40512, 16),
54209 => conv_std_logic_vector(40723, 16),
54210 => conv_std_logic_vector(40934, 16),
54211 => conv_std_logic_vector(41145, 16),
54212 => conv_std_logic_vector(41356, 16),
54213 => conv_std_logic_vector(41567, 16),
54214 => conv_std_logic_vector(41778, 16),
54215 => conv_std_logic_vector(41989, 16),
54216 => conv_std_logic_vector(42200, 16),
54217 => conv_std_logic_vector(42411, 16),
54218 => conv_std_logic_vector(42622, 16),
54219 => conv_std_logic_vector(42833, 16),
54220 => conv_std_logic_vector(43044, 16),
54221 => conv_std_logic_vector(43255, 16),
54222 => conv_std_logic_vector(43466, 16),
54223 => conv_std_logic_vector(43677, 16),
54224 => conv_std_logic_vector(43888, 16),
54225 => conv_std_logic_vector(44099, 16),
54226 => conv_std_logic_vector(44310, 16),
54227 => conv_std_logic_vector(44521, 16),
54228 => conv_std_logic_vector(44732, 16),
54229 => conv_std_logic_vector(44943, 16),
54230 => conv_std_logic_vector(45154, 16),
54231 => conv_std_logic_vector(45365, 16),
54232 => conv_std_logic_vector(45576, 16),
54233 => conv_std_logic_vector(45787, 16),
54234 => conv_std_logic_vector(45998, 16),
54235 => conv_std_logic_vector(46209, 16),
54236 => conv_std_logic_vector(46420, 16),
54237 => conv_std_logic_vector(46631, 16),
54238 => conv_std_logic_vector(46842, 16),
54239 => conv_std_logic_vector(47053, 16),
54240 => conv_std_logic_vector(47264, 16),
54241 => conv_std_logic_vector(47475, 16),
54242 => conv_std_logic_vector(47686, 16),
54243 => conv_std_logic_vector(47897, 16),
54244 => conv_std_logic_vector(48108, 16),
54245 => conv_std_logic_vector(48319, 16),
54246 => conv_std_logic_vector(48530, 16),
54247 => conv_std_logic_vector(48741, 16),
54248 => conv_std_logic_vector(48952, 16),
54249 => conv_std_logic_vector(49163, 16),
54250 => conv_std_logic_vector(49374, 16),
54251 => conv_std_logic_vector(49585, 16),
54252 => conv_std_logic_vector(49796, 16),
54253 => conv_std_logic_vector(50007, 16),
54254 => conv_std_logic_vector(50218, 16),
54255 => conv_std_logic_vector(50429, 16),
54256 => conv_std_logic_vector(50640, 16),
54257 => conv_std_logic_vector(50851, 16),
54258 => conv_std_logic_vector(51062, 16),
54259 => conv_std_logic_vector(51273, 16),
54260 => conv_std_logic_vector(51484, 16),
54261 => conv_std_logic_vector(51695, 16),
54262 => conv_std_logic_vector(51906, 16),
54263 => conv_std_logic_vector(52117, 16),
54264 => conv_std_logic_vector(52328, 16),
54265 => conv_std_logic_vector(52539, 16),
54266 => conv_std_logic_vector(52750, 16),
54267 => conv_std_logic_vector(52961, 16),
54268 => conv_std_logic_vector(53172, 16),
54269 => conv_std_logic_vector(53383, 16),
54270 => conv_std_logic_vector(53594, 16),
54271 => conv_std_logic_vector(53805, 16),
54272 => conv_std_logic_vector(0, 16),
54273 => conv_std_logic_vector(212, 16),
54274 => conv_std_logic_vector(424, 16),
54275 => conv_std_logic_vector(636, 16),
54276 => conv_std_logic_vector(848, 16),
54277 => conv_std_logic_vector(1060, 16),
54278 => conv_std_logic_vector(1272, 16),
54279 => conv_std_logic_vector(1484, 16),
54280 => conv_std_logic_vector(1696, 16),
54281 => conv_std_logic_vector(1908, 16),
54282 => conv_std_logic_vector(2120, 16),
54283 => conv_std_logic_vector(2332, 16),
54284 => conv_std_logic_vector(2544, 16),
54285 => conv_std_logic_vector(2756, 16),
54286 => conv_std_logic_vector(2968, 16),
54287 => conv_std_logic_vector(3180, 16),
54288 => conv_std_logic_vector(3392, 16),
54289 => conv_std_logic_vector(3604, 16),
54290 => conv_std_logic_vector(3816, 16),
54291 => conv_std_logic_vector(4028, 16),
54292 => conv_std_logic_vector(4240, 16),
54293 => conv_std_logic_vector(4452, 16),
54294 => conv_std_logic_vector(4664, 16),
54295 => conv_std_logic_vector(4876, 16),
54296 => conv_std_logic_vector(5088, 16),
54297 => conv_std_logic_vector(5300, 16),
54298 => conv_std_logic_vector(5512, 16),
54299 => conv_std_logic_vector(5724, 16),
54300 => conv_std_logic_vector(5936, 16),
54301 => conv_std_logic_vector(6148, 16),
54302 => conv_std_logic_vector(6360, 16),
54303 => conv_std_logic_vector(6572, 16),
54304 => conv_std_logic_vector(6784, 16),
54305 => conv_std_logic_vector(6996, 16),
54306 => conv_std_logic_vector(7208, 16),
54307 => conv_std_logic_vector(7420, 16),
54308 => conv_std_logic_vector(7632, 16),
54309 => conv_std_logic_vector(7844, 16),
54310 => conv_std_logic_vector(8056, 16),
54311 => conv_std_logic_vector(8268, 16),
54312 => conv_std_logic_vector(8480, 16),
54313 => conv_std_logic_vector(8692, 16),
54314 => conv_std_logic_vector(8904, 16),
54315 => conv_std_logic_vector(9116, 16),
54316 => conv_std_logic_vector(9328, 16),
54317 => conv_std_logic_vector(9540, 16),
54318 => conv_std_logic_vector(9752, 16),
54319 => conv_std_logic_vector(9964, 16),
54320 => conv_std_logic_vector(10176, 16),
54321 => conv_std_logic_vector(10388, 16),
54322 => conv_std_logic_vector(10600, 16),
54323 => conv_std_logic_vector(10812, 16),
54324 => conv_std_logic_vector(11024, 16),
54325 => conv_std_logic_vector(11236, 16),
54326 => conv_std_logic_vector(11448, 16),
54327 => conv_std_logic_vector(11660, 16),
54328 => conv_std_logic_vector(11872, 16),
54329 => conv_std_logic_vector(12084, 16),
54330 => conv_std_logic_vector(12296, 16),
54331 => conv_std_logic_vector(12508, 16),
54332 => conv_std_logic_vector(12720, 16),
54333 => conv_std_logic_vector(12932, 16),
54334 => conv_std_logic_vector(13144, 16),
54335 => conv_std_logic_vector(13356, 16),
54336 => conv_std_logic_vector(13568, 16),
54337 => conv_std_logic_vector(13780, 16),
54338 => conv_std_logic_vector(13992, 16),
54339 => conv_std_logic_vector(14204, 16),
54340 => conv_std_logic_vector(14416, 16),
54341 => conv_std_logic_vector(14628, 16),
54342 => conv_std_logic_vector(14840, 16),
54343 => conv_std_logic_vector(15052, 16),
54344 => conv_std_logic_vector(15264, 16),
54345 => conv_std_logic_vector(15476, 16),
54346 => conv_std_logic_vector(15688, 16),
54347 => conv_std_logic_vector(15900, 16),
54348 => conv_std_logic_vector(16112, 16),
54349 => conv_std_logic_vector(16324, 16),
54350 => conv_std_logic_vector(16536, 16),
54351 => conv_std_logic_vector(16748, 16),
54352 => conv_std_logic_vector(16960, 16),
54353 => conv_std_logic_vector(17172, 16),
54354 => conv_std_logic_vector(17384, 16),
54355 => conv_std_logic_vector(17596, 16),
54356 => conv_std_logic_vector(17808, 16),
54357 => conv_std_logic_vector(18020, 16),
54358 => conv_std_logic_vector(18232, 16),
54359 => conv_std_logic_vector(18444, 16),
54360 => conv_std_logic_vector(18656, 16),
54361 => conv_std_logic_vector(18868, 16),
54362 => conv_std_logic_vector(19080, 16),
54363 => conv_std_logic_vector(19292, 16),
54364 => conv_std_logic_vector(19504, 16),
54365 => conv_std_logic_vector(19716, 16),
54366 => conv_std_logic_vector(19928, 16),
54367 => conv_std_logic_vector(20140, 16),
54368 => conv_std_logic_vector(20352, 16),
54369 => conv_std_logic_vector(20564, 16),
54370 => conv_std_logic_vector(20776, 16),
54371 => conv_std_logic_vector(20988, 16),
54372 => conv_std_logic_vector(21200, 16),
54373 => conv_std_logic_vector(21412, 16),
54374 => conv_std_logic_vector(21624, 16),
54375 => conv_std_logic_vector(21836, 16),
54376 => conv_std_logic_vector(22048, 16),
54377 => conv_std_logic_vector(22260, 16),
54378 => conv_std_logic_vector(22472, 16),
54379 => conv_std_logic_vector(22684, 16),
54380 => conv_std_logic_vector(22896, 16),
54381 => conv_std_logic_vector(23108, 16),
54382 => conv_std_logic_vector(23320, 16),
54383 => conv_std_logic_vector(23532, 16),
54384 => conv_std_logic_vector(23744, 16),
54385 => conv_std_logic_vector(23956, 16),
54386 => conv_std_logic_vector(24168, 16),
54387 => conv_std_logic_vector(24380, 16),
54388 => conv_std_logic_vector(24592, 16),
54389 => conv_std_logic_vector(24804, 16),
54390 => conv_std_logic_vector(25016, 16),
54391 => conv_std_logic_vector(25228, 16),
54392 => conv_std_logic_vector(25440, 16),
54393 => conv_std_logic_vector(25652, 16),
54394 => conv_std_logic_vector(25864, 16),
54395 => conv_std_logic_vector(26076, 16),
54396 => conv_std_logic_vector(26288, 16),
54397 => conv_std_logic_vector(26500, 16),
54398 => conv_std_logic_vector(26712, 16),
54399 => conv_std_logic_vector(26924, 16),
54400 => conv_std_logic_vector(27136, 16),
54401 => conv_std_logic_vector(27348, 16),
54402 => conv_std_logic_vector(27560, 16),
54403 => conv_std_logic_vector(27772, 16),
54404 => conv_std_logic_vector(27984, 16),
54405 => conv_std_logic_vector(28196, 16),
54406 => conv_std_logic_vector(28408, 16),
54407 => conv_std_logic_vector(28620, 16),
54408 => conv_std_logic_vector(28832, 16),
54409 => conv_std_logic_vector(29044, 16),
54410 => conv_std_logic_vector(29256, 16),
54411 => conv_std_logic_vector(29468, 16),
54412 => conv_std_logic_vector(29680, 16),
54413 => conv_std_logic_vector(29892, 16),
54414 => conv_std_logic_vector(30104, 16),
54415 => conv_std_logic_vector(30316, 16),
54416 => conv_std_logic_vector(30528, 16),
54417 => conv_std_logic_vector(30740, 16),
54418 => conv_std_logic_vector(30952, 16),
54419 => conv_std_logic_vector(31164, 16),
54420 => conv_std_logic_vector(31376, 16),
54421 => conv_std_logic_vector(31588, 16),
54422 => conv_std_logic_vector(31800, 16),
54423 => conv_std_logic_vector(32012, 16),
54424 => conv_std_logic_vector(32224, 16),
54425 => conv_std_logic_vector(32436, 16),
54426 => conv_std_logic_vector(32648, 16),
54427 => conv_std_logic_vector(32860, 16),
54428 => conv_std_logic_vector(33072, 16),
54429 => conv_std_logic_vector(33284, 16),
54430 => conv_std_logic_vector(33496, 16),
54431 => conv_std_logic_vector(33708, 16),
54432 => conv_std_logic_vector(33920, 16),
54433 => conv_std_logic_vector(34132, 16),
54434 => conv_std_logic_vector(34344, 16),
54435 => conv_std_logic_vector(34556, 16),
54436 => conv_std_logic_vector(34768, 16),
54437 => conv_std_logic_vector(34980, 16),
54438 => conv_std_logic_vector(35192, 16),
54439 => conv_std_logic_vector(35404, 16),
54440 => conv_std_logic_vector(35616, 16),
54441 => conv_std_logic_vector(35828, 16),
54442 => conv_std_logic_vector(36040, 16),
54443 => conv_std_logic_vector(36252, 16),
54444 => conv_std_logic_vector(36464, 16),
54445 => conv_std_logic_vector(36676, 16),
54446 => conv_std_logic_vector(36888, 16),
54447 => conv_std_logic_vector(37100, 16),
54448 => conv_std_logic_vector(37312, 16),
54449 => conv_std_logic_vector(37524, 16),
54450 => conv_std_logic_vector(37736, 16),
54451 => conv_std_logic_vector(37948, 16),
54452 => conv_std_logic_vector(38160, 16),
54453 => conv_std_logic_vector(38372, 16),
54454 => conv_std_logic_vector(38584, 16),
54455 => conv_std_logic_vector(38796, 16),
54456 => conv_std_logic_vector(39008, 16),
54457 => conv_std_logic_vector(39220, 16),
54458 => conv_std_logic_vector(39432, 16),
54459 => conv_std_logic_vector(39644, 16),
54460 => conv_std_logic_vector(39856, 16),
54461 => conv_std_logic_vector(40068, 16),
54462 => conv_std_logic_vector(40280, 16),
54463 => conv_std_logic_vector(40492, 16),
54464 => conv_std_logic_vector(40704, 16),
54465 => conv_std_logic_vector(40916, 16),
54466 => conv_std_logic_vector(41128, 16),
54467 => conv_std_logic_vector(41340, 16),
54468 => conv_std_logic_vector(41552, 16),
54469 => conv_std_logic_vector(41764, 16),
54470 => conv_std_logic_vector(41976, 16),
54471 => conv_std_logic_vector(42188, 16),
54472 => conv_std_logic_vector(42400, 16),
54473 => conv_std_logic_vector(42612, 16),
54474 => conv_std_logic_vector(42824, 16),
54475 => conv_std_logic_vector(43036, 16),
54476 => conv_std_logic_vector(43248, 16),
54477 => conv_std_logic_vector(43460, 16),
54478 => conv_std_logic_vector(43672, 16),
54479 => conv_std_logic_vector(43884, 16),
54480 => conv_std_logic_vector(44096, 16),
54481 => conv_std_logic_vector(44308, 16),
54482 => conv_std_logic_vector(44520, 16),
54483 => conv_std_logic_vector(44732, 16),
54484 => conv_std_logic_vector(44944, 16),
54485 => conv_std_logic_vector(45156, 16),
54486 => conv_std_logic_vector(45368, 16),
54487 => conv_std_logic_vector(45580, 16),
54488 => conv_std_logic_vector(45792, 16),
54489 => conv_std_logic_vector(46004, 16),
54490 => conv_std_logic_vector(46216, 16),
54491 => conv_std_logic_vector(46428, 16),
54492 => conv_std_logic_vector(46640, 16),
54493 => conv_std_logic_vector(46852, 16),
54494 => conv_std_logic_vector(47064, 16),
54495 => conv_std_logic_vector(47276, 16),
54496 => conv_std_logic_vector(47488, 16),
54497 => conv_std_logic_vector(47700, 16),
54498 => conv_std_logic_vector(47912, 16),
54499 => conv_std_logic_vector(48124, 16),
54500 => conv_std_logic_vector(48336, 16),
54501 => conv_std_logic_vector(48548, 16),
54502 => conv_std_logic_vector(48760, 16),
54503 => conv_std_logic_vector(48972, 16),
54504 => conv_std_logic_vector(49184, 16),
54505 => conv_std_logic_vector(49396, 16),
54506 => conv_std_logic_vector(49608, 16),
54507 => conv_std_logic_vector(49820, 16),
54508 => conv_std_logic_vector(50032, 16),
54509 => conv_std_logic_vector(50244, 16),
54510 => conv_std_logic_vector(50456, 16),
54511 => conv_std_logic_vector(50668, 16),
54512 => conv_std_logic_vector(50880, 16),
54513 => conv_std_logic_vector(51092, 16),
54514 => conv_std_logic_vector(51304, 16),
54515 => conv_std_logic_vector(51516, 16),
54516 => conv_std_logic_vector(51728, 16),
54517 => conv_std_logic_vector(51940, 16),
54518 => conv_std_logic_vector(52152, 16),
54519 => conv_std_logic_vector(52364, 16),
54520 => conv_std_logic_vector(52576, 16),
54521 => conv_std_logic_vector(52788, 16),
54522 => conv_std_logic_vector(53000, 16),
54523 => conv_std_logic_vector(53212, 16),
54524 => conv_std_logic_vector(53424, 16),
54525 => conv_std_logic_vector(53636, 16),
54526 => conv_std_logic_vector(53848, 16),
54527 => conv_std_logic_vector(54060, 16),
54528 => conv_std_logic_vector(0, 16),
54529 => conv_std_logic_vector(213, 16),
54530 => conv_std_logic_vector(426, 16),
54531 => conv_std_logic_vector(639, 16),
54532 => conv_std_logic_vector(852, 16),
54533 => conv_std_logic_vector(1065, 16),
54534 => conv_std_logic_vector(1278, 16),
54535 => conv_std_logic_vector(1491, 16),
54536 => conv_std_logic_vector(1704, 16),
54537 => conv_std_logic_vector(1917, 16),
54538 => conv_std_logic_vector(2130, 16),
54539 => conv_std_logic_vector(2343, 16),
54540 => conv_std_logic_vector(2556, 16),
54541 => conv_std_logic_vector(2769, 16),
54542 => conv_std_logic_vector(2982, 16),
54543 => conv_std_logic_vector(3195, 16),
54544 => conv_std_logic_vector(3408, 16),
54545 => conv_std_logic_vector(3621, 16),
54546 => conv_std_logic_vector(3834, 16),
54547 => conv_std_logic_vector(4047, 16),
54548 => conv_std_logic_vector(4260, 16),
54549 => conv_std_logic_vector(4473, 16),
54550 => conv_std_logic_vector(4686, 16),
54551 => conv_std_logic_vector(4899, 16),
54552 => conv_std_logic_vector(5112, 16),
54553 => conv_std_logic_vector(5325, 16),
54554 => conv_std_logic_vector(5538, 16),
54555 => conv_std_logic_vector(5751, 16),
54556 => conv_std_logic_vector(5964, 16),
54557 => conv_std_logic_vector(6177, 16),
54558 => conv_std_logic_vector(6390, 16),
54559 => conv_std_logic_vector(6603, 16),
54560 => conv_std_logic_vector(6816, 16),
54561 => conv_std_logic_vector(7029, 16),
54562 => conv_std_logic_vector(7242, 16),
54563 => conv_std_logic_vector(7455, 16),
54564 => conv_std_logic_vector(7668, 16),
54565 => conv_std_logic_vector(7881, 16),
54566 => conv_std_logic_vector(8094, 16),
54567 => conv_std_logic_vector(8307, 16),
54568 => conv_std_logic_vector(8520, 16),
54569 => conv_std_logic_vector(8733, 16),
54570 => conv_std_logic_vector(8946, 16),
54571 => conv_std_logic_vector(9159, 16),
54572 => conv_std_logic_vector(9372, 16),
54573 => conv_std_logic_vector(9585, 16),
54574 => conv_std_logic_vector(9798, 16),
54575 => conv_std_logic_vector(10011, 16),
54576 => conv_std_logic_vector(10224, 16),
54577 => conv_std_logic_vector(10437, 16),
54578 => conv_std_logic_vector(10650, 16),
54579 => conv_std_logic_vector(10863, 16),
54580 => conv_std_logic_vector(11076, 16),
54581 => conv_std_logic_vector(11289, 16),
54582 => conv_std_logic_vector(11502, 16),
54583 => conv_std_logic_vector(11715, 16),
54584 => conv_std_logic_vector(11928, 16),
54585 => conv_std_logic_vector(12141, 16),
54586 => conv_std_logic_vector(12354, 16),
54587 => conv_std_logic_vector(12567, 16),
54588 => conv_std_logic_vector(12780, 16),
54589 => conv_std_logic_vector(12993, 16),
54590 => conv_std_logic_vector(13206, 16),
54591 => conv_std_logic_vector(13419, 16),
54592 => conv_std_logic_vector(13632, 16),
54593 => conv_std_logic_vector(13845, 16),
54594 => conv_std_logic_vector(14058, 16),
54595 => conv_std_logic_vector(14271, 16),
54596 => conv_std_logic_vector(14484, 16),
54597 => conv_std_logic_vector(14697, 16),
54598 => conv_std_logic_vector(14910, 16),
54599 => conv_std_logic_vector(15123, 16),
54600 => conv_std_logic_vector(15336, 16),
54601 => conv_std_logic_vector(15549, 16),
54602 => conv_std_logic_vector(15762, 16),
54603 => conv_std_logic_vector(15975, 16),
54604 => conv_std_logic_vector(16188, 16),
54605 => conv_std_logic_vector(16401, 16),
54606 => conv_std_logic_vector(16614, 16),
54607 => conv_std_logic_vector(16827, 16),
54608 => conv_std_logic_vector(17040, 16),
54609 => conv_std_logic_vector(17253, 16),
54610 => conv_std_logic_vector(17466, 16),
54611 => conv_std_logic_vector(17679, 16),
54612 => conv_std_logic_vector(17892, 16),
54613 => conv_std_logic_vector(18105, 16),
54614 => conv_std_logic_vector(18318, 16),
54615 => conv_std_logic_vector(18531, 16),
54616 => conv_std_logic_vector(18744, 16),
54617 => conv_std_logic_vector(18957, 16),
54618 => conv_std_logic_vector(19170, 16),
54619 => conv_std_logic_vector(19383, 16),
54620 => conv_std_logic_vector(19596, 16),
54621 => conv_std_logic_vector(19809, 16),
54622 => conv_std_logic_vector(20022, 16),
54623 => conv_std_logic_vector(20235, 16),
54624 => conv_std_logic_vector(20448, 16),
54625 => conv_std_logic_vector(20661, 16),
54626 => conv_std_logic_vector(20874, 16),
54627 => conv_std_logic_vector(21087, 16),
54628 => conv_std_logic_vector(21300, 16),
54629 => conv_std_logic_vector(21513, 16),
54630 => conv_std_logic_vector(21726, 16),
54631 => conv_std_logic_vector(21939, 16),
54632 => conv_std_logic_vector(22152, 16),
54633 => conv_std_logic_vector(22365, 16),
54634 => conv_std_logic_vector(22578, 16),
54635 => conv_std_logic_vector(22791, 16),
54636 => conv_std_logic_vector(23004, 16),
54637 => conv_std_logic_vector(23217, 16),
54638 => conv_std_logic_vector(23430, 16),
54639 => conv_std_logic_vector(23643, 16),
54640 => conv_std_logic_vector(23856, 16),
54641 => conv_std_logic_vector(24069, 16),
54642 => conv_std_logic_vector(24282, 16),
54643 => conv_std_logic_vector(24495, 16),
54644 => conv_std_logic_vector(24708, 16),
54645 => conv_std_logic_vector(24921, 16),
54646 => conv_std_logic_vector(25134, 16),
54647 => conv_std_logic_vector(25347, 16),
54648 => conv_std_logic_vector(25560, 16),
54649 => conv_std_logic_vector(25773, 16),
54650 => conv_std_logic_vector(25986, 16),
54651 => conv_std_logic_vector(26199, 16),
54652 => conv_std_logic_vector(26412, 16),
54653 => conv_std_logic_vector(26625, 16),
54654 => conv_std_logic_vector(26838, 16),
54655 => conv_std_logic_vector(27051, 16),
54656 => conv_std_logic_vector(27264, 16),
54657 => conv_std_logic_vector(27477, 16),
54658 => conv_std_logic_vector(27690, 16),
54659 => conv_std_logic_vector(27903, 16),
54660 => conv_std_logic_vector(28116, 16),
54661 => conv_std_logic_vector(28329, 16),
54662 => conv_std_logic_vector(28542, 16),
54663 => conv_std_logic_vector(28755, 16),
54664 => conv_std_logic_vector(28968, 16),
54665 => conv_std_logic_vector(29181, 16),
54666 => conv_std_logic_vector(29394, 16),
54667 => conv_std_logic_vector(29607, 16),
54668 => conv_std_logic_vector(29820, 16),
54669 => conv_std_logic_vector(30033, 16),
54670 => conv_std_logic_vector(30246, 16),
54671 => conv_std_logic_vector(30459, 16),
54672 => conv_std_logic_vector(30672, 16),
54673 => conv_std_logic_vector(30885, 16),
54674 => conv_std_logic_vector(31098, 16),
54675 => conv_std_logic_vector(31311, 16),
54676 => conv_std_logic_vector(31524, 16),
54677 => conv_std_logic_vector(31737, 16),
54678 => conv_std_logic_vector(31950, 16),
54679 => conv_std_logic_vector(32163, 16),
54680 => conv_std_logic_vector(32376, 16),
54681 => conv_std_logic_vector(32589, 16),
54682 => conv_std_logic_vector(32802, 16),
54683 => conv_std_logic_vector(33015, 16),
54684 => conv_std_logic_vector(33228, 16),
54685 => conv_std_logic_vector(33441, 16),
54686 => conv_std_logic_vector(33654, 16),
54687 => conv_std_logic_vector(33867, 16),
54688 => conv_std_logic_vector(34080, 16),
54689 => conv_std_logic_vector(34293, 16),
54690 => conv_std_logic_vector(34506, 16),
54691 => conv_std_logic_vector(34719, 16),
54692 => conv_std_logic_vector(34932, 16),
54693 => conv_std_logic_vector(35145, 16),
54694 => conv_std_logic_vector(35358, 16),
54695 => conv_std_logic_vector(35571, 16),
54696 => conv_std_logic_vector(35784, 16),
54697 => conv_std_logic_vector(35997, 16),
54698 => conv_std_logic_vector(36210, 16),
54699 => conv_std_logic_vector(36423, 16),
54700 => conv_std_logic_vector(36636, 16),
54701 => conv_std_logic_vector(36849, 16),
54702 => conv_std_logic_vector(37062, 16),
54703 => conv_std_logic_vector(37275, 16),
54704 => conv_std_logic_vector(37488, 16),
54705 => conv_std_logic_vector(37701, 16),
54706 => conv_std_logic_vector(37914, 16),
54707 => conv_std_logic_vector(38127, 16),
54708 => conv_std_logic_vector(38340, 16),
54709 => conv_std_logic_vector(38553, 16),
54710 => conv_std_logic_vector(38766, 16),
54711 => conv_std_logic_vector(38979, 16),
54712 => conv_std_logic_vector(39192, 16),
54713 => conv_std_logic_vector(39405, 16),
54714 => conv_std_logic_vector(39618, 16),
54715 => conv_std_logic_vector(39831, 16),
54716 => conv_std_logic_vector(40044, 16),
54717 => conv_std_logic_vector(40257, 16),
54718 => conv_std_logic_vector(40470, 16),
54719 => conv_std_logic_vector(40683, 16),
54720 => conv_std_logic_vector(40896, 16),
54721 => conv_std_logic_vector(41109, 16),
54722 => conv_std_logic_vector(41322, 16),
54723 => conv_std_logic_vector(41535, 16),
54724 => conv_std_logic_vector(41748, 16),
54725 => conv_std_logic_vector(41961, 16),
54726 => conv_std_logic_vector(42174, 16),
54727 => conv_std_logic_vector(42387, 16),
54728 => conv_std_logic_vector(42600, 16),
54729 => conv_std_logic_vector(42813, 16),
54730 => conv_std_logic_vector(43026, 16),
54731 => conv_std_logic_vector(43239, 16),
54732 => conv_std_logic_vector(43452, 16),
54733 => conv_std_logic_vector(43665, 16),
54734 => conv_std_logic_vector(43878, 16),
54735 => conv_std_logic_vector(44091, 16),
54736 => conv_std_logic_vector(44304, 16),
54737 => conv_std_logic_vector(44517, 16),
54738 => conv_std_logic_vector(44730, 16),
54739 => conv_std_logic_vector(44943, 16),
54740 => conv_std_logic_vector(45156, 16),
54741 => conv_std_logic_vector(45369, 16),
54742 => conv_std_logic_vector(45582, 16),
54743 => conv_std_logic_vector(45795, 16),
54744 => conv_std_logic_vector(46008, 16),
54745 => conv_std_logic_vector(46221, 16),
54746 => conv_std_logic_vector(46434, 16),
54747 => conv_std_logic_vector(46647, 16),
54748 => conv_std_logic_vector(46860, 16),
54749 => conv_std_logic_vector(47073, 16),
54750 => conv_std_logic_vector(47286, 16),
54751 => conv_std_logic_vector(47499, 16),
54752 => conv_std_logic_vector(47712, 16),
54753 => conv_std_logic_vector(47925, 16),
54754 => conv_std_logic_vector(48138, 16),
54755 => conv_std_logic_vector(48351, 16),
54756 => conv_std_logic_vector(48564, 16),
54757 => conv_std_logic_vector(48777, 16),
54758 => conv_std_logic_vector(48990, 16),
54759 => conv_std_logic_vector(49203, 16),
54760 => conv_std_logic_vector(49416, 16),
54761 => conv_std_logic_vector(49629, 16),
54762 => conv_std_logic_vector(49842, 16),
54763 => conv_std_logic_vector(50055, 16),
54764 => conv_std_logic_vector(50268, 16),
54765 => conv_std_logic_vector(50481, 16),
54766 => conv_std_logic_vector(50694, 16),
54767 => conv_std_logic_vector(50907, 16),
54768 => conv_std_logic_vector(51120, 16),
54769 => conv_std_logic_vector(51333, 16),
54770 => conv_std_logic_vector(51546, 16),
54771 => conv_std_logic_vector(51759, 16),
54772 => conv_std_logic_vector(51972, 16),
54773 => conv_std_logic_vector(52185, 16),
54774 => conv_std_logic_vector(52398, 16),
54775 => conv_std_logic_vector(52611, 16),
54776 => conv_std_logic_vector(52824, 16),
54777 => conv_std_logic_vector(53037, 16),
54778 => conv_std_logic_vector(53250, 16),
54779 => conv_std_logic_vector(53463, 16),
54780 => conv_std_logic_vector(53676, 16),
54781 => conv_std_logic_vector(53889, 16),
54782 => conv_std_logic_vector(54102, 16),
54783 => conv_std_logic_vector(54315, 16),
54784 => conv_std_logic_vector(0, 16),
54785 => conv_std_logic_vector(214, 16),
54786 => conv_std_logic_vector(428, 16),
54787 => conv_std_logic_vector(642, 16),
54788 => conv_std_logic_vector(856, 16),
54789 => conv_std_logic_vector(1070, 16),
54790 => conv_std_logic_vector(1284, 16),
54791 => conv_std_logic_vector(1498, 16),
54792 => conv_std_logic_vector(1712, 16),
54793 => conv_std_logic_vector(1926, 16),
54794 => conv_std_logic_vector(2140, 16),
54795 => conv_std_logic_vector(2354, 16),
54796 => conv_std_logic_vector(2568, 16),
54797 => conv_std_logic_vector(2782, 16),
54798 => conv_std_logic_vector(2996, 16),
54799 => conv_std_logic_vector(3210, 16),
54800 => conv_std_logic_vector(3424, 16),
54801 => conv_std_logic_vector(3638, 16),
54802 => conv_std_logic_vector(3852, 16),
54803 => conv_std_logic_vector(4066, 16),
54804 => conv_std_logic_vector(4280, 16),
54805 => conv_std_logic_vector(4494, 16),
54806 => conv_std_logic_vector(4708, 16),
54807 => conv_std_logic_vector(4922, 16),
54808 => conv_std_logic_vector(5136, 16),
54809 => conv_std_logic_vector(5350, 16),
54810 => conv_std_logic_vector(5564, 16),
54811 => conv_std_logic_vector(5778, 16),
54812 => conv_std_logic_vector(5992, 16),
54813 => conv_std_logic_vector(6206, 16),
54814 => conv_std_logic_vector(6420, 16),
54815 => conv_std_logic_vector(6634, 16),
54816 => conv_std_logic_vector(6848, 16),
54817 => conv_std_logic_vector(7062, 16),
54818 => conv_std_logic_vector(7276, 16),
54819 => conv_std_logic_vector(7490, 16),
54820 => conv_std_logic_vector(7704, 16),
54821 => conv_std_logic_vector(7918, 16),
54822 => conv_std_logic_vector(8132, 16),
54823 => conv_std_logic_vector(8346, 16),
54824 => conv_std_logic_vector(8560, 16),
54825 => conv_std_logic_vector(8774, 16),
54826 => conv_std_logic_vector(8988, 16),
54827 => conv_std_logic_vector(9202, 16),
54828 => conv_std_logic_vector(9416, 16),
54829 => conv_std_logic_vector(9630, 16),
54830 => conv_std_logic_vector(9844, 16),
54831 => conv_std_logic_vector(10058, 16),
54832 => conv_std_logic_vector(10272, 16),
54833 => conv_std_logic_vector(10486, 16),
54834 => conv_std_logic_vector(10700, 16),
54835 => conv_std_logic_vector(10914, 16),
54836 => conv_std_logic_vector(11128, 16),
54837 => conv_std_logic_vector(11342, 16),
54838 => conv_std_logic_vector(11556, 16),
54839 => conv_std_logic_vector(11770, 16),
54840 => conv_std_logic_vector(11984, 16),
54841 => conv_std_logic_vector(12198, 16),
54842 => conv_std_logic_vector(12412, 16),
54843 => conv_std_logic_vector(12626, 16),
54844 => conv_std_logic_vector(12840, 16),
54845 => conv_std_logic_vector(13054, 16),
54846 => conv_std_logic_vector(13268, 16),
54847 => conv_std_logic_vector(13482, 16),
54848 => conv_std_logic_vector(13696, 16),
54849 => conv_std_logic_vector(13910, 16),
54850 => conv_std_logic_vector(14124, 16),
54851 => conv_std_logic_vector(14338, 16),
54852 => conv_std_logic_vector(14552, 16),
54853 => conv_std_logic_vector(14766, 16),
54854 => conv_std_logic_vector(14980, 16),
54855 => conv_std_logic_vector(15194, 16),
54856 => conv_std_logic_vector(15408, 16),
54857 => conv_std_logic_vector(15622, 16),
54858 => conv_std_logic_vector(15836, 16),
54859 => conv_std_logic_vector(16050, 16),
54860 => conv_std_logic_vector(16264, 16),
54861 => conv_std_logic_vector(16478, 16),
54862 => conv_std_logic_vector(16692, 16),
54863 => conv_std_logic_vector(16906, 16),
54864 => conv_std_logic_vector(17120, 16),
54865 => conv_std_logic_vector(17334, 16),
54866 => conv_std_logic_vector(17548, 16),
54867 => conv_std_logic_vector(17762, 16),
54868 => conv_std_logic_vector(17976, 16),
54869 => conv_std_logic_vector(18190, 16),
54870 => conv_std_logic_vector(18404, 16),
54871 => conv_std_logic_vector(18618, 16),
54872 => conv_std_logic_vector(18832, 16),
54873 => conv_std_logic_vector(19046, 16),
54874 => conv_std_logic_vector(19260, 16),
54875 => conv_std_logic_vector(19474, 16),
54876 => conv_std_logic_vector(19688, 16),
54877 => conv_std_logic_vector(19902, 16),
54878 => conv_std_logic_vector(20116, 16),
54879 => conv_std_logic_vector(20330, 16),
54880 => conv_std_logic_vector(20544, 16),
54881 => conv_std_logic_vector(20758, 16),
54882 => conv_std_logic_vector(20972, 16),
54883 => conv_std_logic_vector(21186, 16),
54884 => conv_std_logic_vector(21400, 16),
54885 => conv_std_logic_vector(21614, 16),
54886 => conv_std_logic_vector(21828, 16),
54887 => conv_std_logic_vector(22042, 16),
54888 => conv_std_logic_vector(22256, 16),
54889 => conv_std_logic_vector(22470, 16),
54890 => conv_std_logic_vector(22684, 16),
54891 => conv_std_logic_vector(22898, 16),
54892 => conv_std_logic_vector(23112, 16),
54893 => conv_std_logic_vector(23326, 16),
54894 => conv_std_logic_vector(23540, 16),
54895 => conv_std_logic_vector(23754, 16),
54896 => conv_std_logic_vector(23968, 16),
54897 => conv_std_logic_vector(24182, 16),
54898 => conv_std_logic_vector(24396, 16),
54899 => conv_std_logic_vector(24610, 16),
54900 => conv_std_logic_vector(24824, 16),
54901 => conv_std_logic_vector(25038, 16),
54902 => conv_std_logic_vector(25252, 16),
54903 => conv_std_logic_vector(25466, 16),
54904 => conv_std_logic_vector(25680, 16),
54905 => conv_std_logic_vector(25894, 16),
54906 => conv_std_logic_vector(26108, 16),
54907 => conv_std_logic_vector(26322, 16),
54908 => conv_std_logic_vector(26536, 16),
54909 => conv_std_logic_vector(26750, 16),
54910 => conv_std_logic_vector(26964, 16),
54911 => conv_std_logic_vector(27178, 16),
54912 => conv_std_logic_vector(27392, 16),
54913 => conv_std_logic_vector(27606, 16),
54914 => conv_std_logic_vector(27820, 16),
54915 => conv_std_logic_vector(28034, 16),
54916 => conv_std_logic_vector(28248, 16),
54917 => conv_std_logic_vector(28462, 16),
54918 => conv_std_logic_vector(28676, 16),
54919 => conv_std_logic_vector(28890, 16),
54920 => conv_std_logic_vector(29104, 16),
54921 => conv_std_logic_vector(29318, 16),
54922 => conv_std_logic_vector(29532, 16),
54923 => conv_std_logic_vector(29746, 16),
54924 => conv_std_logic_vector(29960, 16),
54925 => conv_std_logic_vector(30174, 16),
54926 => conv_std_logic_vector(30388, 16),
54927 => conv_std_logic_vector(30602, 16),
54928 => conv_std_logic_vector(30816, 16),
54929 => conv_std_logic_vector(31030, 16),
54930 => conv_std_logic_vector(31244, 16),
54931 => conv_std_logic_vector(31458, 16),
54932 => conv_std_logic_vector(31672, 16),
54933 => conv_std_logic_vector(31886, 16),
54934 => conv_std_logic_vector(32100, 16),
54935 => conv_std_logic_vector(32314, 16),
54936 => conv_std_logic_vector(32528, 16),
54937 => conv_std_logic_vector(32742, 16),
54938 => conv_std_logic_vector(32956, 16),
54939 => conv_std_logic_vector(33170, 16),
54940 => conv_std_logic_vector(33384, 16),
54941 => conv_std_logic_vector(33598, 16),
54942 => conv_std_logic_vector(33812, 16),
54943 => conv_std_logic_vector(34026, 16),
54944 => conv_std_logic_vector(34240, 16),
54945 => conv_std_logic_vector(34454, 16),
54946 => conv_std_logic_vector(34668, 16),
54947 => conv_std_logic_vector(34882, 16),
54948 => conv_std_logic_vector(35096, 16),
54949 => conv_std_logic_vector(35310, 16),
54950 => conv_std_logic_vector(35524, 16),
54951 => conv_std_logic_vector(35738, 16),
54952 => conv_std_logic_vector(35952, 16),
54953 => conv_std_logic_vector(36166, 16),
54954 => conv_std_logic_vector(36380, 16),
54955 => conv_std_logic_vector(36594, 16),
54956 => conv_std_logic_vector(36808, 16),
54957 => conv_std_logic_vector(37022, 16),
54958 => conv_std_logic_vector(37236, 16),
54959 => conv_std_logic_vector(37450, 16),
54960 => conv_std_logic_vector(37664, 16),
54961 => conv_std_logic_vector(37878, 16),
54962 => conv_std_logic_vector(38092, 16),
54963 => conv_std_logic_vector(38306, 16),
54964 => conv_std_logic_vector(38520, 16),
54965 => conv_std_logic_vector(38734, 16),
54966 => conv_std_logic_vector(38948, 16),
54967 => conv_std_logic_vector(39162, 16),
54968 => conv_std_logic_vector(39376, 16),
54969 => conv_std_logic_vector(39590, 16),
54970 => conv_std_logic_vector(39804, 16),
54971 => conv_std_logic_vector(40018, 16),
54972 => conv_std_logic_vector(40232, 16),
54973 => conv_std_logic_vector(40446, 16),
54974 => conv_std_logic_vector(40660, 16),
54975 => conv_std_logic_vector(40874, 16),
54976 => conv_std_logic_vector(41088, 16),
54977 => conv_std_logic_vector(41302, 16),
54978 => conv_std_logic_vector(41516, 16),
54979 => conv_std_logic_vector(41730, 16),
54980 => conv_std_logic_vector(41944, 16),
54981 => conv_std_logic_vector(42158, 16),
54982 => conv_std_logic_vector(42372, 16),
54983 => conv_std_logic_vector(42586, 16),
54984 => conv_std_logic_vector(42800, 16),
54985 => conv_std_logic_vector(43014, 16),
54986 => conv_std_logic_vector(43228, 16),
54987 => conv_std_logic_vector(43442, 16),
54988 => conv_std_logic_vector(43656, 16),
54989 => conv_std_logic_vector(43870, 16),
54990 => conv_std_logic_vector(44084, 16),
54991 => conv_std_logic_vector(44298, 16),
54992 => conv_std_logic_vector(44512, 16),
54993 => conv_std_logic_vector(44726, 16),
54994 => conv_std_logic_vector(44940, 16),
54995 => conv_std_logic_vector(45154, 16),
54996 => conv_std_logic_vector(45368, 16),
54997 => conv_std_logic_vector(45582, 16),
54998 => conv_std_logic_vector(45796, 16),
54999 => conv_std_logic_vector(46010, 16),
55000 => conv_std_logic_vector(46224, 16),
55001 => conv_std_logic_vector(46438, 16),
55002 => conv_std_logic_vector(46652, 16),
55003 => conv_std_logic_vector(46866, 16),
55004 => conv_std_logic_vector(47080, 16),
55005 => conv_std_logic_vector(47294, 16),
55006 => conv_std_logic_vector(47508, 16),
55007 => conv_std_logic_vector(47722, 16),
55008 => conv_std_logic_vector(47936, 16),
55009 => conv_std_logic_vector(48150, 16),
55010 => conv_std_logic_vector(48364, 16),
55011 => conv_std_logic_vector(48578, 16),
55012 => conv_std_logic_vector(48792, 16),
55013 => conv_std_logic_vector(49006, 16),
55014 => conv_std_logic_vector(49220, 16),
55015 => conv_std_logic_vector(49434, 16),
55016 => conv_std_logic_vector(49648, 16),
55017 => conv_std_logic_vector(49862, 16),
55018 => conv_std_logic_vector(50076, 16),
55019 => conv_std_logic_vector(50290, 16),
55020 => conv_std_logic_vector(50504, 16),
55021 => conv_std_logic_vector(50718, 16),
55022 => conv_std_logic_vector(50932, 16),
55023 => conv_std_logic_vector(51146, 16),
55024 => conv_std_logic_vector(51360, 16),
55025 => conv_std_logic_vector(51574, 16),
55026 => conv_std_logic_vector(51788, 16),
55027 => conv_std_logic_vector(52002, 16),
55028 => conv_std_logic_vector(52216, 16),
55029 => conv_std_logic_vector(52430, 16),
55030 => conv_std_logic_vector(52644, 16),
55031 => conv_std_logic_vector(52858, 16),
55032 => conv_std_logic_vector(53072, 16),
55033 => conv_std_logic_vector(53286, 16),
55034 => conv_std_logic_vector(53500, 16),
55035 => conv_std_logic_vector(53714, 16),
55036 => conv_std_logic_vector(53928, 16),
55037 => conv_std_logic_vector(54142, 16),
55038 => conv_std_logic_vector(54356, 16),
55039 => conv_std_logic_vector(54570, 16),
55040 => conv_std_logic_vector(0, 16),
55041 => conv_std_logic_vector(215, 16),
55042 => conv_std_logic_vector(430, 16),
55043 => conv_std_logic_vector(645, 16),
55044 => conv_std_logic_vector(860, 16),
55045 => conv_std_logic_vector(1075, 16),
55046 => conv_std_logic_vector(1290, 16),
55047 => conv_std_logic_vector(1505, 16),
55048 => conv_std_logic_vector(1720, 16),
55049 => conv_std_logic_vector(1935, 16),
55050 => conv_std_logic_vector(2150, 16),
55051 => conv_std_logic_vector(2365, 16),
55052 => conv_std_logic_vector(2580, 16),
55053 => conv_std_logic_vector(2795, 16),
55054 => conv_std_logic_vector(3010, 16),
55055 => conv_std_logic_vector(3225, 16),
55056 => conv_std_logic_vector(3440, 16),
55057 => conv_std_logic_vector(3655, 16),
55058 => conv_std_logic_vector(3870, 16),
55059 => conv_std_logic_vector(4085, 16),
55060 => conv_std_logic_vector(4300, 16),
55061 => conv_std_logic_vector(4515, 16),
55062 => conv_std_logic_vector(4730, 16),
55063 => conv_std_logic_vector(4945, 16),
55064 => conv_std_logic_vector(5160, 16),
55065 => conv_std_logic_vector(5375, 16),
55066 => conv_std_logic_vector(5590, 16),
55067 => conv_std_logic_vector(5805, 16),
55068 => conv_std_logic_vector(6020, 16),
55069 => conv_std_logic_vector(6235, 16),
55070 => conv_std_logic_vector(6450, 16),
55071 => conv_std_logic_vector(6665, 16),
55072 => conv_std_logic_vector(6880, 16),
55073 => conv_std_logic_vector(7095, 16),
55074 => conv_std_logic_vector(7310, 16),
55075 => conv_std_logic_vector(7525, 16),
55076 => conv_std_logic_vector(7740, 16),
55077 => conv_std_logic_vector(7955, 16),
55078 => conv_std_logic_vector(8170, 16),
55079 => conv_std_logic_vector(8385, 16),
55080 => conv_std_logic_vector(8600, 16),
55081 => conv_std_logic_vector(8815, 16),
55082 => conv_std_logic_vector(9030, 16),
55083 => conv_std_logic_vector(9245, 16),
55084 => conv_std_logic_vector(9460, 16),
55085 => conv_std_logic_vector(9675, 16),
55086 => conv_std_logic_vector(9890, 16),
55087 => conv_std_logic_vector(10105, 16),
55088 => conv_std_logic_vector(10320, 16),
55089 => conv_std_logic_vector(10535, 16),
55090 => conv_std_logic_vector(10750, 16),
55091 => conv_std_logic_vector(10965, 16),
55092 => conv_std_logic_vector(11180, 16),
55093 => conv_std_logic_vector(11395, 16),
55094 => conv_std_logic_vector(11610, 16),
55095 => conv_std_logic_vector(11825, 16),
55096 => conv_std_logic_vector(12040, 16),
55097 => conv_std_logic_vector(12255, 16),
55098 => conv_std_logic_vector(12470, 16),
55099 => conv_std_logic_vector(12685, 16),
55100 => conv_std_logic_vector(12900, 16),
55101 => conv_std_logic_vector(13115, 16),
55102 => conv_std_logic_vector(13330, 16),
55103 => conv_std_logic_vector(13545, 16),
55104 => conv_std_logic_vector(13760, 16),
55105 => conv_std_logic_vector(13975, 16),
55106 => conv_std_logic_vector(14190, 16),
55107 => conv_std_logic_vector(14405, 16),
55108 => conv_std_logic_vector(14620, 16),
55109 => conv_std_logic_vector(14835, 16),
55110 => conv_std_logic_vector(15050, 16),
55111 => conv_std_logic_vector(15265, 16),
55112 => conv_std_logic_vector(15480, 16),
55113 => conv_std_logic_vector(15695, 16),
55114 => conv_std_logic_vector(15910, 16),
55115 => conv_std_logic_vector(16125, 16),
55116 => conv_std_logic_vector(16340, 16),
55117 => conv_std_logic_vector(16555, 16),
55118 => conv_std_logic_vector(16770, 16),
55119 => conv_std_logic_vector(16985, 16),
55120 => conv_std_logic_vector(17200, 16),
55121 => conv_std_logic_vector(17415, 16),
55122 => conv_std_logic_vector(17630, 16),
55123 => conv_std_logic_vector(17845, 16),
55124 => conv_std_logic_vector(18060, 16),
55125 => conv_std_logic_vector(18275, 16),
55126 => conv_std_logic_vector(18490, 16),
55127 => conv_std_logic_vector(18705, 16),
55128 => conv_std_logic_vector(18920, 16),
55129 => conv_std_logic_vector(19135, 16),
55130 => conv_std_logic_vector(19350, 16),
55131 => conv_std_logic_vector(19565, 16),
55132 => conv_std_logic_vector(19780, 16),
55133 => conv_std_logic_vector(19995, 16),
55134 => conv_std_logic_vector(20210, 16),
55135 => conv_std_logic_vector(20425, 16),
55136 => conv_std_logic_vector(20640, 16),
55137 => conv_std_logic_vector(20855, 16),
55138 => conv_std_logic_vector(21070, 16),
55139 => conv_std_logic_vector(21285, 16),
55140 => conv_std_logic_vector(21500, 16),
55141 => conv_std_logic_vector(21715, 16),
55142 => conv_std_logic_vector(21930, 16),
55143 => conv_std_logic_vector(22145, 16),
55144 => conv_std_logic_vector(22360, 16),
55145 => conv_std_logic_vector(22575, 16),
55146 => conv_std_logic_vector(22790, 16),
55147 => conv_std_logic_vector(23005, 16),
55148 => conv_std_logic_vector(23220, 16),
55149 => conv_std_logic_vector(23435, 16),
55150 => conv_std_logic_vector(23650, 16),
55151 => conv_std_logic_vector(23865, 16),
55152 => conv_std_logic_vector(24080, 16),
55153 => conv_std_logic_vector(24295, 16),
55154 => conv_std_logic_vector(24510, 16),
55155 => conv_std_logic_vector(24725, 16),
55156 => conv_std_logic_vector(24940, 16),
55157 => conv_std_logic_vector(25155, 16),
55158 => conv_std_logic_vector(25370, 16),
55159 => conv_std_logic_vector(25585, 16),
55160 => conv_std_logic_vector(25800, 16),
55161 => conv_std_logic_vector(26015, 16),
55162 => conv_std_logic_vector(26230, 16),
55163 => conv_std_logic_vector(26445, 16),
55164 => conv_std_logic_vector(26660, 16),
55165 => conv_std_logic_vector(26875, 16),
55166 => conv_std_logic_vector(27090, 16),
55167 => conv_std_logic_vector(27305, 16),
55168 => conv_std_logic_vector(27520, 16),
55169 => conv_std_logic_vector(27735, 16),
55170 => conv_std_logic_vector(27950, 16),
55171 => conv_std_logic_vector(28165, 16),
55172 => conv_std_logic_vector(28380, 16),
55173 => conv_std_logic_vector(28595, 16),
55174 => conv_std_logic_vector(28810, 16),
55175 => conv_std_logic_vector(29025, 16),
55176 => conv_std_logic_vector(29240, 16),
55177 => conv_std_logic_vector(29455, 16),
55178 => conv_std_logic_vector(29670, 16),
55179 => conv_std_logic_vector(29885, 16),
55180 => conv_std_logic_vector(30100, 16),
55181 => conv_std_logic_vector(30315, 16),
55182 => conv_std_logic_vector(30530, 16),
55183 => conv_std_logic_vector(30745, 16),
55184 => conv_std_logic_vector(30960, 16),
55185 => conv_std_logic_vector(31175, 16),
55186 => conv_std_logic_vector(31390, 16),
55187 => conv_std_logic_vector(31605, 16),
55188 => conv_std_logic_vector(31820, 16),
55189 => conv_std_logic_vector(32035, 16),
55190 => conv_std_logic_vector(32250, 16),
55191 => conv_std_logic_vector(32465, 16),
55192 => conv_std_logic_vector(32680, 16),
55193 => conv_std_logic_vector(32895, 16),
55194 => conv_std_logic_vector(33110, 16),
55195 => conv_std_logic_vector(33325, 16),
55196 => conv_std_logic_vector(33540, 16),
55197 => conv_std_logic_vector(33755, 16),
55198 => conv_std_logic_vector(33970, 16),
55199 => conv_std_logic_vector(34185, 16),
55200 => conv_std_logic_vector(34400, 16),
55201 => conv_std_logic_vector(34615, 16),
55202 => conv_std_logic_vector(34830, 16),
55203 => conv_std_logic_vector(35045, 16),
55204 => conv_std_logic_vector(35260, 16),
55205 => conv_std_logic_vector(35475, 16),
55206 => conv_std_logic_vector(35690, 16),
55207 => conv_std_logic_vector(35905, 16),
55208 => conv_std_logic_vector(36120, 16),
55209 => conv_std_logic_vector(36335, 16),
55210 => conv_std_logic_vector(36550, 16),
55211 => conv_std_logic_vector(36765, 16),
55212 => conv_std_logic_vector(36980, 16),
55213 => conv_std_logic_vector(37195, 16),
55214 => conv_std_logic_vector(37410, 16),
55215 => conv_std_logic_vector(37625, 16),
55216 => conv_std_logic_vector(37840, 16),
55217 => conv_std_logic_vector(38055, 16),
55218 => conv_std_logic_vector(38270, 16),
55219 => conv_std_logic_vector(38485, 16),
55220 => conv_std_logic_vector(38700, 16),
55221 => conv_std_logic_vector(38915, 16),
55222 => conv_std_logic_vector(39130, 16),
55223 => conv_std_logic_vector(39345, 16),
55224 => conv_std_logic_vector(39560, 16),
55225 => conv_std_logic_vector(39775, 16),
55226 => conv_std_logic_vector(39990, 16),
55227 => conv_std_logic_vector(40205, 16),
55228 => conv_std_logic_vector(40420, 16),
55229 => conv_std_logic_vector(40635, 16),
55230 => conv_std_logic_vector(40850, 16),
55231 => conv_std_logic_vector(41065, 16),
55232 => conv_std_logic_vector(41280, 16),
55233 => conv_std_logic_vector(41495, 16),
55234 => conv_std_logic_vector(41710, 16),
55235 => conv_std_logic_vector(41925, 16),
55236 => conv_std_logic_vector(42140, 16),
55237 => conv_std_logic_vector(42355, 16),
55238 => conv_std_logic_vector(42570, 16),
55239 => conv_std_logic_vector(42785, 16),
55240 => conv_std_logic_vector(43000, 16),
55241 => conv_std_logic_vector(43215, 16),
55242 => conv_std_logic_vector(43430, 16),
55243 => conv_std_logic_vector(43645, 16),
55244 => conv_std_logic_vector(43860, 16),
55245 => conv_std_logic_vector(44075, 16),
55246 => conv_std_logic_vector(44290, 16),
55247 => conv_std_logic_vector(44505, 16),
55248 => conv_std_logic_vector(44720, 16),
55249 => conv_std_logic_vector(44935, 16),
55250 => conv_std_logic_vector(45150, 16),
55251 => conv_std_logic_vector(45365, 16),
55252 => conv_std_logic_vector(45580, 16),
55253 => conv_std_logic_vector(45795, 16),
55254 => conv_std_logic_vector(46010, 16),
55255 => conv_std_logic_vector(46225, 16),
55256 => conv_std_logic_vector(46440, 16),
55257 => conv_std_logic_vector(46655, 16),
55258 => conv_std_logic_vector(46870, 16),
55259 => conv_std_logic_vector(47085, 16),
55260 => conv_std_logic_vector(47300, 16),
55261 => conv_std_logic_vector(47515, 16),
55262 => conv_std_logic_vector(47730, 16),
55263 => conv_std_logic_vector(47945, 16),
55264 => conv_std_logic_vector(48160, 16),
55265 => conv_std_logic_vector(48375, 16),
55266 => conv_std_logic_vector(48590, 16),
55267 => conv_std_logic_vector(48805, 16),
55268 => conv_std_logic_vector(49020, 16),
55269 => conv_std_logic_vector(49235, 16),
55270 => conv_std_logic_vector(49450, 16),
55271 => conv_std_logic_vector(49665, 16),
55272 => conv_std_logic_vector(49880, 16),
55273 => conv_std_logic_vector(50095, 16),
55274 => conv_std_logic_vector(50310, 16),
55275 => conv_std_logic_vector(50525, 16),
55276 => conv_std_logic_vector(50740, 16),
55277 => conv_std_logic_vector(50955, 16),
55278 => conv_std_logic_vector(51170, 16),
55279 => conv_std_logic_vector(51385, 16),
55280 => conv_std_logic_vector(51600, 16),
55281 => conv_std_logic_vector(51815, 16),
55282 => conv_std_logic_vector(52030, 16),
55283 => conv_std_logic_vector(52245, 16),
55284 => conv_std_logic_vector(52460, 16),
55285 => conv_std_logic_vector(52675, 16),
55286 => conv_std_logic_vector(52890, 16),
55287 => conv_std_logic_vector(53105, 16),
55288 => conv_std_logic_vector(53320, 16),
55289 => conv_std_logic_vector(53535, 16),
55290 => conv_std_logic_vector(53750, 16),
55291 => conv_std_logic_vector(53965, 16),
55292 => conv_std_logic_vector(54180, 16),
55293 => conv_std_logic_vector(54395, 16),
55294 => conv_std_logic_vector(54610, 16),
55295 => conv_std_logic_vector(54825, 16),
55296 => conv_std_logic_vector(0, 16),
55297 => conv_std_logic_vector(216, 16),
55298 => conv_std_logic_vector(432, 16),
55299 => conv_std_logic_vector(648, 16),
55300 => conv_std_logic_vector(864, 16),
55301 => conv_std_logic_vector(1080, 16),
55302 => conv_std_logic_vector(1296, 16),
55303 => conv_std_logic_vector(1512, 16),
55304 => conv_std_logic_vector(1728, 16),
55305 => conv_std_logic_vector(1944, 16),
55306 => conv_std_logic_vector(2160, 16),
55307 => conv_std_logic_vector(2376, 16),
55308 => conv_std_logic_vector(2592, 16),
55309 => conv_std_logic_vector(2808, 16),
55310 => conv_std_logic_vector(3024, 16),
55311 => conv_std_logic_vector(3240, 16),
55312 => conv_std_logic_vector(3456, 16),
55313 => conv_std_logic_vector(3672, 16),
55314 => conv_std_logic_vector(3888, 16),
55315 => conv_std_logic_vector(4104, 16),
55316 => conv_std_logic_vector(4320, 16),
55317 => conv_std_logic_vector(4536, 16),
55318 => conv_std_logic_vector(4752, 16),
55319 => conv_std_logic_vector(4968, 16),
55320 => conv_std_logic_vector(5184, 16),
55321 => conv_std_logic_vector(5400, 16),
55322 => conv_std_logic_vector(5616, 16),
55323 => conv_std_logic_vector(5832, 16),
55324 => conv_std_logic_vector(6048, 16),
55325 => conv_std_logic_vector(6264, 16),
55326 => conv_std_logic_vector(6480, 16),
55327 => conv_std_logic_vector(6696, 16),
55328 => conv_std_logic_vector(6912, 16),
55329 => conv_std_logic_vector(7128, 16),
55330 => conv_std_logic_vector(7344, 16),
55331 => conv_std_logic_vector(7560, 16),
55332 => conv_std_logic_vector(7776, 16),
55333 => conv_std_logic_vector(7992, 16),
55334 => conv_std_logic_vector(8208, 16),
55335 => conv_std_logic_vector(8424, 16),
55336 => conv_std_logic_vector(8640, 16),
55337 => conv_std_logic_vector(8856, 16),
55338 => conv_std_logic_vector(9072, 16),
55339 => conv_std_logic_vector(9288, 16),
55340 => conv_std_logic_vector(9504, 16),
55341 => conv_std_logic_vector(9720, 16),
55342 => conv_std_logic_vector(9936, 16),
55343 => conv_std_logic_vector(10152, 16),
55344 => conv_std_logic_vector(10368, 16),
55345 => conv_std_logic_vector(10584, 16),
55346 => conv_std_logic_vector(10800, 16),
55347 => conv_std_logic_vector(11016, 16),
55348 => conv_std_logic_vector(11232, 16),
55349 => conv_std_logic_vector(11448, 16),
55350 => conv_std_logic_vector(11664, 16),
55351 => conv_std_logic_vector(11880, 16),
55352 => conv_std_logic_vector(12096, 16),
55353 => conv_std_logic_vector(12312, 16),
55354 => conv_std_logic_vector(12528, 16),
55355 => conv_std_logic_vector(12744, 16),
55356 => conv_std_logic_vector(12960, 16),
55357 => conv_std_logic_vector(13176, 16),
55358 => conv_std_logic_vector(13392, 16),
55359 => conv_std_logic_vector(13608, 16),
55360 => conv_std_logic_vector(13824, 16),
55361 => conv_std_logic_vector(14040, 16),
55362 => conv_std_logic_vector(14256, 16),
55363 => conv_std_logic_vector(14472, 16),
55364 => conv_std_logic_vector(14688, 16),
55365 => conv_std_logic_vector(14904, 16),
55366 => conv_std_logic_vector(15120, 16),
55367 => conv_std_logic_vector(15336, 16),
55368 => conv_std_logic_vector(15552, 16),
55369 => conv_std_logic_vector(15768, 16),
55370 => conv_std_logic_vector(15984, 16),
55371 => conv_std_logic_vector(16200, 16),
55372 => conv_std_logic_vector(16416, 16),
55373 => conv_std_logic_vector(16632, 16),
55374 => conv_std_logic_vector(16848, 16),
55375 => conv_std_logic_vector(17064, 16),
55376 => conv_std_logic_vector(17280, 16),
55377 => conv_std_logic_vector(17496, 16),
55378 => conv_std_logic_vector(17712, 16),
55379 => conv_std_logic_vector(17928, 16),
55380 => conv_std_logic_vector(18144, 16),
55381 => conv_std_logic_vector(18360, 16),
55382 => conv_std_logic_vector(18576, 16),
55383 => conv_std_logic_vector(18792, 16),
55384 => conv_std_logic_vector(19008, 16),
55385 => conv_std_logic_vector(19224, 16),
55386 => conv_std_logic_vector(19440, 16),
55387 => conv_std_logic_vector(19656, 16),
55388 => conv_std_logic_vector(19872, 16),
55389 => conv_std_logic_vector(20088, 16),
55390 => conv_std_logic_vector(20304, 16),
55391 => conv_std_logic_vector(20520, 16),
55392 => conv_std_logic_vector(20736, 16),
55393 => conv_std_logic_vector(20952, 16),
55394 => conv_std_logic_vector(21168, 16),
55395 => conv_std_logic_vector(21384, 16),
55396 => conv_std_logic_vector(21600, 16),
55397 => conv_std_logic_vector(21816, 16),
55398 => conv_std_logic_vector(22032, 16),
55399 => conv_std_logic_vector(22248, 16),
55400 => conv_std_logic_vector(22464, 16),
55401 => conv_std_logic_vector(22680, 16),
55402 => conv_std_logic_vector(22896, 16),
55403 => conv_std_logic_vector(23112, 16),
55404 => conv_std_logic_vector(23328, 16),
55405 => conv_std_logic_vector(23544, 16),
55406 => conv_std_logic_vector(23760, 16),
55407 => conv_std_logic_vector(23976, 16),
55408 => conv_std_logic_vector(24192, 16),
55409 => conv_std_logic_vector(24408, 16),
55410 => conv_std_logic_vector(24624, 16),
55411 => conv_std_logic_vector(24840, 16),
55412 => conv_std_logic_vector(25056, 16),
55413 => conv_std_logic_vector(25272, 16),
55414 => conv_std_logic_vector(25488, 16),
55415 => conv_std_logic_vector(25704, 16),
55416 => conv_std_logic_vector(25920, 16),
55417 => conv_std_logic_vector(26136, 16),
55418 => conv_std_logic_vector(26352, 16),
55419 => conv_std_logic_vector(26568, 16),
55420 => conv_std_logic_vector(26784, 16),
55421 => conv_std_logic_vector(27000, 16),
55422 => conv_std_logic_vector(27216, 16),
55423 => conv_std_logic_vector(27432, 16),
55424 => conv_std_logic_vector(27648, 16),
55425 => conv_std_logic_vector(27864, 16),
55426 => conv_std_logic_vector(28080, 16),
55427 => conv_std_logic_vector(28296, 16),
55428 => conv_std_logic_vector(28512, 16),
55429 => conv_std_logic_vector(28728, 16),
55430 => conv_std_logic_vector(28944, 16),
55431 => conv_std_logic_vector(29160, 16),
55432 => conv_std_logic_vector(29376, 16),
55433 => conv_std_logic_vector(29592, 16),
55434 => conv_std_logic_vector(29808, 16),
55435 => conv_std_logic_vector(30024, 16),
55436 => conv_std_logic_vector(30240, 16),
55437 => conv_std_logic_vector(30456, 16),
55438 => conv_std_logic_vector(30672, 16),
55439 => conv_std_logic_vector(30888, 16),
55440 => conv_std_logic_vector(31104, 16),
55441 => conv_std_logic_vector(31320, 16),
55442 => conv_std_logic_vector(31536, 16),
55443 => conv_std_logic_vector(31752, 16),
55444 => conv_std_logic_vector(31968, 16),
55445 => conv_std_logic_vector(32184, 16),
55446 => conv_std_logic_vector(32400, 16),
55447 => conv_std_logic_vector(32616, 16),
55448 => conv_std_logic_vector(32832, 16),
55449 => conv_std_logic_vector(33048, 16),
55450 => conv_std_logic_vector(33264, 16),
55451 => conv_std_logic_vector(33480, 16),
55452 => conv_std_logic_vector(33696, 16),
55453 => conv_std_logic_vector(33912, 16),
55454 => conv_std_logic_vector(34128, 16),
55455 => conv_std_logic_vector(34344, 16),
55456 => conv_std_logic_vector(34560, 16),
55457 => conv_std_logic_vector(34776, 16),
55458 => conv_std_logic_vector(34992, 16),
55459 => conv_std_logic_vector(35208, 16),
55460 => conv_std_logic_vector(35424, 16),
55461 => conv_std_logic_vector(35640, 16),
55462 => conv_std_logic_vector(35856, 16),
55463 => conv_std_logic_vector(36072, 16),
55464 => conv_std_logic_vector(36288, 16),
55465 => conv_std_logic_vector(36504, 16),
55466 => conv_std_logic_vector(36720, 16),
55467 => conv_std_logic_vector(36936, 16),
55468 => conv_std_logic_vector(37152, 16),
55469 => conv_std_logic_vector(37368, 16),
55470 => conv_std_logic_vector(37584, 16),
55471 => conv_std_logic_vector(37800, 16),
55472 => conv_std_logic_vector(38016, 16),
55473 => conv_std_logic_vector(38232, 16),
55474 => conv_std_logic_vector(38448, 16),
55475 => conv_std_logic_vector(38664, 16),
55476 => conv_std_logic_vector(38880, 16),
55477 => conv_std_logic_vector(39096, 16),
55478 => conv_std_logic_vector(39312, 16),
55479 => conv_std_logic_vector(39528, 16),
55480 => conv_std_logic_vector(39744, 16),
55481 => conv_std_logic_vector(39960, 16),
55482 => conv_std_logic_vector(40176, 16),
55483 => conv_std_logic_vector(40392, 16),
55484 => conv_std_logic_vector(40608, 16),
55485 => conv_std_logic_vector(40824, 16),
55486 => conv_std_logic_vector(41040, 16),
55487 => conv_std_logic_vector(41256, 16),
55488 => conv_std_logic_vector(41472, 16),
55489 => conv_std_logic_vector(41688, 16),
55490 => conv_std_logic_vector(41904, 16),
55491 => conv_std_logic_vector(42120, 16),
55492 => conv_std_logic_vector(42336, 16),
55493 => conv_std_logic_vector(42552, 16),
55494 => conv_std_logic_vector(42768, 16),
55495 => conv_std_logic_vector(42984, 16),
55496 => conv_std_logic_vector(43200, 16),
55497 => conv_std_logic_vector(43416, 16),
55498 => conv_std_logic_vector(43632, 16),
55499 => conv_std_logic_vector(43848, 16),
55500 => conv_std_logic_vector(44064, 16),
55501 => conv_std_logic_vector(44280, 16),
55502 => conv_std_logic_vector(44496, 16),
55503 => conv_std_logic_vector(44712, 16),
55504 => conv_std_logic_vector(44928, 16),
55505 => conv_std_logic_vector(45144, 16),
55506 => conv_std_logic_vector(45360, 16),
55507 => conv_std_logic_vector(45576, 16),
55508 => conv_std_logic_vector(45792, 16),
55509 => conv_std_logic_vector(46008, 16),
55510 => conv_std_logic_vector(46224, 16),
55511 => conv_std_logic_vector(46440, 16),
55512 => conv_std_logic_vector(46656, 16),
55513 => conv_std_logic_vector(46872, 16),
55514 => conv_std_logic_vector(47088, 16),
55515 => conv_std_logic_vector(47304, 16),
55516 => conv_std_logic_vector(47520, 16),
55517 => conv_std_logic_vector(47736, 16),
55518 => conv_std_logic_vector(47952, 16),
55519 => conv_std_logic_vector(48168, 16),
55520 => conv_std_logic_vector(48384, 16),
55521 => conv_std_logic_vector(48600, 16),
55522 => conv_std_logic_vector(48816, 16),
55523 => conv_std_logic_vector(49032, 16),
55524 => conv_std_logic_vector(49248, 16),
55525 => conv_std_logic_vector(49464, 16),
55526 => conv_std_logic_vector(49680, 16),
55527 => conv_std_logic_vector(49896, 16),
55528 => conv_std_logic_vector(50112, 16),
55529 => conv_std_logic_vector(50328, 16),
55530 => conv_std_logic_vector(50544, 16),
55531 => conv_std_logic_vector(50760, 16),
55532 => conv_std_logic_vector(50976, 16),
55533 => conv_std_logic_vector(51192, 16),
55534 => conv_std_logic_vector(51408, 16),
55535 => conv_std_logic_vector(51624, 16),
55536 => conv_std_logic_vector(51840, 16),
55537 => conv_std_logic_vector(52056, 16),
55538 => conv_std_logic_vector(52272, 16),
55539 => conv_std_logic_vector(52488, 16),
55540 => conv_std_logic_vector(52704, 16),
55541 => conv_std_logic_vector(52920, 16),
55542 => conv_std_logic_vector(53136, 16),
55543 => conv_std_logic_vector(53352, 16),
55544 => conv_std_logic_vector(53568, 16),
55545 => conv_std_logic_vector(53784, 16),
55546 => conv_std_logic_vector(54000, 16),
55547 => conv_std_logic_vector(54216, 16),
55548 => conv_std_logic_vector(54432, 16),
55549 => conv_std_logic_vector(54648, 16),
55550 => conv_std_logic_vector(54864, 16),
55551 => conv_std_logic_vector(55080, 16),
55552 => conv_std_logic_vector(0, 16),
55553 => conv_std_logic_vector(217, 16),
55554 => conv_std_logic_vector(434, 16),
55555 => conv_std_logic_vector(651, 16),
55556 => conv_std_logic_vector(868, 16),
55557 => conv_std_logic_vector(1085, 16),
55558 => conv_std_logic_vector(1302, 16),
55559 => conv_std_logic_vector(1519, 16),
55560 => conv_std_logic_vector(1736, 16),
55561 => conv_std_logic_vector(1953, 16),
55562 => conv_std_logic_vector(2170, 16),
55563 => conv_std_logic_vector(2387, 16),
55564 => conv_std_logic_vector(2604, 16),
55565 => conv_std_logic_vector(2821, 16),
55566 => conv_std_logic_vector(3038, 16),
55567 => conv_std_logic_vector(3255, 16),
55568 => conv_std_logic_vector(3472, 16),
55569 => conv_std_logic_vector(3689, 16),
55570 => conv_std_logic_vector(3906, 16),
55571 => conv_std_logic_vector(4123, 16),
55572 => conv_std_logic_vector(4340, 16),
55573 => conv_std_logic_vector(4557, 16),
55574 => conv_std_logic_vector(4774, 16),
55575 => conv_std_logic_vector(4991, 16),
55576 => conv_std_logic_vector(5208, 16),
55577 => conv_std_logic_vector(5425, 16),
55578 => conv_std_logic_vector(5642, 16),
55579 => conv_std_logic_vector(5859, 16),
55580 => conv_std_logic_vector(6076, 16),
55581 => conv_std_logic_vector(6293, 16),
55582 => conv_std_logic_vector(6510, 16),
55583 => conv_std_logic_vector(6727, 16),
55584 => conv_std_logic_vector(6944, 16),
55585 => conv_std_logic_vector(7161, 16),
55586 => conv_std_logic_vector(7378, 16),
55587 => conv_std_logic_vector(7595, 16),
55588 => conv_std_logic_vector(7812, 16),
55589 => conv_std_logic_vector(8029, 16),
55590 => conv_std_logic_vector(8246, 16),
55591 => conv_std_logic_vector(8463, 16),
55592 => conv_std_logic_vector(8680, 16),
55593 => conv_std_logic_vector(8897, 16),
55594 => conv_std_logic_vector(9114, 16),
55595 => conv_std_logic_vector(9331, 16),
55596 => conv_std_logic_vector(9548, 16),
55597 => conv_std_logic_vector(9765, 16),
55598 => conv_std_logic_vector(9982, 16),
55599 => conv_std_logic_vector(10199, 16),
55600 => conv_std_logic_vector(10416, 16),
55601 => conv_std_logic_vector(10633, 16),
55602 => conv_std_logic_vector(10850, 16),
55603 => conv_std_logic_vector(11067, 16),
55604 => conv_std_logic_vector(11284, 16),
55605 => conv_std_logic_vector(11501, 16),
55606 => conv_std_logic_vector(11718, 16),
55607 => conv_std_logic_vector(11935, 16),
55608 => conv_std_logic_vector(12152, 16),
55609 => conv_std_logic_vector(12369, 16),
55610 => conv_std_logic_vector(12586, 16),
55611 => conv_std_logic_vector(12803, 16),
55612 => conv_std_logic_vector(13020, 16),
55613 => conv_std_logic_vector(13237, 16),
55614 => conv_std_logic_vector(13454, 16),
55615 => conv_std_logic_vector(13671, 16),
55616 => conv_std_logic_vector(13888, 16),
55617 => conv_std_logic_vector(14105, 16),
55618 => conv_std_logic_vector(14322, 16),
55619 => conv_std_logic_vector(14539, 16),
55620 => conv_std_logic_vector(14756, 16),
55621 => conv_std_logic_vector(14973, 16),
55622 => conv_std_logic_vector(15190, 16),
55623 => conv_std_logic_vector(15407, 16),
55624 => conv_std_logic_vector(15624, 16),
55625 => conv_std_logic_vector(15841, 16),
55626 => conv_std_logic_vector(16058, 16),
55627 => conv_std_logic_vector(16275, 16),
55628 => conv_std_logic_vector(16492, 16),
55629 => conv_std_logic_vector(16709, 16),
55630 => conv_std_logic_vector(16926, 16),
55631 => conv_std_logic_vector(17143, 16),
55632 => conv_std_logic_vector(17360, 16),
55633 => conv_std_logic_vector(17577, 16),
55634 => conv_std_logic_vector(17794, 16),
55635 => conv_std_logic_vector(18011, 16),
55636 => conv_std_logic_vector(18228, 16),
55637 => conv_std_logic_vector(18445, 16),
55638 => conv_std_logic_vector(18662, 16),
55639 => conv_std_logic_vector(18879, 16),
55640 => conv_std_logic_vector(19096, 16),
55641 => conv_std_logic_vector(19313, 16),
55642 => conv_std_logic_vector(19530, 16),
55643 => conv_std_logic_vector(19747, 16),
55644 => conv_std_logic_vector(19964, 16),
55645 => conv_std_logic_vector(20181, 16),
55646 => conv_std_logic_vector(20398, 16),
55647 => conv_std_logic_vector(20615, 16),
55648 => conv_std_logic_vector(20832, 16),
55649 => conv_std_logic_vector(21049, 16),
55650 => conv_std_logic_vector(21266, 16),
55651 => conv_std_logic_vector(21483, 16),
55652 => conv_std_logic_vector(21700, 16),
55653 => conv_std_logic_vector(21917, 16),
55654 => conv_std_logic_vector(22134, 16),
55655 => conv_std_logic_vector(22351, 16),
55656 => conv_std_logic_vector(22568, 16),
55657 => conv_std_logic_vector(22785, 16),
55658 => conv_std_logic_vector(23002, 16),
55659 => conv_std_logic_vector(23219, 16),
55660 => conv_std_logic_vector(23436, 16),
55661 => conv_std_logic_vector(23653, 16),
55662 => conv_std_logic_vector(23870, 16),
55663 => conv_std_logic_vector(24087, 16),
55664 => conv_std_logic_vector(24304, 16),
55665 => conv_std_logic_vector(24521, 16),
55666 => conv_std_logic_vector(24738, 16),
55667 => conv_std_logic_vector(24955, 16),
55668 => conv_std_logic_vector(25172, 16),
55669 => conv_std_logic_vector(25389, 16),
55670 => conv_std_logic_vector(25606, 16),
55671 => conv_std_logic_vector(25823, 16),
55672 => conv_std_logic_vector(26040, 16),
55673 => conv_std_logic_vector(26257, 16),
55674 => conv_std_logic_vector(26474, 16),
55675 => conv_std_logic_vector(26691, 16),
55676 => conv_std_logic_vector(26908, 16),
55677 => conv_std_logic_vector(27125, 16),
55678 => conv_std_logic_vector(27342, 16),
55679 => conv_std_logic_vector(27559, 16),
55680 => conv_std_logic_vector(27776, 16),
55681 => conv_std_logic_vector(27993, 16),
55682 => conv_std_logic_vector(28210, 16),
55683 => conv_std_logic_vector(28427, 16),
55684 => conv_std_logic_vector(28644, 16),
55685 => conv_std_logic_vector(28861, 16),
55686 => conv_std_logic_vector(29078, 16),
55687 => conv_std_logic_vector(29295, 16),
55688 => conv_std_logic_vector(29512, 16),
55689 => conv_std_logic_vector(29729, 16),
55690 => conv_std_logic_vector(29946, 16),
55691 => conv_std_logic_vector(30163, 16),
55692 => conv_std_logic_vector(30380, 16),
55693 => conv_std_logic_vector(30597, 16),
55694 => conv_std_logic_vector(30814, 16),
55695 => conv_std_logic_vector(31031, 16),
55696 => conv_std_logic_vector(31248, 16),
55697 => conv_std_logic_vector(31465, 16),
55698 => conv_std_logic_vector(31682, 16),
55699 => conv_std_logic_vector(31899, 16),
55700 => conv_std_logic_vector(32116, 16),
55701 => conv_std_logic_vector(32333, 16),
55702 => conv_std_logic_vector(32550, 16),
55703 => conv_std_logic_vector(32767, 16),
55704 => conv_std_logic_vector(32984, 16),
55705 => conv_std_logic_vector(33201, 16),
55706 => conv_std_logic_vector(33418, 16),
55707 => conv_std_logic_vector(33635, 16),
55708 => conv_std_logic_vector(33852, 16),
55709 => conv_std_logic_vector(34069, 16),
55710 => conv_std_logic_vector(34286, 16),
55711 => conv_std_logic_vector(34503, 16),
55712 => conv_std_logic_vector(34720, 16),
55713 => conv_std_logic_vector(34937, 16),
55714 => conv_std_logic_vector(35154, 16),
55715 => conv_std_logic_vector(35371, 16),
55716 => conv_std_logic_vector(35588, 16),
55717 => conv_std_logic_vector(35805, 16),
55718 => conv_std_logic_vector(36022, 16),
55719 => conv_std_logic_vector(36239, 16),
55720 => conv_std_logic_vector(36456, 16),
55721 => conv_std_logic_vector(36673, 16),
55722 => conv_std_logic_vector(36890, 16),
55723 => conv_std_logic_vector(37107, 16),
55724 => conv_std_logic_vector(37324, 16),
55725 => conv_std_logic_vector(37541, 16),
55726 => conv_std_logic_vector(37758, 16),
55727 => conv_std_logic_vector(37975, 16),
55728 => conv_std_logic_vector(38192, 16),
55729 => conv_std_logic_vector(38409, 16),
55730 => conv_std_logic_vector(38626, 16),
55731 => conv_std_logic_vector(38843, 16),
55732 => conv_std_logic_vector(39060, 16),
55733 => conv_std_logic_vector(39277, 16),
55734 => conv_std_logic_vector(39494, 16),
55735 => conv_std_logic_vector(39711, 16),
55736 => conv_std_logic_vector(39928, 16),
55737 => conv_std_logic_vector(40145, 16),
55738 => conv_std_logic_vector(40362, 16),
55739 => conv_std_logic_vector(40579, 16),
55740 => conv_std_logic_vector(40796, 16),
55741 => conv_std_logic_vector(41013, 16),
55742 => conv_std_logic_vector(41230, 16),
55743 => conv_std_logic_vector(41447, 16),
55744 => conv_std_logic_vector(41664, 16),
55745 => conv_std_logic_vector(41881, 16),
55746 => conv_std_logic_vector(42098, 16),
55747 => conv_std_logic_vector(42315, 16),
55748 => conv_std_logic_vector(42532, 16),
55749 => conv_std_logic_vector(42749, 16),
55750 => conv_std_logic_vector(42966, 16),
55751 => conv_std_logic_vector(43183, 16),
55752 => conv_std_logic_vector(43400, 16),
55753 => conv_std_logic_vector(43617, 16),
55754 => conv_std_logic_vector(43834, 16),
55755 => conv_std_logic_vector(44051, 16),
55756 => conv_std_logic_vector(44268, 16),
55757 => conv_std_logic_vector(44485, 16),
55758 => conv_std_logic_vector(44702, 16),
55759 => conv_std_logic_vector(44919, 16),
55760 => conv_std_logic_vector(45136, 16),
55761 => conv_std_logic_vector(45353, 16),
55762 => conv_std_logic_vector(45570, 16),
55763 => conv_std_logic_vector(45787, 16),
55764 => conv_std_logic_vector(46004, 16),
55765 => conv_std_logic_vector(46221, 16),
55766 => conv_std_logic_vector(46438, 16),
55767 => conv_std_logic_vector(46655, 16),
55768 => conv_std_logic_vector(46872, 16),
55769 => conv_std_logic_vector(47089, 16),
55770 => conv_std_logic_vector(47306, 16),
55771 => conv_std_logic_vector(47523, 16),
55772 => conv_std_logic_vector(47740, 16),
55773 => conv_std_logic_vector(47957, 16),
55774 => conv_std_logic_vector(48174, 16),
55775 => conv_std_logic_vector(48391, 16),
55776 => conv_std_logic_vector(48608, 16),
55777 => conv_std_logic_vector(48825, 16),
55778 => conv_std_logic_vector(49042, 16),
55779 => conv_std_logic_vector(49259, 16),
55780 => conv_std_logic_vector(49476, 16),
55781 => conv_std_logic_vector(49693, 16),
55782 => conv_std_logic_vector(49910, 16),
55783 => conv_std_logic_vector(50127, 16),
55784 => conv_std_logic_vector(50344, 16),
55785 => conv_std_logic_vector(50561, 16),
55786 => conv_std_logic_vector(50778, 16),
55787 => conv_std_logic_vector(50995, 16),
55788 => conv_std_logic_vector(51212, 16),
55789 => conv_std_logic_vector(51429, 16),
55790 => conv_std_logic_vector(51646, 16),
55791 => conv_std_logic_vector(51863, 16),
55792 => conv_std_logic_vector(52080, 16),
55793 => conv_std_logic_vector(52297, 16),
55794 => conv_std_logic_vector(52514, 16),
55795 => conv_std_logic_vector(52731, 16),
55796 => conv_std_logic_vector(52948, 16),
55797 => conv_std_logic_vector(53165, 16),
55798 => conv_std_logic_vector(53382, 16),
55799 => conv_std_logic_vector(53599, 16),
55800 => conv_std_logic_vector(53816, 16),
55801 => conv_std_logic_vector(54033, 16),
55802 => conv_std_logic_vector(54250, 16),
55803 => conv_std_logic_vector(54467, 16),
55804 => conv_std_logic_vector(54684, 16),
55805 => conv_std_logic_vector(54901, 16),
55806 => conv_std_logic_vector(55118, 16),
55807 => conv_std_logic_vector(55335, 16),
55808 => conv_std_logic_vector(0, 16),
55809 => conv_std_logic_vector(218, 16),
55810 => conv_std_logic_vector(436, 16),
55811 => conv_std_logic_vector(654, 16),
55812 => conv_std_logic_vector(872, 16),
55813 => conv_std_logic_vector(1090, 16),
55814 => conv_std_logic_vector(1308, 16),
55815 => conv_std_logic_vector(1526, 16),
55816 => conv_std_logic_vector(1744, 16),
55817 => conv_std_logic_vector(1962, 16),
55818 => conv_std_logic_vector(2180, 16),
55819 => conv_std_logic_vector(2398, 16),
55820 => conv_std_logic_vector(2616, 16),
55821 => conv_std_logic_vector(2834, 16),
55822 => conv_std_logic_vector(3052, 16),
55823 => conv_std_logic_vector(3270, 16),
55824 => conv_std_logic_vector(3488, 16),
55825 => conv_std_logic_vector(3706, 16),
55826 => conv_std_logic_vector(3924, 16),
55827 => conv_std_logic_vector(4142, 16),
55828 => conv_std_logic_vector(4360, 16),
55829 => conv_std_logic_vector(4578, 16),
55830 => conv_std_logic_vector(4796, 16),
55831 => conv_std_logic_vector(5014, 16),
55832 => conv_std_logic_vector(5232, 16),
55833 => conv_std_logic_vector(5450, 16),
55834 => conv_std_logic_vector(5668, 16),
55835 => conv_std_logic_vector(5886, 16),
55836 => conv_std_logic_vector(6104, 16),
55837 => conv_std_logic_vector(6322, 16),
55838 => conv_std_logic_vector(6540, 16),
55839 => conv_std_logic_vector(6758, 16),
55840 => conv_std_logic_vector(6976, 16),
55841 => conv_std_logic_vector(7194, 16),
55842 => conv_std_logic_vector(7412, 16),
55843 => conv_std_logic_vector(7630, 16),
55844 => conv_std_logic_vector(7848, 16),
55845 => conv_std_logic_vector(8066, 16),
55846 => conv_std_logic_vector(8284, 16),
55847 => conv_std_logic_vector(8502, 16),
55848 => conv_std_logic_vector(8720, 16),
55849 => conv_std_logic_vector(8938, 16),
55850 => conv_std_logic_vector(9156, 16),
55851 => conv_std_logic_vector(9374, 16),
55852 => conv_std_logic_vector(9592, 16),
55853 => conv_std_logic_vector(9810, 16),
55854 => conv_std_logic_vector(10028, 16),
55855 => conv_std_logic_vector(10246, 16),
55856 => conv_std_logic_vector(10464, 16),
55857 => conv_std_logic_vector(10682, 16),
55858 => conv_std_logic_vector(10900, 16),
55859 => conv_std_logic_vector(11118, 16),
55860 => conv_std_logic_vector(11336, 16),
55861 => conv_std_logic_vector(11554, 16),
55862 => conv_std_logic_vector(11772, 16),
55863 => conv_std_logic_vector(11990, 16),
55864 => conv_std_logic_vector(12208, 16),
55865 => conv_std_logic_vector(12426, 16),
55866 => conv_std_logic_vector(12644, 16),
55867 => conv_std_logic_vector(12862, 16),
55868 => conv_std_logic_vector(13080, 16),
55869 => conv_std_logic_vector(13298, 16),
55870 => conv_std_logic_vector(13516, 16),
55871 => conv_std_logic_vector(13734, 16),
55872 => conv_std_logic_vector(13952, 16),
55873 => conv_std_logic_vector(14170, 16),
55874 => conv_std_logic_vector(14388, 16),
55875 => conv_std_logic_vector(14606, 16),
55876 => conv_std_logic_vector(14824, 16),
55877 => conv_std_logic_vector(15042, 16),
55878 => conv_std_logic_vector(15260, 16),
55879 => conv_std_logic_vector(15478, 16),
55880 => conv_std_logic_vector(15696, 16),
55881 => conv_std_logic_vector(15914, 16),
55882 => conv_std_logic_vector(16132, 16),
55883 => conv_std_logic_vector(16350, 16),
55884 => conv_std_logic_vector(16568, 16),
55885 => conv_std_logic_vector(16786, 16),
55886 => conv_std_logic_vector(17004, 16),
55887 => conv_std_logic_vector(17222, 16),
55888 => conv_std_logic_vector(17440, 16),
55889 => conv_std_logic_vector(17658, 16),
55890 => conv_std_logic_vector(17876, 16),
55891 => conv_std_logic_vector(18094, 16),
55892 => conv_std_logic_vector(18312, 16),
55893 => conv_std_logic_vector(18530, 16),
55894 => conv_std_logic_vector(18748, 16),
55895 => conv_std_logic_vector(18966, 16),
55896 => conv_std_logic_vector(19184, 16),
55897 => conv_std_logic_vector(19402, 16),
55898 => conv_std_logic_vector(19620, 16),
55899 => conv_std_logic_vector(19838, 16),
55900 => conv_std_logic_vector(20056, 16),
55901 => conv_std_logic_vector(20274, 16),
55902 => conv_std_logic_vector(20492, 16),
55903 => conv_std_logic_vector(20710, 16),
55904 => conv_std_logic_vector(20928, 16),
55905 => conv_std_logic_vector(21146, 16),
55906 => conv_std_logic_vector(21364, 16),
55907 => conv_std_logic_vector(21582, 16),
55908 => conv_std_logic_vector(21800, 16),
55909 => conv_std_logic_vector(22018, 16),
55910 => conv_std_logic_vector(22236, 16),
55911 => conv_std_logic_vector(22454, 16),
55912 => conv_std_logic_vector(22672, 16),
55913 => conv_std_logic_vector(22890, 16),
55914 => conv_std_logic_vector(23108, 16),
55915 => conv_std_logic_vector(23326, 16),
55916 => conv_std_logic_vector(23544, 16),
55917 => conv_std_logic_vector(23762, 16),
55918 => conv_std_logic_vector(23980, 16),
55919 => conv_std_logic_vector(24198, 16),
55920 => conv_std_logic_vector(24416, 16),
55921 => conv_std_logic_vector(24634, 16),
55922 => conv_std_logic_vector(24852, 16),
55923 => conv_std_logic_vector(25070, 16),
55924 => conv_std_logic_vector(25288, 16),
55925 => conv_std_logic_vector(25506, 16),
55926 => conv_std_logic_vector(25724, 16),
55927 => conv_std_logic_vector(25942, 16),
55928 => conv_std_logic_vector(26160, 16),
55929 => conv_std_logic_vector(26378, 16),
55930 => conv_std_logic_vector(26596, 16),
55931 => conv_std_logic_vector(26814, 16),
55932 => conv_std_logic_vector(27032, 16),
55933 => conv_std_logic_vector(27250, 16),
55934 => conv_std_logic_vector(27468, 16),
55935 => conv_std_logic_vector(27686, 16),
55936 => conv_std_logic_vector(27904, 16),
55937 => conv_std_logic_vector(28122, 16),
55938 => conv_std_logic_vector(28340, 16),
55939 => conv_std_logic_vector(28558, 16),
55940 => conv_std_logic_vector(28776, 16),
55941 => conv_std_logic_vector(28994, 16),
55942 => conv_std_logic_vector(29212, 16),
55943 => conv_std_logic_vector(29430, 16),
55944 => conv_std_logic_vector(29648, 16),
55945 => conv_std_logic_vector(29866, 16),
55946 => conv_std_logic_vector(30084, 16),
55947 => conv_std_logic_vector(30302, 16),
55948 => conv_std_logic_vector(30520, 16),
55949 => conv_std_logic_vector(30738, 16),
55950 => conv_std_logic_vector(30956, 16),
55951 => conv_std_logic_vector(31174, 16),
55952 => conv_std_logic_vector(31392, 16),
55953 => conv_std_logic_vector(31610, 16),
55954 => conv_std_logic_vector(31828, 16),
55955 => conv_std_logic_vector(32046, 16),
55956 => conv_std_logic_vector(32264, 16),
55957 => conv_std_logic_vector(32482, 16),
55958 => conv_std_logic_vector(32700, 16),
55959 => conv_std_logic_vector(32918, 16),
55960 => conv_std_logic_vector(33136, 16),
55961 => conv_std_logic_vector(33354, 16),
55962 => conv_std_logic_vector(33572, 16),
55963 => conv_std_logic_vector(33790, 16),
55964 => conv_std_logic_vector(34008, 16),
55965 => conv_std_logic_vector(34226, 16),
55966 => conv_std_logic_vector(34444, 16),
55967 => conv_std_logic_vector(34662, 16),
55968 => conv_std_logic_vector(34880, 16),
55969 => conv_std_logic_vector(35098, 16),
55970 => conv_std_logic_vector(35316, 16),
55971 => conv_std_logic_vector(35534, 16),
55972 => conv_std_logic_vector(35752, 16),
55973 => conv_std_logic_vector(35970, 16),
55974 => conv_std_logic_vector(36188, 16),
55975 => conv_std_logic_vector(36406, 16),
55976 => conv_std_logic_vector(36624, 16),
55977 => conv_std_logic_vector(36842, 16),
55978 => conv_std_logic_vector(37060, 16),
55979 => conv_std_logic_vector(37278, 16),
55980 => conv_std_logic_vector(37496, 16),
55981 => conv_std_logic_vector(37714, 16),
55982 => conv_std_logic_vector(37932, 16),
55983 => conv_std_logic_vector(38150, 16),
55984 => conv_std_logic_vector(38368, 16),
55985 => conv_std_logic_vector(38586, 16),
55986 => conv_std_logic_vector(38804, 16),
55987 => conv_std_logic_vector(39022, 16),
55988 => conv_std_logic_vector(39240, 16),
55989 => conv_std_logic_vector(39458, 16),
55990 => conv_std_logic_vector(39676, 16),
55991 => conv_std_logic_vector(39894, 16),
55992 => conv_std_logic_vector(40112, 16),
55993 => conv_std_logic_vector(40330, 16),
55994 => conv_std_logic_vector(40548, 16),
55995 => conv_std_logic_vector(40766, 16),
55996 => conv_std_logic_vector(40984, 16),
55997 => conv_std_logic_vector(41202, 16),
55998 => conv_std_logic_vector(41420, 16),
55999 => conv_std_logic_vector(41638, 16),
56000 => conv_std_logic_vector(41856, 16),
56001 => conv_std_logic_vector(42074, 16),
56002 => conv_std_logic_vector(42292, 16),
56003 => conv_std_logic_vector(42510, 16),
56004 => conv_std_logic_vector(42728, 16),
56005 => conv_std_logic_vector(42946, 16),
56006 => conv_std_logic_vector(43164, 16),
56007 => conv_std_logic_vector(43382, 16),
56008 => conv_std_logic_vector(43600, 16),
56009 => conv_std_logic_vector(43818, 16),
56010 => conv_std_logic_vector(44036, 16),
56011 => conv_std_logic_vector(44254, 16),
56012 => conv_std_logic_vector(44472, 16),
56013 => conv_std_logic_vector(44690, 16),
56014 => conv_std_logic_vector(44908, 16),
56015 => conv_std_logic_vector(45126, 16),
56016 => conv_std_logic_vector(45344, 16),
56017 => conv_std_logic_vector(45562, 16),
56018 => conv_std_logic_vector(45780, 16),
56019 => conv_std_logic_vector(45998, 16),
56020 => conv_std_logic_vector(46216, 16),
56021 => conv_std_logic_vector(46434, 16),
56022 => conv_std_logic_vector(46652, 16),
56023 => conv_std_logic_vector(46870, 16),
56024 => conv_std_logic_vector(47088, 16),
56025 => conv_std_logic_vector(47306, 16),
56026 => conv_std_logic_vector(47524, 16),
56027 => conv_std_logic_vector(47742, 16),
56028 => conv_std_logic_vector(47960, 16),
56029 => conv_std_logic_vector(48178, 16),
56030 => conv_std_logic_vector(48396, 16),
56031 => conv_std_logic_vector(48614, 16),
56032 => conv_std_logic_vector(48832, 16),
56033 => conv_std_logic_vector(49050, 16),
56034 => conv_std_logic_vector(49268, 16),
56035 => conv_std_logic_vector(49486, 16),
56036 => conv_std_logic_vector(49704, 16),
56037 => conv_std_logic_vector(49922, 16),
56038 => conv_std_logic_vector(50140, 16),
56039 => conv_std_logic_vector(50358, 16),
56040 => conv_std_logic_vector(50576, 16),
56041 => conv_std_logic_vector(50794, 16),
56042 => conv_std_logic_vector(51012, 16),
56043 => conv_std_logic_vector(51230, 16),
56044 => conv_std_logic_vector(51448, 16),
56045 => conv_std_logic_vector(51666, 16),
56046 => conv_std_logic_vector(51884, 16),
56047 => conv_std_logic_vector(52102, 16),
56048 => conv_std_logic_vector(52320, 16),
56049 => conv_std_logic_vector(52538, 16),
56050 => conv_std_logic_vector(52756, 16),
56051 => conv_std_logic_vector(52974, 16),
56052 => conv_std_logic_vector(53192, 16),
56053 => conv_std_logic_vector(53410, 16),
56054 => conv_std_logic_vector(53628, 16),
56055 => conv_std_logic_vector(53846, 16),
56056 => conv_std_logic_vector(54064, 16),
56057 => conv_std_logic_vector(54282, 16),
56058 => conv_std_logic_vector(54500, 16),
56059 => conv_std_logic_vector(54718, 16),
56060 => conv_std_logic_vector(54936, 16),
56061 => conv_std_logic_vector(55154, 16),
56062 => conv_std_logic_vector(55372, 16),
56063 => conv_std_logic_vector(55590, 16),
56064 => conv_std_logic_vector(0, 16),
56065 => conv_std_logic_vector(219, 16),
56066 => conv_std_logic_vector(438, 16),
56067 => conv_std_logic_vector(657, 16),
56068 => conv_std_logic_vector(876, 16),
56069 => conv_std_logic_vector(1095, 16),
56070 => conv_std_logic_vector(1314, 16),
56071 => conv_std_logic_vector(1533, 16),
56072 => conv_std_logic_vector(1752, 16),
56073 => conv_std_logic_vector(1971, 16),
56074 => conv_std_logic_vector(2190, 16),
56075 => conv_std_logic_vector(2409, 16),
56076 => conv_std_logic_vector(2628, 16),
56077 => conv_std_logic_vector(2847, 16),
56078 => conv_std_logic_vector(3066, 16),
56079 => conv_std_logic_vector(3285, 16),
56080 => conv_std_logic_vector(3504, 16),
56081 => conv_std_logic_vector(3723, 16),
56082 => conv_std_logic_vector(3942, 16),
56083 => conv_std_logic_vector(4161, 16),
56084 => conv_std_logic_vector(4380, 16),
56085 => conv_std_logic_vector(4599, 16),
56086 => conv_std_logic_vector(4818, 16),
56087 => conv_std_logic_vector(5037, 16),
56088 => conv_std_logic_vector(5256, 16),
56089 => conv_std_logic_vector(5475, 16),
56090 => conv_std_logic_vector(5694, 16),
56091 => conv_std_logic_vector(5913, 16),
56092 => conv_std_logic_vector(6132, 16),
56093 => conv_std_logic_vector(6351, 16),
56094 => conv_std_logic_vector(6570, 16),
56095 => conv_std_logic_vector(6789, 16),
56096 => conv_std_logic_vector(7008, 16),
56097 => conv_std_logic_vector(7227, 16),
56098 => conv_std_logic_vector(7446, 16),
56099 => conv_std_logic_vector(7665, 16),
56100 => conv_std_logic_vector(7884, 16),
56101 => conv_std_logic_vector(8103, 16),
56102 => conv_std_logic_vector(8322, 16),
56103 => conv_std_logic_vector(8541, 16),
56104 => conv_std_logic_vector(8760, 16),
56105 => conv_std_logic_vector(8979, 16),
56106 => conv_std_logic_vector(9198, 16),
56107 => conv_std_logic_vector(9417, 16),
56108 => conv_std_logic_vector(9636, 16),
56109 => conv_std_logic_vector(9855, 16),
56110 => conv_std_logic_vector(10074, 16),
56111 => conv_std_logic_vector(10293, 16),
56112 => conv_std_logic_vector(10512, 16),
56113 => conv_std_logic_vector(10731, 16),
56114 => conv_std_logic_vector(10950, 16),
56115 => conv_std_logic_vector(11169, 16),
56116 => conv_std_logic_vector(11388, 16),
56117 => conv_std_logic_vector(11607, 16),
56118 => conv_std_logic_vector(11826, 16),
56119 => conv_std_logic_vector(12045, 16),
56120 => conv_std_logic_vector(12264, 16),
56121 => conv_std_logic_vector(12483, 16),
56122 => conv_std_logic_vector(12702, 16),
56123 => conv_std_logic_vector(12921, 16),
56124 => conv_std_logic_vector(13140, 16),
56125 => conv_std_logic_vector(13359, 16),
56126 => conv_std_logic_vector(13578, 16),
56127 => conv_std_logic_vector(13797, 16),
56128 => conv_std_logic_vector(14016, 16),
56129 => conv_std_logic_vector(14235, 16),
56130 => conv_std_logic_vector(14454, 16),
56131 => conv_std_logic_vector(14673, 16),
56132 => conv_std_logic_vector(14892, 16),
56133 => conv_std_logic_vector(15111, 16),
56134 => conv_std_logic_vector(15330, 16),
56135 => conv_std_logic_vector(15549, 16),
56136 => conv_std_logic_vector(15768, 16),
56137 => conv_std_logic_vector(15987, 16),
56138 => conv_std_logic_vector(16206, 16),
56139 => conv_std_logic_vector(16425, 16),
56140 => conv_std_logic_vector(16644, 16),
56141 => conv_std_logic_vector(16863, 16),
56142 => conv_std_logic_vector(17082, 16),
56143 => conv_std_logic_vector(17301, 16),
56144 => conv_std_logic_vector(17520, 16),
56145 => conv_std_logic_vector(17739, 16),
56146 => conv_std_logic_vector(17958, 16),
56147 => conv_std_logic_vector(18177, 16),
56148 => conv_std_logic_vector(18396, 16),
56149 => conv_std_logic_vector(18615, 16),
56150 => conv_std_logic_vector(18834, 16),
56151 => conv_std_logic_vector(19053, 16),
56152 => conv_std_logic_vector(19272, 16),
56153 => conv_std_logic_vector(19491, 16),
56154 => conv_std_logic_vector(19710, 16),
56155 => conv_std_logic_vector(19929, 16),
56156 => conv_std_logic_vector(20148, 16),
56157 => conv_std_logic_vector(20367, 16),
56158 => conv_std_logic_vector(20586, 16),
56159 => conv_std_logic_vector(20805, 16),
56160 => conv_std_logic_vector(21024, 16),
56161 => conv_std_logic_vector(21243, 16),
56162 => conv_std_logic_vector(21462, 16),
56163 => conv_std_logic_vector(21681, 16),
56164 => conv_std_logic_vector(21900, 16),
56165 => conv_std_logic_vector(22119, 16),
56166 => conv_std_logic_vector(22338, 16),
56167 => conv_std_logic_vector(22557, 16),
56168 => conv_std_logic_vector(22776, 16),
56169 => conv_std_logic_vector(22995, 16),
56170 => conv_std_logic_vector(23214, 16),
56171 => conv_std_logic_vector(23433, 16),
56172 => conv_std_logic_vector(23652, 16),
56173 => conv_std_logic_vector(23871, 16),
56174 => conv_std_logic_vector(24090, 16),
56175 => conv_std_logic_vector(24309, 16),
56176 => conv_std_logic_vector(24528, 16),
56177 => conv_std_logic_vector(24747, 16),
56178 => conv_std_logic_vector(24966, 16),
56179 => conv_std_logic_vector(25185, 16),
56180 => conv_std_logic_vector(25404, 16),
56181 => conv_std_logic_vector(25623, 16),
56182 => conv_std_logic_vector(25842, 16),
56183 => conv_std_logic_vector(26061, 16),
56184 => conv_std_logic_vector(26280, 16),
56185 => conv_std_logic_vector(26499, 16),
56186 => conv_std_logic_vector(26718, 16),
56187 => conv_std_logic_vector(26937, 16),
56188 => conv_std_logic_vector(27156, 16),
56189 => conv_std_logic_vector(27375, 16),
56190 => conv_std_logic_vector(27594, 16),
56191 => conv_std_logic_vector(27813, 16),
56192 => conv_std_logic_vector(28032, 16),
56193 => conv_std_logic_vector(28251, 16),
56194 => conv_std_logic_vector(28470, 16),
56195 => conv_std_logic_vector(28689, 16),
56196 => conv_std_logic_vector(28908, 16),
56197 => conv_std_logic_vector(29127, 16),
56198 => conv_std_logic_vector(29346, 16),
56199 => conv_std_logic_vector(29565, 16),
56200 => conv_std_logic_vector(29784, 16),
56201 => conv_std_logic_vector(30003, 16),
56202 => conv_std_logic_vector(30222, 16),
56203 => conv_std_logic_vector(30441, 16),
56204 => conv_std_logic_vector(30660, 16),
56205 => conv_std_logic_vector(30879, 16),
56206 => conv_std_logic_vector(31098, 16),
56207 => conv_std_logic_vector(31317, 16),
56208 => conv_std_logic_vector(31536, 16),
56209 => conv_std_logic_vector(31755, 16),
56210 => conv_std_logic_vector(31974, 16),
56211 => conv_std_logic_vector(32193, 16),
56212 => conv_std_logic_vector(32412, 16),
56213 => conv_std_logic_vector(32631, 16),
56214 => conv_std_logic_vector(32850, 16),
56215 => conv_std_logic_vector(33069, 16),
56216 => conv_std_logic_vector(33288, 16),
56217 => conv_std_logic_vector(33507, 16),
56218 => conv_std_logic_vector(33726, 16),
56219 => conv_std_logic_vector(33945, 16),
56220 => conv_std_logic_vector(34164, 16),
56221 => conv_std_logic_vector(34383, 16),
56222 => conv_std_logic_vector(34602, 16),
56223 => conv_std_logic_vector(34821, 16),
56224 => conv_std_logic_vector(35040, 16),
56225 => conv_std_logic_vector(35259, 16),
56226 => conv_std_logic_vector(35478, 16),
56227 => conv_std_logic_vector(35697, 16),
56228 => conv_std_logic_vector(35916, 16),
56229 => conv_std_logic_vector(36135, 16),
56230 => conv_std_logic_vector(36354, 16),
56231 => conv_std_logic_vector(36573, 16),
56232 => conv_std_logic_vector(36792, 16),
56233 => conv_std_logic_vector(37011, 16),
56234 => conv_std_logic_vector(37230, 16),
56235 => conv_std_logic_vector(37449, 16),
56236 => conv_std_logic_vector(37668, 16),
56237 => conv_std_logic_vector(37887, 16),
56238 => conv_std_logic_vector(38106, 16),
56239 => conv_std_logic_vector(38325, 16),
56240 => conv_std_logic_vector(38544, 16),
56241 => conv_std_logic_vector(38763, 16),
56242 => conv_std_logic_vector(38982, 16),
56243 => conv_std_logic_vector(39201, 16),
56244 => conv_std_logic_vector(39420, 16),
56245 => conv_std_logic_vector(39639, 16),
56246 => conv_std_logic_vector(39858, 16),
56247 => conv_std_logic_vector(40077, 16),
56248 => conv_std_logic_vector(40296, 16),
56249 => conv_std_logic_vector(40515, 16),
56250 => conv_std_logic_vector(40734, 16),
56251 => conv_std_logic_vector(40953, 16),
56252 => conv_std_logic_vector(41172, 16),
56253 => conv_std_logic_vector(41391, 16),
56254 => conv_std_logic_vector(41610, 16),
56255 => conv_std_logic_vector(41829, 16),
56256 => conv_std_logic_vector(42048, 16),
56257 => conv_std_logic_vector(42267, 16),
56258 => conv_std_logic_vector(42486, 16),
56259 => conv_std_logic_vector(42705, 16),
56260 => conv_std_logic_vector(42924, 16),
56261 => conv_std_logic_vector(43143, 16),
56262 => conv_std_logic_vector(43362, 16),
56263 => conv_std_logic_vector(43581, 16),
56264 => conv_std_logic_vector(43800, 16),
56265 => conv_std_logic_vector(44019, 16),
56266 => conv_std_logic_vector(44238, 16),
56267 => conv_std_logic_vector(44457, 16),
56268 => conv_std_logic_vector(44676, 16),
56269 => conv_std_logic_vector(44895, 16),
56270 => conv_std_logic_vector(45114, 16),
56271 => conv_std_logic_vector(45333, 16),
56272 => conv_std_logic_vector(45552, 16),
56273 => conv_std_logic_vector(45771, 16),
56274 => conv_std_logic_vector(45990, 16),
56275 => conv_std_logic_vector(46209, 16),
56276 => conv_std_logic_vector(46428, 16),
56277 => conv_std_logic_vector(46647, 16),
56278 => conv_std_logic_vector(46866, 16),
56279 => conv_std_logic_vector(47085, 16),
56280 => conv_std_logic_vector(47304, 16),
56281 => conv_std_logic_vector(47523, 16),
56282 => conv_std_logic_vector(47742, 16),
56283 => conv_std_logic_vector(47961, 16),
56284 => conv_std_logic_vector(48180, 16),
56285 => conv_std_logic_vector(48399, 16),
56286 => conv_std_logic_vector(48618, 16),
56287 => conv_std_logic_vector(48837, 16),
56288 => conv_std_logic_vector(49056, 16),
56289 => conv_std_logic_vector(49275, 16),
56290 => conv_std_logic_vector(49494, 16),
56291 => conv_std_logic_vector(49713, 16),
56292 => conv_std_logic_vector(49932, 16),
56293 => conv_std_logic_vector(50151, 16),
56294 => conv_std_logic_vector(50370, 16),
56295 => conv_std_logic_vector(50589, 16),
56296 => conv_std_logic_vector(50808, 16),
56297 => conv_std_logic_vector(51027, 16),
56298 => conv_std_logic_vector(51246, 16),
56299 => conv_std_logic_vector(51465, 16),
56300 => conv_std_logic_vector(51684, 16),
56301 => conv_std_logic_vector(51903, 16),
56302 => conv_std_logic_vector(52122, 16),
56303 => conv_std_logic_vector(52341, 16),
56304 => conv_std_logic_vector(52560, 16),
56305 => conv_std_logic_vector(52779, 16),
56306 => conv_std_logic_vector(52998, 16),
56307 => conv_std_logic_vector(53217, 16),
56308 => conv_std_logic_vector(53436, 16),
56309 => conv_std_logic_vector(53655, 16),
56310 => conv_std_logic_vector(53874, 16),
56311 => conv_std_logic_vector(54093, 16),
56312 => conv_std_logic_vector(54312, 16),
56313 => conv_std_logic_vector(54531, 16),
56314 => conv_std_logic_vector(54750, 16),
56315 => conv_std_logic_vector(54969, 16),
56316 => conv_std_logic_vector(55188, 16),
56317 => conv_std_logic_vector(55407, 16),
56318 => conv_std_logic_vector(55626, 16),
56319 => conv_std_logic_vector(55845, 16),
56320 => conv_std_logic_vector(0, 16),
56321 => conv_std_logic_vector(220, 16),
56322 => conv_std_logic_vector(440, 16),
56323 => conv_std_logic_vector(660, 16),
56324 => conv_std_logic_vector(880, 16),
56325 => conv_std_logic_vector(1100, 16),
56326 => conv_std_logic_vector(1320, 16),
56327 => conv_std_logic_vector(1540, 16),
56328 => conv_std_logic_vector(1760, 16),
56329 => conv_std_logic_vector(1980, 16),
56330 => conv_std_logic_vector(2200, 16),
56331 => conv_std_logic_vector(2420, 16),
56332 => conv_std_logic_vector(2640, 16),
56333 => conv_std_logic_vector(2860, 16),
56334 => conv_std_logic_vector(3080, 16),
56335 => conv_std_logic_vector(3300, 16),
56336 => conv_std_logic_vector(3520, 16),
56337 => conv_std_logic_vector(3740, 16),
56338 => conv_std_logic_vector(3960, 16),
56339 => conv_std_logic_vector(4180, 16),
56340 => conv_std_logic_vector(4400, 16),
56341 => conv_std_logic_vector(4620, 16),
56342 => conv_std_logic_vector(4840, 16),
56343 => conv_std_logic_vector(5060, 16),
56344 => conv_std_logic_vector(5280, 16),
56345 => conv_std_logic_vector(5500, 16),
56346 => conv_std_logic_vector(5720, 16),
56347 => conv_std_logic_vector(5940, 16),
56348 => conv_std_logic_vector(6160, 16),
56349 => conv_std_logic_vector(6380, 16),
56350 => conv_std_logic_vector(6600, 16),
56351 => conv_std_logic_vector(6820, 16),
56352 => conv_std_logic_vector(7040, 16),
56353 => conv_std_logic_vector(7260, 16),
56354 => conv_std_logic_vector(7480, 16),
56355 => conv_std_logic_vector(7700, 16),
56356 => conv_std_logic_vector(7920, 16),
56357 => conv_std_logic_vector(8140, 16),
56358 => conv_std_logic_vector(8360, 16),
56359 => conv_std_logic_vector(8580, 16),
56360 => conv_std_logic_vector(8800, 16),
56361 => conv_std_logic_vector(9020, 16),
56362 => conv_std_logic_vector(9240, 16),
56363 => conv_std_logic_vector(9460, 16),
56364 => conv_std_logic_vector(9680, 16),
56365 => conv_std_logic_vector(9900, 16),
56366 => conv_std_logic_vector(10120, 16),
56367 => conv_std_logic_vector(10340, 16),
56368 => conv_std_logic_vector(10560, 16),
56369 => conv_std_logic_vector(10780, 16),
56370 => conv_std_logic_vector(11000, 16),
56371 => conv_std_logic_vector(11220, 16),
56372 => conv_std_logic_vector(11440, 16),
56373 => conv_std_logic_vector(11660, 16),
56374 => conv_std_logic_vector(11880, 16),
56375 => conv_std_logic_vector(12100, 16),
56376 => conv_std_logic_vector(12320, 16),
56377 => conv_std_logic_vector(12540, 16),
56378 => conv_std_logic_vector(12760, 16),
56379 => conv_std_logic_vector(12980, 16),
56380 => conv_std_logic_vector(13200, 16),
56381 => conv_std_logic_vector(13420, 16),
56382 => conv_std_logic_vector(13640, 16),
56383 => conv_std_logic_vector(13860, 16),
56384 => conv_std_logic_vector(14080, 16),
56385 => conv_std_logic_vector(14300, 16),
56386 => conv_std_logic_vector(14520, 16),
56387 => conv_std_logic_vector(14740, 16),
56388 => conv_std_logic_vector(14960, 16),
56389 => conv_std_logic_vector(15180, 16),
56390 => conv_std_logic_vector(15400, 16),
56391 => conv_std_logic_vector(15620, 16),
56392 => conv_std_logic_vector(15840, 16),
56393 => conv_std_logic_vector(16060, 16),
56394 => conv_std_logic_vector(16280, 16),
56395 => conv_std_logic_vector(16500, 16),
56396 => conv_std_logic_vector(16720, 16),
56397 => conv_std_logic_vector(16940, 16),
56398 => conv_std_logic_vector(17160, 16),
56399 => conv_std_logic_vector(17380, 16),
56400 => conv_std_logic_vector(17600, 16),
56401 => conv_std_logic_vector(17820, 16),
56402 => conv_std_logic_vector(18040, 16),
56403 => conv_std_logic_vector(18260, 16),
56404 => conv_std_logic_vector(18480, 16),
56405 => conv_std_logic_vector(18700, 16),
56406 => conv_std_logic_vector(18920, 16),
56407 => conv_std_logic_vector(19140, 16),
56408 => conv_std_logic_vector(19360, 16),
56409 => conv_std_logic_vector(19580, 16),
56410 => conv_std_logic_vector(19800, 16),
56411 => conv_std_logic_vector(20020, 16),
56412 => conv_std_logic_vector(20240, 16),
56413 => conv_std_logic_vector(20460, 16),
56414 => conv_std_logic_vector(20680, 16),
56415 => conv_std_logic_vector(20900, 16),
56416 => conv_std_logic_vector(21120, 16),
56417 => conv_std_logic_vector(21340, 16),
56418 => conv_std_logic_vector(21560, 16),
56419 => conv_std_logic_vector(21780, 16),
56420 => conv_std_logic_vector(22000, 16),
56421 => conv_std_logic_vector(22220, 16),
56422 => conv_std_logic_vector(22440, 16),
56423 => conv_std_logic_vector(22660, 16),
56424 => conv_std_logic_vector(22880, 16),
56425 => conv_std_logic_vector(23100, 16),
56426 => conv_std_logic_vector(23320, 16),
56427 => conv_std_logic_vector(23540, 16),
56428 => conv_std_logic_vector(23760, 16),
56429 => conv_std_logic_vector(23980, 16),
56430 => conv_std_logic_vector(24200, 16),
56431 => conv_std_logic_vector(24420, 16),
56432 => conv_std_logic_vector(24640, 16),
56433 => conv_std_logic_vector(24860, 16),
56434 => conv_std_logic_vector(25080, 16),
56435 => conv_std_logic_vector(25300, 16),
56436 => conv_std_logic_vector(25520, 16),
56437 => conv_std_logic_vector(25740, 16),
56438 => conv_std_logic_vector(25960, 16),
56439 => conv_std_logic_vector(26180, 16),
56440 => conv_std_logic_vector(26400, 16),
56441 => conv_std_logic_vector(26620, 16),
56442 => conv_std_logic_vector(26840, 16),
56443 => conv_std_logic_vector(27060, 16),
56444 => conv_std_logic_vector(27280, 16),
56445 => conv_std_logic_vector(27500, 16),
56446 => conv_std_logic_vector(27720, 16),
56447 => conv_std_logic_vector(27940, 16),
56448 => conv_std_logic_vector(28160, 16),
56449 => conv_std_logic_vector(28380, 16),
56450 => conv_std_logic_vector(28600, 16),
56451 => conv_std_logic_vector(28820, 16),
56452 => conv_std_logic_vector(29040, 16),
56453 => conv_std_logic_vector(29260, 16),
56454 => conv_std_logic_vector(29480, 16),
56455 => conv_std_logic_vector(29700, 16),
56456 => conv_std_logic_vector(29920, 16),
56457 => conv_std_logic_vector(30140, 16),
56458 => conv_std_logic_vector(30360, 16),
56459 => conv_std_logic_vector(30580, 16),
56460 => conv_std_logic_vector(30800, 16),
56461 => conv_std_logic_vector(31020, 16),
56462 => conv_std_logic_vector(31240, 16),
56463 => conv_std_logic_vector(31460, 16),
56464 => conv_std_logic_vector(31680, 16),
56465 => conv_std_logic_vector(31900, 16),
56466 => conv_std_logic_vector(32120, 16),
56467 => conv_std_logic_vector(32340, 16),
56468 => conv_std_logic_vector(32560, 16),
56469 => conv_std_logic_vector(32780, 16),
56470 => conv_std_logic_vector(33000, 16),
56471 => conv_std_logic_vector(33220, 16),
56472 => conv_std_logic_vector(33440, 16),
56473 => conv_std_logic_vector(33660, 16),
56474 => conv_std_logic_vector(33880, 16),
56475 => conv_std_logic_vector(34100, 16),
56476 => conv_std_logic_vector(34320, 16),
56477 => conv_std_logic_vector(34540, 16),
56478 => conv_std_logic_vector(34760, 16),
56479 => conv_std_logic_vector(34980, 16),
56480 => conv_std_logic_vector(35200, 16),
56481 => conv_std_logic_vector(35420, 16),
56482 => conv_std_logic_vector(35640, 16),
56483 => conv_std_logic_vector(35860, 16),
56484 => conv_std_logic_vector(36080, 16),
56485 => conv_std_logic_vector(36300, 16),
56486 => conv_std_logic_vector(36520, 16),
56487 => conv_std_logic_vector(36740, 16),
56488 => conv_std_logic_vector(36960, 16),
56489 => conv_std_logic_vector(37180, 16),
56490 => conv_std_logic_vector(37400, 16),
56491 => conv_std_logic_vector(37620, 16),
56492 => conv_std_logic_vector(37840, 16),
56493 => conv_std_logic_vector(38060, 16),
56494 => conv_std_logic_vector(38280, 16),
56495 => conv_std_logic_vector(38500, 16),
56496 => conv_std_logic_vector(38720, 16),
56497 => conv_std_logic_vector(38940, 16),
56498 => conv_std_logic_vector(39160, 16),
56499 => conv_std_logic_vector(39380, 16),
56500 => conv_std_logic_vector(39600, 16),
56501 => conv_std_logic_vector(39820, 16),
56502 => conv_std_logic_vector(40040, 16),
56503 => conv_std_logic_vector(40260, 16),
56504 => conv_std_logic_vector(40480, 16),
56505 => conv_std_logic_vector(40700, 16),
56506 => conv_std_logic_vector(40920, 16),
56507 => conv_std_logic_vector(41140, 16),
56508 => conv_std_logic_vector(41360, 16),
56509 => conv_std_logic_vector(41580, 16),
56510 => conv_std_logic_vector(41800, 16),
56511 => conv_std_logic_vector(42020, 16),
56512 => conv_std_logic_vector(42240, 16),
56513 => conv_std_logic_vector(42460, 16),
56514 => conv_std_logic_vector(42680, 16),
56515 => conv_std_logic_vector(42900, 16),
56516 => conv_std_logic_vector(43120, 16),
56517 => conv_std_logic_vector(43340, 16),
56518 => conv_std_logic_vector(43560, 16),
56519 => conv_std_logic_vector(43780, 16),
56520 => conv_std_logic_vector(44000, 16),
56521 => conv_std_logic_vector(44220, 16),
56522 => conv_std_logic_vector(44440, 16),
56523 => conv_std_logic_vector(44660, 16),
56524 => conv_std_logic_vector(44880, 16),
56525 => conv_std_logic_vector(45100, 16),
56526 => conv_std_logic_vector(45320, 16),
56527 => conv_std_logic_vector(45540, 16),
56528 => conv_std_logic_vector(45760, 16),
56529 => conv_std_logic_vector(45980, 16),
56530 => conv_std_logic_vector(46200, 16),
56531 => conv_std_logic_vector(46420, 16),
56532 => conv_std_logic_vector(46640, 16),
56533 => conv_std_logic_vector(46860, 16),
56534 => conv_std_logic_vector(47080, 16),
56535 => conv_std_logic_vector(47300, 16),
56536 => conv_std_logic_vector(47520, 16),
56537 => conv_std_logic_vector(47740, 16),
56538 => conv_std_logic_vector(47960, 16),
56539 => conv_std_logic_vector(48180, 16),
56540 => conv_std_logic_vector(48400, 16),
56541 => conv_std_logic_vector(48620, 16),
56542 => conv_std_logic_vector(48840, 16),
56543 => conv_std_logic_vector(49060, 16),
56544 => conv_std_logic_vector(49280, 16),
56545 => conv_std_logic_vector(49500, 16),
56546 => conv_std_logic_vector(49720, 16),
56547 => conv_std_logic_vector(49940, 16),
56548 => conv_std_logic_vector(50160, 16),
56549 => conv_std_logic_vector(50380, 16),
56550 => conv_std_logic_vector(50600, 16),
56551 => conv_std_logic_vector(50820, 16),
56552 => conv_std_logic_vector(51040, 16),
56553 => conv_std_logic_vector(51260, 16),
56554 => conv_std_logic_vector(51480, 16),
56555 => conv_std_logic_vector(51700, 16),
56556 => conv_std_logic_vector(51920, 16),
56557 => conv_std_logic_vector(52140, 16),
56558 => conv_std_logic_vector(52360, 16),
56559 => conv_std_logic_vector(52580, 16),
56560 => conv_std_logic_vector(52800, 16),
56561 => conv_std_logic_vector(53020, 16),
56562 => conv_std_logic_vector(53240, 16),
56563 => conv_std_logic_vector(53460, 16),
56564 => conv_std_logic_vector(53680, 16),
56565 => conv_std_logic_vector(53900, 16),
56566 => conv_std_logic_vector(54120, 16),
56567 => conv_std_logic_vector(54340, 16),
56568 => conv_std_logic_vector(54560, 16),
56569 => conv_std_logic_vector(54780, 16),
56570 => conv_std_logic_vector(55000, 16),
56571 => conv_std_logic_vector(55220, 16),
56572 => conv_std_logic_vector(55440, 16),
56573 => conv_std_logic_vector(55660, 16),
56574 => conv_std_logic_vector(55880, 16),
56575 => conv_std_logic_vector(56100, 16),
56576 => conv_std_logic_vector(0, 16),
56577 => conv_std_logic_vector(221, 16),
56578 => conv_std_logic_vector(442, 16),
56579 => conv_std_logic_vector(663, 16),
56580 => conv_std_logic_vector(884, 16),
56581 => conv_std_logic_vector(1105, 16),
56582 => conv_std_logic_vector(1326, 16),
56583 => conv_std_logic_vector(1547, 16),
56584 => conv_std_logic_vector(1768, 16),
56585 => conv_std_logic_vector(1989, 16),
56586 => conv_std_logic_vector(2210, 16),
56587 => conv_std_logic_vector(2431, 16),
56588 => conv_std_logic_vector(2652, 16),
56589 => conv_std_logic_vector(2873, 16),
56590 => conv_std_logic_vector(3094, 16),
56591 => conv_std_logic_vector(3315, 16),
56592 => conv_std_logic_vector(3536, 16),
56593 => conv_std_logic_vector(3757, 16),
56594 => conv_std_logic_vector(3978, 16),
56595 => conv_std_logic_vector(4199, 16),
56596 => conv_std_logic_vector(4420, 16),
56597 => conv_std_logic_vector(4641, 16),
56598 => conv_std_logic_vector(4862, 16),
56599 => conv_std_logic_vector(5083, 16),
56600 => conv_std_logic_vector(5304, 16),
56601 => conv_std_logic_vector(5525, 16),
56602 => conv_std_logic_vector(5746, 16),
56603 => conv_std_logic_vector(5967, 16),
56604 => conv_std_logic_vector(6188, 16),
56605 => conv_std_logic_vector(6409, 16),
56606 => conv_std_logic_vector(6630, 16),
56607 => conv_std_logic_vector(6851, 16),
56608 => conv_std_logic_vector(7072, 16),
56609 => conv_std_logic_vector(7293, 16),
56610 => conv_std_logic_vector(7514, 16),
56611 => conv_std_logic_vector(7735, 16),
56612 => conv_std_logic_vector(7956, 16),
56613 => conv_std_logic_vector(8177, 16),
56614 => conv_std_logic_vector(8398, 16),
56615 => conv_std_logic_vector(8619, 16),
56616 => conv_std_logic_vector(8840, 16),
56617 => conv_std_logic_vector(9061, 16),
56618 => conv_std_logic_vector(9282, 16),
56619 => conv_std_logic_vector(9503, 16),
56620 => conv_std_logic_vector(9724, 16),
56621 => conv_std_logic_vector(9945, 16),
56622 => conv_std_logic_vector(10166, 16),
56623 => conv_std_logic_vector(10387, 16),
56624 => conv_std_logic_vector(10608, 16),
56625 => conv_std_logic_vector(10829, 16),
56626 => conv_std_logic_vector(11050, 16),
56627 => conv_std_logic_vector(11271, 16),
56628 => conv_std_logic_vector(11492, 16),
56629 => conv_std_logic_vector(11713, 16),
56630 => conv_std_logic_vector(11934, 16),
56631 => conv_std_logic_vector(12155, 16),
56632 => conv_std_logic_vector(12376, 16),
56633 => conv_std_logic_vector(12597, 16),
56634 => conv_std_logic_vector(12818, 16),
56635 => conv_std_logic_vector(13039, 16),
56636 => conv_std_logic_vector(13260, 16),
56637 => conv_std_logic_vector(13481, 16),
56638 => conv_std_logic_vector(13702, 16),
56639 => conv_std_logic_vector(13923, 16),
56640 => conv_std_logic_vector(14144, 16),
56641 => conv_std_logic_vector(14365, 16),
56642 => conv_std_logic_vector(14586, 16),
56643 => conv_std_logic_vector(14807, 16),
56644 => conv_std_logic_vector(15028, 16),
56645 => conv_std_logic_vector(15249, 16),
56646 => conv_std_logic_vector(15470, 16),
56647 => conv_std_logic_vector(15691, 16),
56648 => conv_std_logic_vector(15912, 16),
56649 => conv_std_logic_vector(16133, 16),
56650 => conv_std_logic_vector(16354, 16),
56651 => conv_std_logic_vector(16575, 16),
56652 => conv_std_logic_vector(16796, 16),
56653 => conv_std_logic_vector(17017, 16),
56654 => conv_std_logic_vector(17238, 16),
56655 => conv_std_logic_vector(17459, 16),
56656 => conv_std_logic_vector(17680, 16),
56657 => conv_std_logic_vector(17901, 16),
56658 => conv_std_logic_vector(18122, 16),
56659 => conv_std_logic_vector(18343, 16),
56660 => conv_std_logic_vector(18564, 16),
56661 => conv_std_logic_vector(18785, 16),
56662 => conv_std_logic_vector(19006, 16),
56663 => conv_std_logic_vector(19227, 16),
56664 => conv_std_logic_vector(19448, 16),
56665 => conv_std_logic_vector(19669, 16),
56666 => conv_std_logic_vector(19890, 16),
56667 => conv_std_logic_vector(20111, 16),
56668 => conv_std_logic_vector(20332, 16),
56669 => conv_std_logic_vector(20553, 16),
56670 => conv_std_logic_vector(20774, 16),
56671 => conv_std_logic_vector(20995, 16),
56672 => conv_std_logic_vector(21216, 16),
56673 => conv_std_logic_vector(21437, 16),
56674 => conv_std_logic_vector(21658, 16),
56675 => conv_std_logic_vector(21879, 16),
56676 => conv_std_logic_vector(22100, 16),
56677 => conv_std_logic_vector(22321, 16),
56678 => conv_std_logic_vector(22542, 16),
56679 => conv_std_logic_vector(22763, 16),
56680 => conv_std_logic_vector(22984, 16),
56681 => conv_std_logic_vector(23205, 16),
56682 => conv_std_logic_vector(23426, 16),
56683 => conv_std_logic_vector(23647, 16),
56684 => conv_std_logic_vector(23868, 16),
56685 => conv_std_logic_vector(24089, 16),
56686 => conv_std_logic_vector(24310, 16),
56687 => conv_std_logic_vector(24531, 16),
56688 => conv_std_logic_vector(24752, 16),
56689 => conv_std_logic_vector(24973, 16),
56690 => conv_std_logic_vector(25194, 16),
56691 => conv_std_logic_vector(25415, 16),
56692 => conv_std_logic_vector(25636, 16),
56693 => conv_std_logic_vector(25857, 16),
56694 => conv_std_logic_vector(26078, 16),
56695 => conv_std_logic_vector(26299, 16),
56696 => conv_std_logic_vector(26520, 16),
56697 => conv_std_logic_vector(26741, 16),
56698 => conv_std_logic_vector(26962, 16),
56699 => conv_std_logic_vector(27183, 16),
56700 => conv_std_logic_vector(27404, 16),
56701 => conv_std_logic_vector(27625, 16),
56702 => conv_std_logic_vector(27846, 16),
56703 => conv_std_logic_vector(28067, 16),
56704 => conv_std_logic_vector(28288, 16),
56705 => conv_std_logic_vector(28509, 16),
56706 => conv_std_logic_vector(28730, 16),
56707 => conv_std_logic_vector(28951, 16),
56708 => conv_std_logic_vector(29172, 16),
56709 => conv_std_logic_vector(29393, 16),
56710 => conv_std_logic_vector(29614, 16),
56711 => conv_std_logic_vector(29835, 16),
56712 => conv_std_logic_vector(30056, 16),
56713 => conv_std_logic_vector(30277, 16),
56714 => conv_std_logic_vector(30498, 16),
56715 => conv_std_logic_vector(30719, 16),
56716 => conv_std_logic_vector(30940, 16),
56717 => conv_std_logic_vector(31161, 16),
56718 => conv_std_logic_vector(31382, 16),
56719 => conv_std_logic_vector(31603, 16),
56720 => conv_std_logic_vector(31824, 16),
56721 => conv_std_logic_vector(32045, 16),
56722 => conv_std_logic_vector(32266, 16),
56723 => conv_std_logic_vector(32487, 16),
56724 => conv_std_logic_vector(32708, 16),
56725 => conv_std_logic_vector(32929, 16),
56726 => conv_std_logic_vector(33150, 16),
56727 => conv_std_logic_vector(33371, 16),
56728 => conv_std_logic_vector(33592, 16),
56729 => conv_std_logic_vector(33813, 16),
56730 => conv_std_logic_vector(34034, 16),
56731 => conv_std_logic_vector(34255, 16),
56732 => conv_std_logic_vector(34476, 16),
56733 => conv_std_logic_vector(34697, 16),
56734 => conv_std_logic_vector(34918, 16),
56735 => conv_std_logic_vector(35139, 16),
56736 => conv_std_logic_vector(35360, 16),
56737 => conv_std_logic_vector(35581, 16),
56738 => conv_std_logic_vector(35802, 16),
56739 => conv_std_logic_vector(36023, 16),
56740 => conv_std_logic_vector(36244, 16),
56741 => conv_std_logic_vector(36465, 16),
56742 => conv_std_logic_vector(36686, 16),
56743 => conv_std_logic_vector(36907, 16),
56744 => conv_std_logic_vector(37128, 16),
56745 => conv_std_logic_vector(37349, 16),
56746 => conv_std_logic_vector(37570, 16),
56747 => conv_std_logic_vector(37791, 16),
56748 => conv_std_logic_vector(38012, 16),
56749 => conv_std_logic_vector(38233, 16),
56750 => conv_std_logic_vector(38454, 16),
56751 => conv_std_logic_vector(38675, 16),
56752 => conv_std_logic_vector(38896, 16),
56753 => conv_std_logic_vector(39117, 16),
56754 => conv_std_logic_vector(39338, 16),
56755 => conv_std_logic_vector(39559, 16),
56756 => conv_std_logic_vector(39780, 16),
56757 => conv_std_logic_vector(40001, 16),
56758 => conv_std_logic_vector(40222, 16),
56759 => conv_std_logic_vector(40443, 16),
56760 => conv_std_logic_vector(40664, 16),
56761 => conv_std_logic_vector(40885, 16),
56762 => conv_std_logic_vector(41106, 16),
56763 => conv_std_logic_vector(41327, 16),
56764 => conv_std_logic_vector(41548, 16),
56765 => conv_std_logic_vector(41769, 16),
56766 => conv_std_logic_vector(41990, 16),
56767 => conv_std_logic_vector(42211, 16),
56768 => conv_std_logic_vector(42432, 16),
56769 => conv_std_logic_vector(42653, 16),
56770 => conv_std_logic_vector(42874, 16),
56771 => conv_std_logic_vector(43095, 16),
56772 => conv_std_logic_vector(43316, 16),
56773 => conv_std_logic_vector(43537, 16),
56774 => conv_std_logic_vector(43758, 16),
56775 => conv_std_logic_vector(43979, 16),
56776 => conv_std_logic_vector(44200, 16),
56777 => conv_std_logic_vector(44421, 16),
56778 => conv_std_logic_vector(44642, 16),
56779 => conv_std_logic_vector(44863, 16),
56780 => conv_std_logic_vector(45084, 16),
56781 => conv_std_logic_vector(45305, 16),
56782 => conv_std_logic_vector(45526, 16),
56783 => conv_std_logic_vector(45747, 16),
56784 => conv_std_logic_vector(45968, 16),
56785 => conv_std_logic_vector(46189, 16),
56786 => conv_std_logic_vector(46410, 16),
56787 => conv_std_logic_vector(46631, 16),
56788 => conv_std_logic_vector(46852, 16),
56789 => conv_std_logic_vector(47073, 16),
56790 => conv_std_logic_vector(47294, 16),
56791 => conv_std_logic_vector(47515, 16),
56792 => conv_std_logic_vector(47736, 16),
56793 => conv_std_logic_vector(47957, 16),
56794 => conv_std_logic_vector(48178, 16),
56795 => conv_std_logic_vector(48399, 16),
56796 => conv_std_logic_vector(48620, 16),
56797 => conv_std_logic_vector(48841, 16),
56798 => conv_std_logic_vector(49062, 16),
56799 => conv_std_logic_vector(49283, 16),
56800 => conv_std_logic_vector(49504, 16),
56801 => conv_std_logic_vector(49725, 16),
56802 => conv_std_logic_vector(49946, 16),
56803 => conv_std_logic_vector(50167, 16),
56804 => conv_std_logic_vector(50388, 16),
56805 => conv_std_logic_vector(50609, 16),
56806 => conv_std_logic_vector(50830, 16),
56807 => conv_std_logic_vector(51051, 16),
56808 => conv_std_logic_vector(51272, 16),
56809 => conv_std_logic_vector(51493, 16),
56810 => conv_std_logic_vector(51714, 16),
56811 => conv_std_logic_vector(51935, 16),
56812 => conv_std_logic_vector(52156, 16),
56813 => conv_std_logic_vector(52377, 16),
56814 => conv_std_logic_vector(52598, 16),
56815 => conv_std_logic_vector(52819, 16),
56816 => conv_std_logic_vector(53040, 16),
56817 => conv_std_logic_vector(53261, 16),
56818 => conv_std_logic_vector(53482, 16),
56819 => conv_std_logic_vector(53703, 16),
56820 => conv_std_logic_vector(53924, 16),
56821 => conv_std_logic_vector(54145, 16),
56822 => conv_std_logic_vector(54366, 16),
56823 => conv_std_logic_vector(54587, 16),
56824 => conv_std_logic_vector(54808, 16),
56825 => conv_std_logic_vector(55029, 16),
56826 => conv_std_logic_vector(55250, 16),
56827 => conv_std_logic_vector(55471, 16),
56828 => conv_std_logic_vector(55692, 16),
56829 => conv_std_logic_vector(55913, 16),
56830 => conv_std_logic_vector(56134, 16),
56831 => conv_std_logic_vector(56355, 16),
56832 => conv_std_logic_vector(0, 16),
56833 => conv_std_logic_vector(222, 16),
56834 => conv_std_logic_vector(444, 16),
56835 => conv_std_logic_vector(666, 16),
56836 => conv_std_logic_vector(888, 16),
56837 => conv_std_logic_vector(1110, 16),
56838 => conv_std_logic_vector(1332, 16),
56839 => conv_std_logic_vector(1554, 16),
56840 => conv_std_logic_vector(1776, 16),
56841 => conv_std_logic_vector(1998, 16),
56842 => conv_std_logic_vector(2220, 16),
56843 => conv_std_logic_vector(2442, 16),
56844 => conv_std_logic_vector(2664, 16),
56845 => conv_std_logic_vector(2886, 16),
56846 => conv_std_logic_vector(3108, 16),
56847 => conv_std_logic_vector(3330, 16),
56848 => conv_std_logic_vector(3552, 16),
56849 => conv_std_logic_vector(3774, 16),
56850 => conv_std_logic_vector(3996, 16),
56851 => conv_std_logic_vector(4218, 16),
56852 => conv_std_logic_vector(4440, 16),
56853 => conv_std_logic_vector(4662, 16),
56854 => conv_std_logic_vector(4884, 16),
56855 => conv_std_logic_vector(5106, 16),
56856 => conv_std_logic_vector(5328, 16),
56857 => conv_std_logic_vector(5550, 16),
56858 => conv_std_logic_vector(5772, 16),
56859 => conv_std_logic_vector(5994, 16),
56860 => conv_std_logic_vector(6216, 16),
56861 => conv_std_logic_vector(6438, 16),
56862 => conv_std_logic_vector(6660, 16),
56863 => conv_std_logic_vector(6882, 16),
56864 => conv_std_logic_vector(7104, 16),
56865 => conv_std_logic_vector(7326, 16),
56866 => conv_std_logic_vector(7548, 16),
56867 => conv_std_logic_vector(7770, 16),
56868 => conv_std_logic_vector(7992, 16),
56869 => conv_std_logic_vector(8214, 16),
56870 => conv_std_logic_vector(8436, 16),
56871 => conv_std_logic_vector(8658, 16),
56872 => conv_std_logic_vector(8880, 16),
56873 => conv_std_logic_vector(9102, 16),
56874 => conv_std_logic_vector(9324, 16),
56875 => conv_std_logic_vector(9546, 16),
56876 => conv_std_logic_vector(9768, 16),
56877 => conv_std_logic_vector(9990, 16),
56878 => conv_std_logic_vector(10212, 16),
56879 => conv_std_logic_vector(10434, 16),
56880 => conv_std_logic_vector(10656, 16),
56881 => conv_std_logic_vector(10878, 16),
56882 => conv_std_logic_vector(11100, 16),
56883 => conv_std_logic_vector(11322, 16),
56884 => conv_std_logic_vector(11544, 16),
56885 => conv_std_logic_vector(11766, 16),
56886 => conv_std_logic_vector(11988, 16),
56887 => conv_std_logic_vector(12210, 16),
56888 => conv_std_logic_vector(12432, 16),
56889 => conv_std_logic_vector(12654, 16),
56890 => conv_std_logic_vector(12876, 16),
56891 => conv_std_logic_vector(13098, 16),
56892 => conv_std_logic_vector(13320, 16),
56893 => conv_std_logic_vector(13542, 16),
56894 => conv_std_logic_vector(13764, 16),
56895 => conv_std_logic_vector(13986, 16),
56896 => conv_std_logic_vector(14208, 16),
56897 => conv_std_logic_vector(14430, 16),
56898 => conv_std_logic_vector(14652, 16),
56899 => conv_std_logic_vector(14874, 16),
56900 => conv_std_logic_vector(15096, 16),
56901 => conv_std_logic_vector(15318, 16),
56902 => conv_std_logic_vector(15540, 16),
56903 => conv_std_logic_vector(15762, 16),
56904 => conv_std_logic_vector(15984, 16),
56905 => conv_std_logic_vector(16206, 16),
56906 => conv_std_logic_vector(16428, 16),
56907 => conv_std_logic_vector(16650, 16),
56908 => conv_std_logic_vector(16872, 16),
56909 => conv_std_logic_vector(17094, 16),
56910 => conv_std_logic_vector(17316, 16),
56911 => conv_std_logic_vector(17538, 16),
56912 => conv_std_logic_vector(17760, 16),
56913 => conv_std_logic_vector(17982, 16),
56914 => conv_std_logic_vector(18204, 16),
56915 => conv_std_logic_vector(18426, 16),
56916 => conv_std_logic_vector(18648, 16),
56917 => conv_std_logic_vector(18870, 16),
56918 => conv_std_logic_vector(19092, 16),
56919 => conv_std_logic_vector(19314, 16),
56920 => conv_std_logic_vector(19536, 16),
56921 => conv_std_logic_vector(19758, 16),
56922 => conv_std_logic_vector(19980, 16),
56923 => conv_std_logic_vector(20202, 16),
56924 => conv_std_logic_vector(20424, 16),
56925 => conv_std_logic_vector(20646, 16),
56926 => conv_std_logic_vector(20868, 16),
56927 => conv_std_logic_vector(21090, 16),
56928 => conv_std_logic_vector(21312, 16),
56929 => conv_std_logic_vector(21534, 16),
56930 => conv_std_logic_vector(21756, 16),
56931 => conv_std_logic_vector(21978, 16),
56932 => conv_std_logic_vector(22200, 16),
56933 => conv_std_logic_vector(22422, 16),
56934 => conv_std_logic_vector(22644, 16),
56935 => conv_std_logic_vector(22866, 16),
56936 => conv_std_logic_vector(23088, 16),
56937 => conv_std_logic_vector(23310, 16),
56938 => conv_std_logic_vector(23532, 16),
56939 => conv_std_logic_vector(23754, 16),
56940 => conv_std_logic_vector(23976, 16),
56941 => conv_std_logic_vector(24198, 16),
56942 => conv_std_logic_vector(24420, 16),
56943 => conv_std_logic_vector(24642, 16),
56944 => conv_std_logic_vector(24864, 16),
56945 => conv_std_logic_vector(25086, 16),
56946 => conv_std_logic_vector(25308, 16),
56947 => conv_std_logic_vector(25530, 16),
56948 => conv_std_logic_vector(25752, 16),
56949 => conv_std_logic_vector(25974, 16),
56950 => conv_std_logic_vector(26196, 16),
56951 => conv_std_logic_vector(26418, 16),
56952 => conv_std_logic_vector(26640, 16),
56953 => conv_std_logic_vector(26862, 16),
56954 => conv_std_logic_vector(27084, 16),
56955 => conv_std_logic_vector(27306, 16),
56956 => conv_std_logic_vector(27528, 16),
56957 => conv_std_logic_vector(27750, 16),
56958 => conv_std_logic_vector(27972, 16),
56959 => conv_std_logic_vector(28194, 16),
56960 => conv_std_logic_vector(28416, 16),
56961 => conv_std_logic_vector(28638, 16),
56962 => conv_std_logic_vector(28860, 16),
56963 => conv_std_logic_vector(29082, 16),
56964 => conv_std_logic_vector(29304, 16),
56965 => conv_std_logic_vector(29526, 16),
56966 => conv_std_logic_vector(29748, 16),
56967 => conv_std_logic_vector(29970, 16),
56968 => conv_std_logic_vector(30192, 16),
56969 => conv_std_logic_vector(30414, 16),
56970 => conv_std_logic_vector(30636, 16),
56971 => conv_std_logic_vector(30858, 16),
56972 => conv_std_logic_vector(31080, 16),
56973 => conv_std_logic_vector(31302, 16),
56974 => conv_std_logic_vector(31524, 16),
56975 => conv_std_logic_vector(31746, 16),
56976 => conv_std_logic_vector(31968, 16),
56977 => conv_std_logic_vector(32190, 16),
56978 => conv_std_logic_vector(32412, 16),
56979 => conv_std_logic_vector(32634, 16),
56980 => conv_std_logic_vector(32856, 16),
56981 => conv_std_logic_vector(33078, 16),
56982 => conv_std_logic_vector(33300, 16),
56983 => conv_std_logic_vector(33522, 16),
56984 => conv_std_logic_vector(33744, 16),
56985 => conv_std_logic_vector(33966, 16),
56986 => conv_std_logic_vector(34188, 16),
56987 => conv_std_logic_vector(34410, 16),
56988 => conv_std_logic_vector(34632, 16),
56989 => conv_std_logic_vector(34854, 16),
56990 => conv_std_logic_vector(35076, 16),
56991 => conv_std_logic_vector(35298, 16),
56992 => conv_std_logic_vector(35520, 16),
56993 => conv_std_logic_vector(35742, 16),
56994 => conv_std_logic_vector(35964, 16),
56995 => conv_std_logic_vector(36186, 16),
56996 => conv_std_logic_vector(36408, 16),
56997 => conv_std_logic_vector(36630, 16),
56998 => conv_std_logic_vector(36852, 16),
56999 => conv_std_logic_vector(37074, 16),
57000 => conv_std_logic_vector(37296, 16),
57001 => conv_std_logic_vector(37518, 16),
57002 => conv_std_logic_vector(37740, 16),
57003 => conv_std_logic_vector(37962, 16),
57004 => conv_std_logic_vector(38184, 16),
57005 => conv_std_logic_vector(38406, 16),
57006 => conv_std_logic_vector(38628, 16),
57007 => conv_std_logic_vector(38850, 16),
57008 => conv_std_logic_vector(39072, 16),
57009 => conv_std_logic_vector(39294, 16),
57010 => conv_std_logic_vector(39516, 16),
57011 => conv_std_logic_vector(39738, 16),
57012 => conv_std_logic_vector(39960, 16),
57013 => conv_std_logic_vector(40182, 16),
57014 => conv_std_logic_vector(40404, 16),
57015 => conv_std_logic_vector(40626, 16),
57016 => conv_std_logic_vector(40848, 16),
57017 => conv_std_logic_vector(41070, 16),
57018 => conv_std_logic_vector(41292, 16),
57019 => conv_std_logic_vector(41514, 16),
57020 => conv_std_logic_vector(41736, 16),
57021 => conv_std_logic_vector(41958, 16),
57022 => conv_std_logic_vector(42180, 16),
57023 => conv_std_logic_vector(42402, 16),
57024 => conv_std_logic_vector(42624, 16),
57025 => conv_std_logic_vector(42846, 16),
57026 => conv_std_logic_vector(43068, 16),
57027 => conv_std_logic_vector(43290, 16),
57028 => conv_std_logic_vector(43512, 16),
57029 => conv_std_logic_vector(43734, 16),
57030 => conv_std_logic_vector(43956, 16),
57031 => conv_std_logic_vector(44178, 16),
57032 => conv_std_logic_vector(44400, 16),
57033 => conv_std_logic_vector(44622, 16),
57034 => conv_std_logic_vector(44844, 16),
57035 => conv_std_logic_vector(45066, 16),
57036 => conv_std_logic_vector(45288, 16),
57037 => conv_std_logic_vector(45510, 16),
57038 => conv_std_logic_vector(45732, 16),
57039 => conv_std_logic_vector(45954, 16),
57040 => conv_std_logic_vector(46176, 16),
57041 => conv_std_logic_vector(46398, 16),
57042 => conv_std_logic_vector(46620, 16),
57043 => conv_std_logic_vector(46842, 16),
57044 => conv_std_logic_vector(47064, 16),
57045 => conv_std_logic_vector(47286, 16),
57046 => conv_std_logic_vector(47508, 16),
57047 => conv_std_logic_vector(47730, 16),
57048 => conv_std_logic_vector(47952, 16),
57049 => conv_std_logic_vector(48174, 16),
57050 => conv_std_logic_vector(48396, 16),
57051 => conv_std_logic_vector(48618, 16),
57052 => conv_std_logic_vector(48840, 16),
57053 => conv_std_logic_vector(49062, 16),
57054 => conv_std_logic_vector(49284, 16),
57055 => conv_std_logic_vector(49506, 16),
57056 => conv_std_logic_vector(49728, 16),
57057 => conv_std_logic_vector(49950, 16),
57058 => conv_std_logic_vector(50172, 16),
57059 => conv_std_logic_vector(50394, 16),
57060 => conv_std_logic_vector(50616, 16),
57061 => conv_std_logic_vector(50838, 16),
57062 => conv_std_logic_vector(51060, 16),
57063 => conv_std_logic_vector(51282, 16),
57064 => conv_std_logic_vector(51504, 16),
57065 => conv_std_logic_vector(51726, 16),
57066 => conv_std_logic_vector(51948, 16),
57067 => conv_std_logic_vector(52170, 16),
57068 => conv_std_logic_vector(52392, 16),
57069 => conv_std_logic_vector(52614, 16),
57070 => conv_std_logic_vector(52836, 16),
57071 => conv_std_logic_vector(53058, 16),
57072 => conv_std_logic_vector(53280, 16),
57073 => conv_std_logic_vector(53502, 16),
57074 => conv_std_logic_vector(53724, 16),
57075 => conv_std_logic_vector(53946, 16),
57076 => conv_std_logic_vector(54168, 16),
57077 => conv_std_logic_vector(54390, 16),
57078 => conv_std_logic_vector(54612, 16),
57079 => conv_std_logic_vector(54834, 16),
57080 => conv_std_logic_vector(55056, 16),
57081 => conv_std_logic_vector(55278, 16),
57082 => conv_std_logic_vector(55500, 16),
57083 => conv_std_logic_vector(55722, 16),
57084 => conv_std_logic_vector(55944, 16),
57085 => conv_std_logic_vector(56166, 16),
57086 => conv_std_logic_vector(56388, 16),
57087 => conv_std_logic_vector(56610, 16),
57088 => conv_std_logic_vector(0, 16),
57089 => conv_std_logic_vector(223, 16),
57090 => conv_std_logic_vector(446, 16),
57091 => conv_std_logic_vector(669, 16),
57092 => conv_std_logic_vector(892, 16),
57093 => conv_std_logic_vector(1115, 16),
57094 => conv_std_logic_vector(1338, 16),
57095 => conv_std_logic_vector(1561, 16),
57096 => conv_std_logic_vector(1784, 16),
57097 => conv_std_logic_vector(2007, 16),
57098 => conv_std_logic_vector(2230, 16),
57099 => conv_std_logic_vector(2453, 16),
57100 => conv_std_logic_vector(2676, 16),
57101 => conv_std_logic_vector(2899, 16),
57102 => conv_std_logic_vector(3122, 16),
57103 => conv_std_logic_vector(3345, 16),
57104 => conv_std_logic_vector(3568, 16),
57105 => conv_std_logic_vector(3791, 16),
57106 => conv_std_logic_vector(4014, 16),
57107 => conv_std_logic_vector(4237, 16),
57108 => conv_std_logic_vector(4460, 16),
57109 => conv_std_logic_vector(4683, 16),
57110 => conv_std_logic_vector(4906, 16),
57111 => conv_std_logic_vector(5129, 16),
57112 => conv_std_logic_vector(5352, 16),
57113 => conv_std_logic_vector(5575, 16),
57114 => conv_std_logic_vector(5798, 16),
57115 => conv_std_logic_vector(6021, 16),
57116 => conv_std_logic_vector(6244, 16),
57117 => conv_std_logic_vector(6467, 16),
57118 => conv_std_logic_vector(6690, 16),
57119 => conv_std_logic_vector(6913, 16),
57120 => conv_std_logic_vector(7136, 16),
57121 => conv_std_logic_vector(7359, 16),
57122 => conv_std_logic_vector(7582, 16),
57123 => conv_std_logic_vector(7805, 16),
57124 => conv_std_logic_vector(8028, 16),
57125 => conv_std_logic_vector(8251, 16),
57126 => conv_std_logic_vector(8474, 16),
57127 => conv_std_logic_vector(8697, 16),
57128 => conv_std_logic_vector(8920, 16),
57129 => conv_std_logic_vector(9143, 16),
57130 => conv_std_logic_vector(9366, 16),
57131 => conv_std_logic_vector(9589, 16),
57132 => conv_std_logic_vector(9812, 16),
57133 => conv_std_logic_vector(10035, 16),
57134 => conv_std_logic_vector(10258, 16),
57135 => conv_std_logic_vector(10481, 16),
57136 => conv_std_logic_vector(10704, 16),
57137 => conv_std_logic_vector(10927, 16),
57138 => conv_std_logic_vector(11150, 16),
57139 => conv_std_logic_vector(11373, 16),
57140 => conv_std_logic_vector(11596, 16),
57141 => conv_std_logic_vector(11819, 16),
57142 => conv_std_logic_vector(12042, 16),
57143 => conv_std_logic_vector(12265, 16),
57144 => conv_std_logic_vector(12488, 16),
57145 => conv_std_logic_vector(12711, 16),
57146 => conv_std_logic_vector(12934, 16),
57147 => conv_std_logic_vector(13157, 16),
57148 => conv_std_logic_vector(13380, 16),
57149 => conv_std_logic_vector(13603, 16),
57150 => conv_std_logic_vector(13826, 16),
57151 => conv_std_logic_vector(14049, 16),
57152 => conv_std_logic_vector(14272, 16),
57153 => conv_std_logic_vector(14495, 16),
57154 => conv_std_logic_vector(14718, 16),
57155 => conv_std_logic_vector(14941, 16),
57156 => conv_std_logic_vector(15164, 16),
57157 => conv_std_logic_vector(15387, 16),
57158 => conv_std_logic_vector(15610, 16),
57159 => conv_std_logic_vector(15833, 16),
57160 => conv_std_logic_vector(16056, 16),
57161 => conv_std_logic_vector(16279, 16),
57162 => conv_std_logic_vector(16502, 16),
57163 => conv_std_logic_vector(16725, 16),
57164 => conv_std_logic_vector(16948, 16),
57165 => conv_std_logic_vector(17171, 16),
57166 => conv_std_logic_vector(17394, 16),
57167 => conv_std_logic_vector(17617, 16),
57168 => conv_std_logic_vector(17840, 16),
57169 => conv_std_logic_vector(18063, 16),
57170 => conv_std_logic_vector(18286, 16),
57171 => conv_std_logic_vector(18509, 16),
57172 => conv_std_logic_vector(18732, 16),
57173 => conv_std_logic_vector(18955, 16),
57174 => conv_std_logic_vector(19178, 16),
57175 => conv_std_logic_vector(19401, 16),
57176 => conv_std_logic_vector(19624, 16),
57177 => conv_std_logic_vector(19847, 16),
57178 => conv_std_logic_vector(20070, 16),
57179 => conv_std_logic_vector(20293, 16),
57180 => conv_std_logic_vector(20516, 16),
57181 => conv_std_logic_vector(20739, 16),
57182 => conv_std_logic_vector(20962, 16),
57183 => conv_std_logic_vector(21185, 16),
57184 => conv_std_logic_vector(21408, 16),
57185 => conv_std_logic_vector(21631, 16),
57186 => conv_std_logic_vector(21854, 16),
57187 => conv_std_logic_vector(22077, 16),
57188 => conv_std_logic_vector(22300, 16),
57189 => conv_std_logic_vector(22523, 16),
57190 => conv_std_logic_vector(22746, 16),
57191 => conv_std_logic_vector(22969, 16),
57192 => conv_std_logic_vector(23192, 16),
57193 => conv_std_logic_vector(23415, 16),
57194 => conv_std_logic_vector(23638, 16),
57195 => conv_std_logic_vector(23861, 16),
57196 => conv_std_logic_vector(24084, 16),
57197 => conv_std_logic_vector(24307, 16),
57198 => conv_std_logic_vector(24530, 16),
57199 => conv_std_logic_vector(24753, 16),
57200 => conv_std_logic_vector(24976, 16),
57201 => conv_std_logic_vector(25199, 16),
57202 => conv_std_logic_vector(25422, 16),
57203 => conv_std_logic_vector(25645, 16),
57204 => conv_std_logic_vector(25868, 16),
57205 => conv_std_logic_vector(26091, 16),
57206 => conv_std_logic_vector(26314, 16),
57207 => conv_std_logic_vector(26537, 16),
57208 => conv_std_logic_vector(26760, 16),
57209 => conv_std_logic_vector(26983, 16),
57210 => conv_std_logic_vector(27206, 16),
57211 => conv_std_logic_vector(27429, 16),
57212 => conv_std_logic_vector(27652, 16),
57213 => conv_std_logic_vector(27875, 16),
57214 => conv_std_logic_vector(28098, 16),
57215 => conv_std_logic_vector(28321, 16),
57216 => conv_std_logic_vector(28544, 16),
57217 => conv_std_logic_vector(28767, 16),
57218 => conv_std_logic_vector(28990, 16),
57219 => conv_std_logic_vector(29213, 16),
57220 => conv_std_logic_vector(29436, 16),
57221 => conv_std_logic_vector(29659, 16),
57222 => conv_std_logic_vector(29882, 16),
57223 => conv_std_logic_vector(30105, 16),
57224 => conv_std_logic_vector(30328, 16),
57225 => conv_std_logic_vector(30551, 16),
57226 => conv_std_logic_vector(30774, 16),
57227 => conv_std_logic_vector(30997, 16),
57228 => conv_std_logic_vector(31220, 16),
57229 => conv_std_logic_vector(31443, 16),
57230 => conv_std_logic_vector(31666, 16),
57231 => conv_std_logic_vector(31889, 16),
57232 => conv_std_logic_vector(32112, 16),
57233 => conv_std_logic_vector(32335, 16),
57234 => conv_std_logic_vector(32558, 16),
57235 => conv_std_logic_vector(32781, 16),
57236 => conv_std_logic_vector(33004, 16),
57237 => conv_std_logic_vector(33227, 16),
57238 => conv_std_logic_vector(33450, 16),
57239 => conv_std_logic_vector(33673, 16),
57240 => conv_std_logic_vector(33896, 16),
57241 => conv_std_logic_vector(34119, 16),
57242 => conv_std_logic_vector(34342, 16),
57243 => conv_std_logic_vector(34565, 16),
57244 => conv_std_logic_vector(34788, 16),
57245 => conv_std_logic_vector(35011, 16),
57246 => conv_std_logic_vector(35234, 16),
57247 => conv_std_logic_vector(35457, 16),
57248 => conv_std_logic_vector(35680, 16),
57249 => conv_std_logic_vector(35903, 16),
57250 => conv_std_logic_vector(36126, 16),
57251 => conv_std_logic_vector(36349, 16),
57252 => conv_std_logic_vector(36572, 16),
57253 => conv_std_logic_vector(36795, 16),
57254 => conv_std_logic_vector(37018, 16),
57255 => conv_std_logic_vector(37241, 16),
57256 => conv_std_logic_vector(37464, 16),
57257 => conv_std_logic_vector(37687, 16),
57258 => conv_std_logic_vector(37910, 16),
57259 => conv_std_logic_vector(38133, 16),
57260 => conv_std_logic_vector(38356, 16),
57261 => conv_std_logic_vector(38579, 16),
57262 => conv_std_logic_vector(38802, 16),
57263 => conv_std_logic_vector(39025, 16),
57264 => conv_std_logic_vector(39248, 16),
57265 => conv_std_logic_vector(39471, 16),
57266 => conv_std_logic_vector(39694, 16),
57267 => conv_std_logic_vector(39917, 16),
57268 => conv_std_logic_vector(40140, 16),
57269 => conv_std_logic_vector(40363, 16),
57270 => conv_std_logic_vector(40586, 16),
57271 => conv_std_logic_vector(40809, 16),
57272 => conv_std_logic_vector(41032, 16),
57273 => conv_std_logic_vector(41255, 16),
57274 => conv_std_logic_vector(41478, 16),
57275 => conv_std_logic_vector(41701, 16),
57276 => conv_std_logic_vector(41924, 16),
57277 => conv_std_logic_vector(42147, 16),
57278 => conv_std_logic_vector(42370, 16),
57279 => conv_std_logic_vector(42593, 16),
57280 => conv_std_logic_vector(42816, 16),
57281 => conv_std_logic_vector(43039, 16),
57282 => conv_std_logic_vector(43262, 16),
57283 => conv_std_logic_vector(43485, 16),
57284 => conv_std_logic_vector(43708, 16),
57285 => conv_std_logic_vector(43931, 16),
57286 => conv_std_logic_vector(44154, 16),
57287 => conv_std_logic_vector(44377, 16),
57288 => conv_std_logic_vector(44600, 16),
57289 => conv_std_logic_vector(44823, 16),
57290 => conv_std_logic_vector(45046, 16),
57291 => conv_std_logic_vector(45269, 16),
57292 => conv_std_logic_vector(45492, 16),
57293 => conv_std_logic_vector(45715, 16),
57294 => conv_std_logic_vector(45938, 16),
57295 => conv_std_logic_vector(46161, 16),
57296 => conv_std_logic_vector(46384, 16),
57297 => conv_std_logic_vector(46607, 16),
57298 => conv_std_logic_vector(46830, 16),
57299 => conv_std_logic_vector(47053, 16),
57300 => conv_std_logic_vector(47276, 16),
57301 => conv_std_logic_vector(47499, 16),
57302 => conv_std_logic_vector(47722, 16),
57303 => conv_std_logic_vector(47945, 16),
57304 => conv_std_logic_vector(48168, 16),
57305 => conv_std_logic_vector(48391, 16),
57306 => conv_std_logic_vector(48614, 16),
57307 => conv_std_logic_vector(48837, 16),
57308 => conv_std_logic_vector(49060, 16),
57309 => conv_std_logic_vector(49283, 16),
57310 => conv_std_logic_vector(49506, 16),
57311 => conv_std_logic_vector(49729, 16),
57312 => conv_std_logic_vector(49952, 16),
57313 => conv_std_logic_vector(50175, 16),
57314 => conv_std_logic_vector(50398, 16),
57315 => conv_std_logic_vector(50621, 16),
57316 => conv_std_logic_vector(50844, 16),
57317 => conv_std_logic_vector(51067, 16),
57318 => conv_std_logic_vector(51290, 16),
57319 => conv_std_logic_vector(51513, 16),
57320 => conv_std_logic_vector(51736, 16),
57321 => conv_std_logic_vector(51959, 16),
57322 => conv_std_logic_vector(52182, 16),
57323 => conv_std_logic_vector(52405, 16),
57324 => conv_std_logic_vector(52628, 16),
57325 => conv_std_logic_vector(52851, 16),
57326 => conv_std_logic_vector(53074, 16),
57327 => conv_std_logic_vector(53297, 16),
57328 => conv_std_logic_vector(53520, 16),
57329 => conv_std_logic_vector(53743, 16),
57330 => conv_std_logic_vector(53966, 16),
57331 => conv_std_logic_vector(54189, 16),
57332 => conv_std_logic_vector(54412, 16),
57333 => conv_std_logic_vector(54635, 16),
57334 => conv_std_logic_vector(54858, 16),
57335 => conv_std_logic_vector(55081, 16),
57336 => conv_std_logic_vector(55304, 16),
57337 => conv_std_logic_vector(55527, 16),
57338 => conv_std_logic_vector(55750, 16),
57339 => conv_std_logic_vector(55973, 16),
57340 => conv_std_logic_vector(56196, 16),
57341 => conv_std_logic_vector(56419, 16),
57342 => conv_std_logic_vector(56642, 16),
57343 => conv_std_logic_vector(56865, 16),
57344 => conv_std_logic_vector(0, 16),
57345 => conv_std_logic_vector(224, 16),
57346 => conv_std_logic_vector(448, 16),
57347 => conv_std_logic_vector(672, 16),
57348 => conv_std_logic_vector(896, 16),
57349 => conv_std_logic_vector(1120, 16),
57350 => conv_std_logic_vector(1344, 16),
57351 => conv_std_logic_vector(1568, 16),
57352 => conv_std_logic_vector(1792, 16),
57353 => conv_std_logic_vector(2016, 16),
57354 => conv_std_logic_vector(2240, 16),
57355 => conv_std_logic_vector(2464, 16),
57356 => conv_std_logic_vector(2688, 16),
57357 => conv_std_logic_vector(2912, 16),
57358 => conv_std_logic_vector(3136, 16),
57359 => conv_std_logic_vector(3360, 16),
57360 => conv_std_logic_vector(3584, 16),
57361 => conv_std_logic_vector(3808, 16),
57362 => conv_std_logic_vector(4032, 16),
57363 => conv_std_logic_vector(4256, 16),
57364 => conv_std_logic_vector(4480, 16),
57365 => conv_std_logic_vector(4704, 16),
57366 => conv_std_logic_vector(4928, 16),
57367 => conv_std_logic_vector(5152, 16),
57368 => conv_std_logic_vector(5376, 16),
57369 => conv_std_logic_vector(5600, 16),
57370 => conv_std_logic_vector(5824, 16),
57371 => conv_std_logic_vector(6048, 16),
57372 => conv_std_logic_vector(6272, 16),
57373 => conv_std_logic_vector(6496, 16),
57374 => conv_std_logic_vector(6720, 16),
57375 => conv_std_logic_vector(6944, 16),
57376 => conv_std_logic_vector(7168, 16),
57377 => conv_std_logic_vector(7392, 16),
57378 => conv_std_logic_vector(7616, 16),
57379 => conv_std_logic_vector(7840, 16),
57380 => conv_std_logic_vector(8064, 16),
57381 => conv_std_logic_vector(8288, 16),
57382 => conv_std_logic_vector(8512, 16),
57383 => conv_std_logic_vector(8736, 16),
57384 => conv_std_logic_vector(8960, 16),
57385 => conv_std_logic_vector(9184, 16),
57386 => conv_std_logic_vector(9408, 16),
57387 => conv_std_logic_vector(9632, 16),
57388 => conv_std_logic_vector(9856, 16),
57389 => conv_std_logic_vector(10080, 16),
57390 => conv_std_logic_vector(10304, 16),
57391 => conv_std_logic_vector(10528, 16),
57392 => conv_std_logic_vector(10752, 16),
57393 => conv_std_logic_vector(10976, 16),
57394 => conv_std_logic_vector(11200, 16),
57395 => conv_std_logic_vector(11424, 16),
57396 => conv_std_logic_vector(11648, 16),
57397 => conv_std_logic_vector(11872, 16),
57398 => conv_std_logic_vector(12096, 16),
57399 => conv_std_logic_vector(12320, 16),
57400 => conv_std_logic_vector(12544, 16),
57401 => conv_std_logic_vector(12768, 16),
57402 => conv_std_logic_vector(12992, 16),
57403 => conv_std_logic_vector(13216, 16),
57404 => conv_std_logic_vector(13440, 16),
57405 => conv_std_logic_vector(13664, 16),
57406 => conv_std_logic_vector(13888, 16),
57407 => conv_std_logic_vector(14112, 16),
57408 => conv_std_logic_vector(14336, 16),
57409 => conv_std_logic_vector(14560, 16),
57410 => conv_std_logic_vector(14784, 16),
57411 => conv_std_logic_vector(15008, 16),
57412 => conv_std_logic_vector(15232, 16),
57413 => conv_std_logic_vector(15456, 16),
57414 => conv_std_logic_vector(15680, 16),
57415 => conv_std_logic_vector(15904, 16),
57416 => conv_std_logic_vector(16128, 16),
57417 => conv_std_logic_vector(16352, 16),
57418 => conv_std_logic_vector(16576, 16),
57419 => conv_std_logic_vector(16800, 16),
57420 => conv_std_logic_vector(17024, 16),
57421 => conv_std_logic_vector(17248, 16),
57422 => conv_std_logic_vector(17472, 16),
57423 => conv_std_logic_vector(17696, 16),
57424 => conv_std_logic_vector(17920, 16),
57425 => conv_std_logic_vector(18144, 16),
57426 => conv_std_logic_vector(18368, 16),
57427 => conv_std_logic_vector(18592, 16),
57428 => conv_std_logic_vector(18816, 16),
57429 => conv_std_logic_vector(19040, 16),
57430 => conv_std_logic_vector(19264, 16),
57431 => conv_std_logic_vector(19488, 16),
57432 => conv_std_logic_vector(19712, 16),
57433 => conv_std_logic_vector(19936, 16),
57434 => conv_std_logic_vector(20160, 16),
57435 => conv_std_logic_vector(20384, 16),
57436 => conv_std_logic_vector(20608, 16),
57437 => conv_std_logic_vector(20832, 16),
57438 => conv_std_logic_vector(21056, 16),
57439 => conv_std_logic_vector(21280, 16),
57440 => conv_std_logic_vector(21504, 16),
57441 => conv_std_logic_vector(21728, 16),
57442 => conv_std_logic_vector(21952, 16),
57443 => conv_std_logic_vector(22176, 16),
57444 => conv_std_logic_vector(22400, 16),
57445 => conv_std_logic_vector(22624, 16),
57446 => conv_std_logic_vector(22848, 16),
57447 => conv_std_logic_vector(23072, 16),
57448 => conv_std_logic_vector(23296, 16),
57449 => conv_std_logic_vector(23520, 16),
57450 => conv_std_logic_vector(23744, 16),
57451 => conv_std_logic_vector(23968, 16),
57452 => conv_std_logic_vector(24192, 16),
57453 => conv_std_logic_vector(24416, 16),
57454 => conv_std_logic_vector(24640, 16),
57455 => conv_std_logic_vector(24864, 16),
57456 => conv_std_logic_vector(25088, 16),
57457 => conv_std_logic_vector(25312, 16),
57458 => conv_std_logic_vector(25536, 16),
57459 => conv_std_logic_vector(25760, 16),
57460 => conv_std_logic_vector(25984, 16),
57461 => conv_std_logic_vector(26208, 16),
57462 => conv_std_logic_vector(26432, 16),
57463 => conv_std_logic_vector(26656, 16),
57464 => conv_std_logic_vector(26880, 16),
57465 => conv_std_logic_vector(27104, 16),
57466 => conv_std_logic_vector(27328, 16),
57467 => conv_std_logic_vector(27552, 16),
57468 => conv_std_logic_vector(27776, 16),
57469 => conv_std_logic_vector(28000, 16),
57470 => conv_std_logic_vector(28224, 16),
57471 => conv_std_logic_vector(28448, 16),
57472 => conv_std_logic_vector(28672, 16),
57473 => conv_std_logic_vector(28896, 16),
57474 => conv_std_logic_vector(29120, 16),
57475 => conv_std_logic_vector(29344, 16),
57476 => conv_std_logic_vector(29568, 16),
57477 => conv_std_logic_vector(29792, 16),
57478 => conv_std_logic_vector(30016, 16),
57479 => conv_std_logic_vector(30240, 16),
57480 => conv_std_logic_vector(30464, 16),
57481 => conv_std_logic_vector(30688, 16),
57482 => conv_std_logic_vector(30912, 16),
57483 => conv_std_logic_vector(31136, 16),
57484 => conv_std_logic_vector(31360, 16),
57485 => conv_std_logic_vector(31584, 16),
57486 => conv_std_logic_vector(31808, 16),
57487 => conv_std_logic_vector(32032, 16),
57488 => conv_std_logic_vector(32256, 16),
57489 => conv_std_logic_vector(32480, 16),
57490 => conv_std_logic_vector(32704, 16),
57491 => conv_std_logic_vector(32928, 16),
57492 => conv_std_logic_vector(33152, 16),
57493 => conv_std_logic_vector(33376, 16),
57494 => conv_std_logic_vector(33600, 16),
57495 => conv_std_logic_vector(33824, 16),
57496 => conv_std_logic_vector(34048, 16),
57497 => conv_std_logic_vector(34272, 16),
57498 => conv_std_logic_vector(34496, 16),
57499 => conv_std_logic_vector(34720, 16),
57500 => conv_std_logic_vector(34944, 16),
57501 => conv_std_logic_vector(35168, 16),
57502 => conv_std_logic_vector(35392, 16),
57503 => conv_std_logic_vector(35616, 16),
57504 => conv_std_logic_vector(35840, 16),
57505 => conv_std_logic_vector(36064, 16),
57506 => conv_std_logic_vector(36288, 16),
57507 => conv_std_logic_vector(36512, 16),
57508 => conv_std_logic_vector(36736, 16),
57509 => conv_std_logic_vector(36960, 16),
57510 => conv_std_logic_vector(37184, 16),
57511 => conv_std_logic_vector(37408, 16),
57512 => conv_std_logic_vector(37632, 16),
57513 => conv_std_logic_vector(37856, 16),
57514 => conv_std_logic_vector(38080, 16),
57515 => conv_std_logic_vector(38304, 16),
57516 => conv_std_logic_vector(38528, 16),
57517 => conv_std_logic_vector(38752, 16),
57518 => conv_std_logic_vector(38976, 16),
57519 => conv_std_logic_vector(39200, 16),
57520 => conv_std_logic_vector(39424, 16),
57521 => conv_std_logic_vector(39648, 16),
57522 => conv_std_logic_vector(39872, 16),
57523 => conv_std_logic_vector(40096, 16),
57524 => conv_std_logic_vector(40320, 16),
57525 => conv_std_logic_vector(40544, 16),
57526 => conv_std_logic_vector(40768, 16),
57527 => conv_std_logic_vector(40992, 16),
57528 => conv_std_logic_vector(41216, 16),
57529 => conv_std_logic_vector(41440, 16),
57530 => conv_std_logic_vector(41664, 16),
57531 => conv_std_logic_vector(41888, 16),
57532 => conv_std_logic_vector(42112, 16),
57533 => conv_std_logic_vector(42336, 16),
57534 => conv_std_logic_vector(42560, 16),
57535 => conv_std_logic_vector(42784, 16),
57536 => conv_std_logic_vector(43008, 16),
57537 => conv_std_logic_vector(43232, 16),
57538 => conv_std_logic_vector(43456, 16),
57539 => conv_std_logic_vector(43680, 16),
57540 => conv_std_logic_vector(43904, 16),
57541 => conv_std_logic_vector(44128, 16),
57542 => conv_std_logic_vector(44352, 16),
57543 => conv_std_logic_vector(44576, 16),
57544 => conv_std_logic_vector(44800, 16),
57545 => conv_std_logic_vector(45024, 16),
57546 => conv_std_logic_vector(45248, 16),
57547 => conv_std_logic_vector(45472, 16),
57548 => conv_std_logic_vector(45696, 16),
57549 => conv_std_logic_vector(45920, 16),
57550 => conv_std_logic_vector(46144, 16),
57551 => conv_std_logic_vector(46368, 16),
57552 => conv_std_logic_vector(46592, 16),
57553 => conv_std_logic_vector(46816, 16),
57554 => conv_std_logic_vector(47040, 16),
57555 => conv_std_logic_vector(47264, 16),
57556 => conv_std_logic_vector(47488, 16),
57557 => conv_std_logic_vector(47712, 16),
57558 => conv_std_logic_vector(47936, 16),
57559 => conv_std_logic_vector(48160, 16),
57560 => conv_std_logic_vector(48384, 16),
57561 => conv_std_logic_vector(48608, 16),
57562 => conv_std_logic_vector(48832, 16),
57563 => conv_std_logic_vector(49056, 16),
57564 => conv_std_logic_vector(49280, 16),
57565 => conv_std_logic_vector(49504, 16),
57566 => conv_std_logic_vector(49728, 16),
57567 => conv_std_logic_vector(49952, 16),
57568 => conv_std_logic_vector(50176, 16),
57569 => conv_std_logic_vector(50400, 16),
57570 => conv_std_logic_vector(50624, 16),
57571 => conv_std_logic_vector(50848, 16),
57572 => conv_std_logic_vector(51072, 16),
57573 => conv_std_logic_vector(51296, 16),
57574 => conv_std_logic_vector(51520, 16),
57575 => conv_std_logic_vector(51744, 16),
57576 => conv_std_logic_vector(51968, 16),
57577 => conv_std_logic_vector(52192, 16),
57578 => conv_std_logic_vector(52416, 16),
57579 => conv_std_logic_vector(52640, 16),
57580 => conv_std_logic_vector(52864, 16),
57581 => conv_std_logic_vector(53088, 16),
57582 => conv_std_logic_vector(53312, 16),
57583 => conv_std_logic_vector(53536, 16),
57584 => conv_std_logic_vector(53760, 16),
57585 => conv_std_logic_vector(53984, 16),
57586 => conv_std_logic_vector(54208, 16),
57587 => conv_std_logic_vector(54432, 16),
57588 => conv_std_logic_vector(54656, 16),
57589 => conv_std_logic_vector(54880, 16),
57590 => conv_std_logic_vector(55104, 16),
57591 => conv_std_logic_vector(55328, 16),
57592 => conv_std_logic_vector(55552, 16),
57593 => conv_std_logic_vector(55776, 16),
57594 => conv_std_logic_vector(56000, 16),
57595 => conv_std_logic_vector(56224, 16),
57596 => conv_std_logic_vector(56448, 16),
57597 => conv_std_logic_vector(56672, 16),
57598 => conv_std_logic_vector(56896, 16),
57599 => conv_std_logic_vector(57120, 16),
57600 => conv_std_logic_vector(0, 16),
57601 => conv_std_logic_vector(225, 16),
57602 => conv_std_logic_vector(450, 16),
57603 => conv_std_logic_vector(675, 16),
57604 => conv_std_logic_vector(900, 16),
57605 => conv_std_logic_vector(1125, 16),
57606 => conv_std_logic_vector(1350, 16),
57607 => conv_std_logic_vector(1575, 16),
57608 => conv_std_logic_vector(1800, 16),
57609 => conv_std_logic_vector(2025, 16),
57610 => conv_std_logic_vector(2250, 16),
57611 => conv_std_logic_vector(2475, 16),
57612 => conv_std_logic_vector(2700, 16),
57613 => conv_std_logic_vector(2925, 16),
57614 => conv_std_logic_vector(3150, 16),
57615 => conv_std_logic_vector(3375, 16),
57616 => conv_std_logic_vector(3600, 16),
57617 => conv_std_logic_vector(3825, 16),
57618 => conv_std_logic_vector(4050, 16),
57619 => conv_std_logic_vector(4275, 16),
57620 => conv_std_logic_vector(4500, 16),
57621 => conv_std_logic_vector(4725, 16),
57622 => conv_std_logic_vector(4950, 16),
57623 => conv_std_logic_vector(5175, 16),
57624 => conv_std_logic_vector(5400, 16),
57625 => conv_std_logic_vector(5625, 16),
57626 => conv_std_logic_vector(5850, 16),
57627 => conv_std_logic_vector(6075, 16),
57628 => conv_std_logic_vector(6300, 16),
57629 => conv_std_logic_vector(6525, 16),
57630 => conv_std_logic_vector(6750, 16),
57631 => conv_std_logic_vector(6975, 16),
57632 => conv_std_logic_vector(7200, 16),
57633 => conv_std_logic_vector(7425, 16),
57634 => conv_std_logic_vector(7650, 16),
57635 => conv_std_logic_vector(7875, 16),
57636 => conv_std_logic_vector(8100, 16),
57637 => conv_std_logic_vector(8325, 16),
57638 => conv_std_logic_vector(8550, 16),
57639 => conv_std_logic_vector(8775, 16),
57640 => conv_std_logic_vector(9000, 16),
57641 => conv_std_logic_vector(9225, 16),
57642 => conv_std_logic_vector(9450, 16),
57643 => conv_std_logic_vector(9675, 16),
57644 => conv_std_logic_vector(9900, 16),
57645 => conv_std_logic_vector(10125, 16),
57646 => conv_std_logic_vector(10350, 16),
57647 => conv_std_logic_vector(10575, 16),
57648 => conv_std_logic_vector(10800, 16),
57649 => conv_std_logic_vector(11025, 16),
57650 => conv_std_logic_vector(11250, 16),
57651 => conv_std_logic_vector(11475, 16),
57652 => conv_std_logic_vector(11700, 16),
57653 => conv_std_logic_vector(11925, 16),
57654 => conv_std_logic_vector(12150, 16),
57655 => conv_std_logic_vector(12375, 16),
57656 => conv_std_logic_vector(12600, 16),
57657 => conv_std_logic_vector(12825, 16),
57658 => conv_std_logic_vector(13050, 16),
57659 => conv_std_logic_vector(13275, 16),
57660 => conv_std_logic_vector(13500, 16),
57661 => conv_std_logic_vector(13725, 16),
57662 => conv_std_logic_vector(13950, 16),
57663 => conv_std_logic_vector(14175, 16),
57664 => conv_std_logic_vector(14400, 16),
57665 => conv_std_logic_vector(14625, 16),
57666 => conv_std_logic_vector(14850, 16),
57667 => conv_std_logic_vector(15075, 16),
57668 => conv_std_logic_vector(15300, 16),
57669 => conv_std_logic_vector(15525, 16),
57670 => conv_std_logic_vector(15750, 16),
57671 => conv_std_logic_vector(15975, 16),
57672 => conv_std_logic_vector(16200, 16),
57673 => conv_std_logic_vector(16425, 16),
57674 => conv_std_logic_vector(16650, 16),
57675 => conv_std_logic_vector(16875, 16),
57676 => conv_std_logic_vector(17100, 16),
57677 => conv_std_logic_vector(17325, 16),
57678 => conv_std_logic_vector(17550, 16),
57679 => conv_std_logic_vector(17775, 16),
57680 => conv_std_logic_vector(18000, 16),
57681 => conv_std_logic_vector(18225, 16),
57682 => conv_std_logic_vector(18450, 16),
57683 => conv_std_logic_vector(18675, 16),
57684 => conv_std_logic_vector(18900, 16),
57685 => conv_std_logic_vector(19125, 16),
57686 => conv_std_logic_vector(19350, 16),
57687 => conv_std_logic_vector(19575, 16),
57688 => conv_std_logic_vector(19800, 16),
57689 => conv_std_logic_vector(20025, 16),
57690 => conv_std_logic_vector(20250, 16),
57691 => conv_std_logic_vector(20475, 16),
57692 => conv_std_logic_vector(20700, 16),
57693 => conv_std_logic_vector(20925, 16),
57694 => conv_std_logic_vector(21150, 16),
57695 => conv_std_logic_vector(21375, 16),
57696 => conv_std_logic_vector(21600, 16),
57697 => conv_std_logic_vector(21825, 16),
57698 => conv_std_logic_vector(22050, 16),
57699 => conv_std_logic_vector(22275, 16),
57700 => conv_std_logic_vector(22500, 16),
57701 => conv_std_logic_vector(22725, 16),
57702 => conv_std_logic_vector(22950, 16),
57703 => conv_std_logic_vector(23175, 16),
57704 => conv_std_logic_vector(23400, 16),
57705 => conv_std_logic_vector(23625, 16),
57706 => conv_std_logic_vector(23850, 16),
57707 => conv_std_logic_vector(24075, 16),
57708 => conv_std_logic_vector(24300, 16),
57709 => conv_std_logic_vector(24525, 16),
57710 => conv_std_logic_vector(24750, 16),
57711 => conv_std_logic_vector(24975, 16),
57712 => conv_std_logic_vector(25200, 16),
57713 => conv_std_logic_vector(25425, 16),
57714 => conv_std_logic_vector(25650, 16),
57715 => conv_std_logic_vector(25875, 16),
57716 => conv_std_logic_vector(26100, 16),
57717 => conv_std_logic_vector(26325, 16),
57718 => conv_std_logic_vector(26550, 16),
57719 => conv_std_logic_vector(26775, 16),
57720 => conv_std_logic_vector(27000, 16),
57721 => conv_std_logic_vector(27225, 16),
57722 => conv_std_logic_vector(27450, 16),
57723 => conv_std_logic_vector(27675, 16),
57724 => conv_std_logic_vector(27900, 16),
57725 => conv_std_logic_vector(28125, 16),
57726 => conv_std_logic_vector(28350, 16),
57727 => conv_std_logic_vector(28575, 16),
57728 => conv_std_logic_vector(28800, 16),
57729 => conv_std_logic_vector(29025, 16),
57730 => conv_std_logic_vector(29250, 16),
57731 => conv_std_logic_vector(29475, 16),
57732 => conv_std_logic_vector(29700, 16),
57733 => conv_std_logic_vector(29925, 16),
57734 => conv_std_logic_vector(30150, 16),
57735 => conv_std_logic_vector(30375, 16),
57736 => conv_std_logic_vector(30600, 16),
57737 => conv_std_logic_vector(30825, 16),
57738 => conv_std_logic_vector(31050, 16),
57739 => conv_std_logic_vector(31275, 16),
57740 => conv_std_logic_vector(31500, 16),
57741 => conv_std_logic_vector(31725, 16),
57742 => conv_std_logic_vector(31950, 16),
57743 => conv_std_logic_vector(32175, 16),
57744 => conv_std_logic_vector(32400, 16),
57745 => conv_std_logic_vector(32625, 16),
57746 => conv_std_logic_vector(32850, 16),
57747 => conv_std_logic_vector(33075, 16),
57748 => conv_std_logic_vector(33300, 16),
57749 => conv_std_logic_vector(33525, 16),
57750 => conv_std_logic_vector(33750, 16),
57751 => conv_std_logic_vector(33975, 16),
57752 => conv_std_logic_vector(34200, 16),
57753 => conv_std_logic_vector(34425, 16),
57754 => conv_std_logic_vector(34650, 16),
57755 => conv_std_logic_vector(34875, 16),
57756 => conv_std_logic_vector(35100, 16),
57757 => conv_std_logic_vector(35325, 16),
57758 => conv_std_logic_vector(35550, 16),
57759 => conv_std_logic_vector(35775, 16),
57760 => conv_std_logic_vector(36000, 16),
57761 => conv_std_logic_vector(36225, 16),
57762 => conv_std_logic_vector(36450, 16),
57763 => conv_std_logic_vector(36675, 16),
57764 => conv_std_logic_vector(36900, 16),
57765 => conv_std_logic_vector(37125, 16),
57766 => conv_std_logic_vector(37350, 16),
57767 => conv_std_logic_vector(37575, 16),
57768 => conv_std_logic_vector(37800, 16),
57769 => conv_std_logic_vector(38025, 16),
57770 => conv_std_logic_vector(38250, 16),
57771 => conv_std_logic_vector(38475, 16),
57772 => conv_std_logic_vector(38700, 16),
57773 => conv_std_logic_vector(38925, 16),
57774 => conv_std_logic_vector(39150, 16),
57775 => conv_std_logic_vector(39375, 16),
57776 => conv_std_logic_vector(39600, 16),
57777 => conv_std_logic_vector(39825, 16),
57778 => conv_std_logic_vector(40050, 16),
57779 => conv_std_logic_vector(40275, 16),
57780 => conv_std_logic_vector(40500, 16),
57781 => conv_std_logic_vector(40725, 16),
57782 => conv_std_logic_vector(40950, 16),
57783 => conv_std_logic_vector(41175, 16),
57784 => conv_std_logic_vector(41400, 16),
57785 => conv_std_logic_vector(41625, 16),
57786 => conv_std_logic_vector(41850, 16),
57787 => conv_std_logic_vector(42075, 16),
57788 => conv_std_logic_vector(42300, 16),
57789 => conv_std_logic_vector(42525, 16),
57790 => conv_std_logic_vector(42750, 16),
57791 => conv_std_logic_vector(42975, 16),
57792 => conv_std_logic_vector(43200, 16),
57793 => conv_std_logic_vector(43425, 16),
57794 => conv_std_logic_vector(43650, 16),
57795 => conv_std_logic_vector(43875, 16),
57796 => conv_std_logic_vector(44100, 16),
57797 => conv_std_logic_vector(44325, 16),
57798 => conv_std_logic_vector(44550, 16),
57799 => conv_std_logic_vector(44775, 16),
57800 => conv_std_logic_vector(45000, 16),
57801 => conv_std_logic_vector(45225, 16),
57802 => conv_std_logic_vector(45450, 16),
57803 => conv_std_logic_vector(45675, 16),
57804 => conv_std_logic_vector(45900, 16),
57805 => conv_std_logic_vector(46125, 16),
57806 => conv_std_logic_vector(46350, 16),
57807 => conv_std_logic_vector(46575, 16),
57808 => conv_std_logic_vector(46800, 16),
57809 => conv_std_logic_vector(47025, 16),
57810 => conv_std_logic_vector(47250, 16),
57811 => conv_std_logic_vector(47475, 16),
57812 => conv_std_logic_vector(47700, 16),
57813 => conv_std_logic_vector(47925, 16),
57814 => conv_std_logic_vector(48150, 16),
57815 => conv_std_logic_vector(48375, 16),
57816 => conv_std_logic_vector(48600, 16),
57817 => conv_std_logic_vector(48825, 16),
57818 => conv_std_logic_vector(49050, 16),
57819 => conv_std_logic_vector(49275, 16),
57820 => conv_std_logic_vector(49500, 16),
57821 => conv_std_logic_vector(49725, 16),
57822 => conv_std_logic_vector(49950, 16),
57823 => conv_std_logic_vector(50175, 16),
57824 => conv_std_logic_vector(50400, 16),
57825 => conv_std_logic_vector(50625, 16),
57826 => conv_std_logic_vector(50850, 16),
57827 => conv_std_logic_vector(51075, 16),
57828 => conv_std_logic_vector(51300, 16),
57829 => conv_std_logic_vector(51525, 16),
57830 => conv_std_logic_vector(51750, 16),
57831 => conv_std_logic_vector(51975, 16),
57832 => conv_std_logic_vector(52200, 16),
57833 => conv_std_logic_vector(52425, 16),
57834 => conv_std_logic_vector(52650, 16),
57835 => conv_std_logic_vector(52875, 16),
57836 => conv_std_logic_vector(53100, 16),
57837 => conv_std_logic_vector(53325, 16),
57838 => conv_std_logic_vector(53550, 16),
57839 => conv_std_logic_vector(53775, 16),
57840 => conv_std_logic_vector(54000, 16),
57841 => conv_std_logic_vector(54225, 16),
57842 => conv_std_logic_vector(54450, 16),
57843 => conv_std_logic_vector(54675, 16),
57844 => conv_std_logic_vector(54900, 16),
57845 => conv_std_logic_vector(55125, 16),
57846 => conv_std_logic_vector(55350, 16),
57847 => conv_std_logic_vector(55575, 16),
57848 => conv_std_logic_vector(55800, 16),
57849 => conv_std_logic_vector(56025, 16),
57850 => conv_std_logic_vector(56250, 16),
57851 => conv_std_logic_vector(56475, 16),
57852 => conv_std_logic_vector(56700, 16),
57853 => conv_std_logic_vector(56925, 16),
57854 => conv_std_logic_vector(57150, 16),
57855 => conv_std_logic_vector(57375, 16),
57856 => conv_std_logic_vector(0, 16),
57857 => conv_std_logic_vector(226, 16),
57858 => conv_std_logic_vector(452, 16),
57859 => conv_std_logic_vector(678, 16),
57860 => conv_std_logic_vector(904, 16),
57861 => conv_std_logic_vector(1130, 16),
57862 => conv_std_logic_vector(1356, 16),
57863 => conv_std_logic_vector(1582, 16),
57864 => conv_std_logic_vector(1808, 16),
57865 => conv_std_logic_vector(2034, 16),
57866 => conv_std_logic_vector(2260, 16),
57867 => conv_std_logic_vector(2486, 16),
57868 => conv_std_logic_vector(2712, 16),
57869 => conv_std_logic_vector(2938, 16),
57870 => conv_std_logic_vector(3164, 16),
57871 => conv_std_logic_vector(3390, 16),
57872 => conv_std_logic_vector(3616, 16),
57873 => conv_std_logic_vector(3842, 16),
57874 => conv_std_logic_vector(4068, 16),
57875 => conv_std_logic_vector(4294, 16),
57876 => conv_std_logic_vector(4520, 16),
57877 => conv_std_logic_vector(4746, 16),
57878 => conv_std_logic_vector(4972, 16),
57879 => conv_std_logic_vector(5198, 16),
57880 => conv_std_logic_vector(5424, 16),
57881 => conv_std_logic_vector(5650, 16),
57882 => conv_std_logic_vector(5876, 16),
57883 => conv_std_logic_vector(6102, 16),
57884 => conv_std_logic_vector(6328, 16),
57885 => conv_std_logic_vector(6554, 16),
57886 => conv_std_logic_vector(6780, 16),
57887 => conv_std_logic_vector(7006, 16),
57888 => conv_std_logic_vector(7232, 16),
57889 => conv_std_logic_vector(7458, 16),
57890 => conv_std_logic_vector(7684, 16),
57891 => conv_std_logic_vector(7910, 16),
57892 => conv_std_logic_vector(8136, 16),
57893 => conv_std_logic_vector(8362, 16),
57894 => conv_std_logic_vector(8588, 16),
57895 => conv_std_logic_vector(8814, 16),
57896 => conv_std_logic_vector(9040, 16),
57897 => conv_std_logic_vector(9266, 16),
57898 => conv_std_logic_vector(9492, 16),
57899 => conv_std_logic_vector(9718, 16),
57900 => conv_std_logic_vector(9944, 16),
57901 => conv_std_logic_vector(10170, 16),
57902 => conv_std_logic_vector(10396, 16),
57903 => conv_std_logic_vector(10622, 16),
57904 => conv_std_logic_vector(10848, 16),
57905 => conv_std_logic_vector(11074, 16),
57906 => conv_std_logic_vector(11300, 16),
57907 => conv_std_logic_vector(11526, 16),
57908 => conv_std_logic_vector(11752, 16),
57909 => conv_std_logic_vector(11978, 16),
57910 => conv_std_logic_vector(12204, 16),
57911 => conv_std_logic_vector(12430, 16),
57912 => conv_std_logic_vector(12656, 16),
57913 => conv_std_logic_vector(12882, 16),
57914 => conv_std_logic_vector(13108, 16),
57915 => conv_std_logic_vector(13334, 16),
57916 => conv_std_logic_vector(13560, 16),
57917 => conv_std_logic_vector(13786, 16),
57918 => conv_std_logic_vector(14012, 16),
57919 => conv_std_logic_vector(14238, 16),
57920 => conv_std_logic_vector(14464, 16),
57921 => conv_std_logic_vector(14690, 16),
57922 => conv_std_logic_vector(14916, 16),
57923 => conv_std_logic_vector(15142, 16),
57924 => conv_std_logic_vector(15368, 16),
57925 => conv_std_logic_vector(15594, 16),
57926 => conv_std_logic_vector(15820, 16),
57927 => conv_std_logic_vector(16046, 16),
57928 => conv_std_logic_vector(16272, 16),
57929 => conv_std_logic_vector(16498, 16),
57930 => conv_std_logic_vector(16724, 16),
57931 => conv_std_logic_vector(16950, 16),
57932 => conv_std_logic_vector(17176, 16),
57933 => conv_std_logic_vector(17402, 16),
57934 => conv_std_logic_vector(17628, 16),
57935 => conv_std_logic_vector(17854, 16),
57936 => conv_std_logic_vector(18080, 16),
57937 => conv_std_logic_vector(18306, 16),
57938 => conv_std_logic_vector(18532, 16),
57939 => conv_std_logic_vector(18758, 16),
57940 => conv_std_logic_vector(18984, 16),
57941 => conv_std_logic_vector(19210, 16),
57942 => conv_std_logic_vector(19436, 16),
57943 => conv_std_logic_vector(19662, 16),
57944 => conv_std_logic_vector(19888, 16),
57945 => conv_std_logic_vector(20114, 16),
57946 => conv_std_logic_vector(20340, 16),
57947 => conv_std_logic_vector(20566, 16),
57948 => conv_std_logic_vector(20792, 16),
57949 => conv_std_logic_vector(21018, 16),
57950 => conv_std_logic_vector(21244, 16),
57951 => conv_std_logic_vector(21470, 16),
57952 => conv_std_logic_vector(21696, 16),
57953 => conv_std_logic_vector(21922, 16),
57954 => conv_std_logic_vector(22148, 16),
57955 => conv_std_logic_vector(22374, 16),
57956 => conv_std_logic_vector(22600, 16),
57957 => conv_std_logic_vector(22826, 16),
57958 => conv_std_logic_vector(23052, 16),
57959 => conv_std_logic_vector(23278, 16),
57960 => conv_std_logic_vector(23504, 16),
57961 => conv_std_logic_vector(23730, 16),
57962 => conv_std_logic_vector(23956, 16),
57963 => conv_std_logic_vector(24182, 16),
57964 => conv_std_logic_vector(24408, 16),
57965 => conv_std_logic_vector(24634, 16),
57966 => conv_std_logic_vector(24860, 16),
57967 => conv_std_logic_vector(25086, 16),
57968 => conv_std_logic_vector(25312, 16),
57969 => conv_std_logic_vector(25538, 16),
57970 => conv_std_logic_vector(25764, 16),
57971 => conv_std_logic_vector(25990, 16),
57972 => conv_std_logic_vector(26216, 16),
57973 => conv_std_logic_vector(26442, 16),
57974 => conv_std_logic_vector(26668, 16),
57975 => conv_std_logic_vector(26894, 16),
57976 => conv_std_logic_vector(27120, 16),
57977 => conv_std_logic_vector(27346, 16),
57978 => conv_std_logic_vector(27572, 16),
57979 => conv_std_logic_vector(27798, 16),
57980 => conv_std_logic_vector(28024, 16),
57981 => conv_std_logic_vector(28250, 16),
57982 => conv_std_logic_vector(28476, 16),
57983 => conv_std_logic_vector(28702, 16),
57984 => conv_std_logic_vector(28928, 16),
57985 => conv_std_logic_vector(29154, 16),
57986 => conv_std_logic_vector(29380, 16),
57987 => conv_std_logic_vector(29606, 16),
57988 => conv_std_logic_vector(29832, 16),
57989 => conv_std_logic_vector(30058, 16),
57990 => conv_std_logic_vector(30284, 16),
57991 => conv_std_logic_vector(30510, 16),
57992 => conv_std_logic_vector(30736, 16),
57993 => conv_std_logic_vector(30962, 16),
57994 => conv_std_logic_vector(31188, 16),
57995 => conv_std_logic_vector(31414, 16),
57996 => conv_std_logic_vector(31640, 16),
57997 => conv_std_logic_vector(31866, 16),
57998 => conv_std_logic_vector(32092, 16),
57999 => conv_std_logic_vector(32318, 16),
58000 => conv_std_logic_vector(32544, 16),
58001 => conv_std_logic_vector(32770, 16),
58002 => conv_std_logic_vector(32996, 16),
58003 => conv_std_logic_vector(33222, 16),
58004 => conv_std_logic_vector(33448, 16),
58005 => conv_std_logic_vector(33674, 16),
58006 => conv_std_logic_vector(33900, 16),
58007 => conv_std_logic_vector(34126, 16),
58008 => conv_std_logic_vector(34352, 16),
58009 => conv_std_logic_vector(34578, 16),
58010 => conv_std_logic_vector(34804, 16),
58011 => conv_std_logic_vector(35030, 16),
58012 => conv_std_logic_vector(35256, 16),
58013 => conv_std_logic_vector(35482, 16),
58014 => conv_std_logic_vector(35708, 16),
58015 => conv_std_logic_vector(35934, 16),
58016 => conv_std_logic_vector(36160, 16),
58017 => conv_std_logic_vector(36386, 16),
58018 => conv_std_logic_vector(36612, 16),
58019 => conv_std_logic_vector(36838, 16),
58020 => conv_std_logic_vector(37064, 16),
58021 => conv_std_logic_vector(37290, 16),
58022 => conv_std_logic_vector(37516, 16),
58023 => conv_std_logic_vector(37742, 16),
58024 => conv_std_logic_vector(37968, 16),
58025 => conv_std_logic_vector(38194, 16),
58026 => conv_std_logic_vector(38420, 16),
58027 => conv_std_logic_vector(38646, 16),
58028 => conv_std_logic_vector(38872, 16),
58029 => conv_std_logic_vector(39098, 16),
58030 => conv_std_logic_vector(39324, 16),
58031 => conv_std_logic_vector(39550, 16),
58032 => conv_std_logic_vector(39776, 16),
58033 => conv_std_logic_vector(40002, 16),
58034 => conv_std_logic_vector(40228, 16),
58035 => conv_std_logic_vector(40454, 16),
58036 => conv_std_logic_vector(40680, 16),
58037 => conv_std_logic_vector(40906, 16),
58038 => conv_std_logic_vector(41132, 16),
58039 => conv_std_logic_vector(41358, 16),
58040 => conv_std_logic_vector(41584, 16),
58041 => conv_std_logic_vector(41810, 16),
58042 => conv_std_logic_vector(42036, 16),
58043 => conv_std_logic_vector(42262, 16),
58044 => conv_std_logic_vector(42488, 16),
58045 => conv_std_logic_vector(42714, 16),
58046 => conv_std_logic_vector(42940, 16),
58047 => conv_std_logic_vector(43166, 16),
58048 => conv_std_logic_vector(43392, 16),
58049 => conv_std_logic_vector(43618, 16),
58050 => conv_std_logic_vector(43844, 16),
58051 => conv_std_logic_vector(44070, 16),
58052 => conv_std_logic_vector(44296, 16),
58053 => conv_std_logic_vector(44522, 16),
58054 => conv_std_logic_vector(44748, 16),
58055 => conv_std_logic_vector(44974, 16),
58056 => conv_std_logic_vector(45200, 16),
58057 => conv_std_logic_vector(45426, 16),
58058 => conv_std_logic_vector(45652, 16),
58059 => conv_std_logic_vector(45878, 16),
58060 => conv_std_logic_vector(46104, 16),
58061 => conv_std_logic_vector(46330, 16),
58062 => conv_std_logic_vector(46556, 16),
58063 => conv_std_logic_vector(46782, 16),
58064 => conv_std_logic_vector(47008, 16),
58065 => conv_std_logic_vector(47234, 16),
58066 => conv_std_logic_vector(47460, 16),
58067 => conv_std_logic_vector(47686, 16),
58068 => conv_std_logic_vector(47912, 16),
58069 => conv_std_logic_vector(48138, 16),
58070 => conv_std_logic_vector(48364, 16),
58071 => conv_std_logic_vector(48590, 16),
58072 => conv_std_logic_vector(48816, 16),
58073 => conv_std_logic_vector(49042, 16),
58074 => conv_std_logic_vector(49268, 16),
58075 => conv_std_logic_vector(49494, 16),
58076 => conv_std_logic_vector(49720, 16),
58077 => conv_std_logic_vector(49946, 16),
58078 => conv_std_logic_vector(50172, 16),
58079 => conv_std_logic_vector(50398, 16),
58080 => conv_std_logic_vector(50624, 16),
58081 => conv_std_logic_vector(50850, 16),
58082 => conv_std_logic_vector(51076, 16),
58083 => conv_std_logic_vector(51302, 16),
58084 => conv_std_logic_vector(51528, 16),
58085 => conv_std_logic_vector(51754, 16),
58086 => conv_std_logic_vector(51980, 16),
58087 => conv_std_logic_vector(52206, 16),
58088 => conv_std_logic_vector(52432, 16),
58089 => conv_std_logic_vector(52658, 16),
58090 => conv_std_logic_vector(52884, 16),
58091 => conv_std_logic_vector(53110, 16),
58092 => conv_std_logic_vector(53336, 16),
58093 => conv_std_logic_vector(53562, 16),
58094 => conv_std_logic_vector(53788, 16),
58095 => conv_std_logic_vector(54014, 16),
58096 => conv_std_logic_vector(54240, 16),
58097 => conv_std_logic_vector(54466, 16),
58098 => conv_std_logic_vector(54692, 16),
58099 => conv_std_logic_vector(54918, 16),
58100 => conv_std_logic_vector(55144, 16),
58101 => conv_std_logic_vector(55370, 16),
58102 => conv_std_logic_vector(55596, 16),
58103 => conv_std_logic_vector(55822, 16),
58104 => conv_std_logic_vector(56048, 16),
58105 => conv_std_logic_vector(56274, 16),
58106 => conv_std_logic_vector(56500, 16),
58107 => conv_std_logic_vector(56726, 16),
58108 => conv_std_logic_vector(56952, 16),
58109 => conv_std_logic_vector(57178, 16),
58110 => conv_std_logic_vector(57404, 16),
58111 => conv_std_logic_vector(57630, 16),
58112 => conv_std_logic_vector(0, 16),
58113 => conv_std_logic_vector(227, 16),
58114 => conv_std_logic_vector(454, 16),
58115 => conv_std_logic_vector(681, 16),
58116 => conv_std_logic_vector(908, 16),
58117 => conv_std_logic_vector(1135, 16),
58118 => conv_std_logic_vector(1362, 16),
58119 => conv_std_logic_vector(1589, 16),
58120 => conv_std_logic_vector(1816, 16),
58121 => conv_std_logic_vector(2043, 16),
58122 => conv_std_logic_vector(2270, 16),
58123 => conv_std_logic_vector(2497, 16),
58124 => conv_std_logic_vector(2724, 16),
58125 => conv_std_logic_vector(2951, 16),
58126 => conv_std_logic_vector(3178, 16),
58127 => conv_std_logic_vector(3405, 16),
58128 => conv_std_logic_vector(3632, 16),
58129 => conv_std_logic_vector(3859, 16),
58130 => conv_std_logic_vector(4086, 16),
58131 => conv_std_logic_vector(4313, 16),
58132 => conv_std_logic_vector(4540, 16),
58133 => conv_std_logic_vector(4767, 16),
58134 => conv_std_logic_vector(4994, 16),
58135 => conv_std_logic_vector(5221, 16),
58136 => conv_std_logic_vector(5448, 16),
58137 => conv_std_logic_vector(5675, 16),
58138 => conv_std_logic_vector(5902, 16),
58139 => conv_std_logic_vector(6129, 16),
58140 => conv_std_logic_vector(6356, 16),
58141 => conv_std_logic_vector(6583, 16),
58142 => conv_std_logic_vector(6810, 16),
58143 => conv_std_logic_vector(7037, 16),
58144 => conv_std_logic_vector(7264, 16),
58145 => conv_std_logic_vector(7491, 16),
58146 => conv_std_logic_vector(7718, 16),
58147 => conv_std_logic_vector(7945, 16),
58148 => conv_std_logic_vector(8172, 16),
58149 => conv_std_logic_vector(8399, 16),
58150 => conv_std_logic_vector(8626, 16),
58151 => conv_std_logic_vector(8853, 16),
58152 => conv_std_logic_vector(9080, 16),
58153 => conv_std_logic_vector(9307, 16),
58154 => conv_std_logic_vector(9534, 16),
58155 => conv_std_logic_vector(9761, 16),
58156 => conv_std_logic_vector(9988, 16),
58157 => conv_std_logic_vector(10215, 16),
58158 => conv_std_logic_vector(10442, 16),
58159 => conv_std_logic_vector(10669, 16),
58160 => conv_std_logic_vector(10896, 16),
58161 => conv_std_logic_vector(11123, 16),
58162 => conv_std_logic_vector(11350, 16),
58163 => conv_std_logic_vector(11577, 16),
58164 => conv_std_logic_vector(11804, 16),
58165 => conv_std_logic_vector(12031, 16),
58166 => conv_std_logic_vector(12258, 16),
58167 => conv_std_logic_vector(12485, 16),
58168 => conv_std_logic_vector(12712, 16),
58169 => conv_std_logic_vector(12939, 16),
58170 => conv_std_logic_vector(13166, 16),
58171 => conv_std_logic_vector(13393, 16),
58172 => conv_std_logic_vector(13620, 16),
58173 => conv_std_logic_vector(13847, 16),
58174 => conv_std_logic_vector(14074, 16),
58175 => conv_std_logic_vector(14301, 16),
58176 => conv_std_logic_vector(14528, 16),
58177 => conv_std_logic_vector(14755, 16),
58178 => conv_std_logic_vector(14982, 16),
58179 => conv_std_logic_vector(15209, 16),
58180 => conv_std_logic_vector(15436, 16),
58181 => conv_std_logic_vector(15663, 16),
58182 => conv_std_logic_vector(15890, 16),
58183 => conv_std_logic_vector(16117, 16),
58184 => conv_std_logic_vector(16344, 16),
58185 => conv_std_logic_vector(16571, 16),
58186 => conv_std_logic_vector(16798, 16),
58187 => conv_std_logic_vector(17025, 16),
58188 => conv_std_logic_vector(17252, 16),
58189 => conv_std_logic_vector(17479, 16),
58190 => conv_std_logic_vector(17706, 16),
58191 => conv_std_logic_vector(17933, 16),
58192 => conv_std_logic_vector(18160, 16),
58193 => conv_std_logic_vector(18387, 16),
58194 => conv_std_logic_vector(18614, 16),
58195 => conv_std_logic_vector(18841, 16),
58196 => conv_std_logic_vector(19068, 16),
58197 => conv_std_logic_vector(19295, 16),
58198 => conv_std_logic_vector(19522, 16),
58199 => conv_std_logic_vector(19749, 16),
58200 => conv_std_logic_vector(19976, 16),
58201 => conv_std_logic_vector(20203, 16),
58202 => conv_std_logic_vector(20430, 16),
58203 => conv_std_logic_vector(20657, 16),
58204 => conv_std_logic_vector(20884, 16),
58205 => conv_std_logic_vector(21111, 16),
58206 => conv_std_logic_vector(21338, 16),
58207 => conv_std_logic_vector(21565, 16),
58208 => conv_std_logic_vector(21792, 16),
58209 => conv_std_logic_vector(22019, 16),
58210 => conv_std_logic_vector(22246, 16),
58211 => conv_std_logic_vector(22473, 16),
58212 => conv_std_logic_vector(22700, 16),
58213 => conv_std_logic_vector(22927, 16),
58214 => conv_std_logic_vector(23154, 16),
58215 => conv_std_logic_vector(23381, 16),
58216 => conv_std_logic_vector(23608, 16),
58217 => conv_std_logic_vector(23835, 16),
58218 => conv_std_logic_vector(24062, 16),
58219 => conv_std_logic_vector(24289, 16),
58220 => conv_std_logic_vector(24516, 16),
58221 => conv_std_logic_vector(24743, 16),
58222 => conv_std_logic_vector(24970, 16),
58223 => conv_std_logic_vector(25197, 16),
58224 => conv_std_logic_vector(25424, 16),
58225 => conv_std_logic_vector(25651, 16),
58226 => conv_std_logic_vector(25878, 16),
58227 => conv_std_logic_vector(26105, 16),
58228 => conv_std_logic_vector(26332, 16),
58229 => conv_std_logic_vector(26559, 16),
58230 => conv_std_logic_vector(26786, 16),
58231 => conv_std_logic_vector(27013, 16),
58232 => conv_std_logic_vector(27240, 16),
58233 => conv_std_logic_vector(27467, 16),
58234 => conv_std_logic_vector(27694, 16),
58235 => conv_std_logic_vector(27921, 16),
58236 => conv_std_logic_vector(28148, 16),
58237 => conv_std_logic_vector(28375, 16),
58238 => conv_std_logic_vector(28602, 16),
58239 => conv_std_logic_vector(28829, 16),
58240 => conv_std_logic_vector(29056, 16),
58241 => conv_std_logic_vector(29283, 16),
58242 => conv_std_logic_vector(29510, 16),
58243 => conv_std_logic_vector(29737, 16),
58244 => conv_std_logic_vector(29964, 16),
58245 => conv_std_logic_vector(30191, 16),
58246 => conv_std_logic_vector(30418, 16),
58247 => conv_std_logic_vector(30645, 16),
58248 => conv_std_logic_vector(30872, 16),
58249 => conv_std_logic_vector(31099, 16),
58250 => conv_std_logic_vector(31326, 16),
58251 => conv_std_logic_vector(31553, 16),
58252 => conv_std_logic_vector(31780, 16),
58253 => conv_std_logic_vector(32007, 16),
58254 => conv_std_logic_vector(32234, 16),
58255 => conv_std_logic_vector(32461, 16),
58256 => conv_std_logic_vector(32688, 16),
58257 => conv_std_logic_vector(32915, 16),
58258 => conv_std_logic_vector(33142, 16),
58259 => conv_std_logic_vector(33369, 16),
58260 => conv_std_logic_vector(33596, 16),
58261 => conv_std_logic_vector(33823, 16),
58262 => conv_std_logic_vector(34050, 16),
58263 => conv_std_logic_vector(34277, 16),
58264 => conv_std_logic_vector(34504, 16),
58265 => conv_std_logic_vector(34731, 16),
58266 => conv_std_logic_vector(34958, 16),
58267 => conv_std_logic_vector(35185, 16),
58268 => conv_std_logic_vector(35412, 16),
58269 => conv_std_logic_vector(35639, 16),
58270 => conv_std_logic_vector(35866, 16),
58271 => conv_std_logic_vector(36093, 16),
58272 => conv_std_logic_vector(36320, 16),
58273 => conv_std_logic_vector(36547, 16),
58274 => conv_std_logic_vector(36774, 16),
58275 => conv_std_logic_vector(37001, 16),
58276 => conv_std_logic_vector(37228, 16),
58277 => conv_std_logic_vector(37455, 16),
58278 => conv_std_logic_vector(37682, 16),
58279 => conv_std_logic_vector(37909, 16),
58280 => conv_std_logic_vector(38136, 16),
58281 => conv_std_logic_vector(38363, 16),
58282 => conv_std_logic_vector(38590, 16),
58283 => conv_std_logic_vector(38817, 16),
58284 => conv_std_logic_vector(39044, 16),
58285 => conv_std_logic_vector(39271, 16),
58286 => conv_std_logic_vector(39498, 16),
58287 => conv_std_logic_vector(39725, 16),
58288 => conv_std_logic_vector(39952, 16),
58289 => conv_std_logic_vector(40179, 16),
58290 => conv_std_logic_vector(40406, 16),
58291 => conv_std_logic_vector(40633, 16),
58292 => conv_std_logic_vector(40860, 16),
58293 => conv_std_logic_vector(41087, 16),
58294 => conv_std_logic_vector(41314, 16),
58295 => conv_std_logic_vector(41541, 16),
58296 => conv_std_logic_vector(41768, 16),
58297 => conv_std_logic_vector(41995, 16),
58298 => conv_std_logic_vector(42222, 16),
58299 => conv_std_logic_vector(42449, 16),
58300 => conv_std_logic_vector(42676, 16),
58301 => conv_std_logic_vector(42903, 16),
58302 => conv_std_logic_vector(43130, 16),
58303 => conv_std_logic_vector(43357, 16),
58304 => conv_std_logic_vector(43584, 16),
58305 => conv_std_logic_vector(43811, 16),
58306 => conv_std_logic_vector(44038, 16),
58307 => conv_std_logic_vector(44265, 16),
58308 => conv_std_logic_vector(44492, 16),
58309 => conv_std_logic_vector(44719, 16),
58310 => conv_std_logic_vector(44946, 16),
58311 => conv_std_logic_vector(45173, 16),
58312 => conv_std_logic_vector(45400, 16),
58313 => conv_std_logic_vector(45627, 16),
58314 => conv_std_logic_vector(45854, 16),
58315 => conv_std_logic_vector(46081, 16),
58316 => conv_std_logic_vector(46308, 16),
58317 => conv_std_logic_vector(46535, 16),
58318 => conv_std_logic_vector(46762, 16),
58319 => conv_std_logic_vector(46989, 16),
58320 => conv_std_logic_vector(47216, 16),
58321 => conv_std_logic_vector(47443, 16),
58322 => conv_std_logic_vector(47670, 16),
58323 => conv_std_logic_vector(47897, 16),
58324 => conv_std_logic_vector(48124, 16),
58325 => conv_std_logic_vector(48351, 16),
58326 => conv_std_logic_vector(48578, 16),
58327 => conv_std_logic_vector(48805, 16),
58328 => conv_std_logic_vector(49032, 16),
58329 => conv_std_logic_vector(49259, 16),
58330 => conv_std_logic_vector(49486, 16),
58331 => conv_std_logic_vector(49713, 16),
58332 => conv_std_logic_vector(49940, 16),
58333 => conv_std_logic_vector(50167, 16),
58334 => conv_std_logic_vector(50394, 16),
58335 => conv_std_logic_vector(50621, 16),
58336 => conv_std_logic_vector(50848, 16),
58337 => conv_std_logic_vector(51075, 16),
58338 => conv_std_logic_vector(51302, 16),
58339 => conv_std_logic_vector(51529, 16),
58340 => conv_std_logic_vector(51756, 16),
58341 => conv_std_logic_vector(51983, 16),
58342 => conv_std_logic_vector(52210, 16),
58343 => conv_std_logic_vector(52437, 16),
58344 => conv_std_logic_vector(52664, 16),
58345 => conv_std_logic_vector(52891, 16),
58346 => conv_std_logic_vector(53118, 16),
58347 => conv_std_logic_vector(53345, 16),
58348 => conv_std_logic_vector(53572, 16),
58349 => conv_std_logic_vector(53799, 16),
58350 => conv_std_logic_vector(54026, 16),
58351 => conv_std_logic_vector(54253, 16),
58352 => conv_std_logic_vector(54480, 16),
58353 => conv_std_logic_vector(54707, 16),
58354 => conv_std_logic_vector(54934, 16),
58355 => conv_std_logic_vector(55161, 16),
58356 => conv_std_logic_vector(55388, 16),
58357 => conv_std_logic_vector(55615, 16),
58358 => conv_std_logic_vector(55842, 16),
58359 => conv_std_logic_vector(56069, 16),
58360 => conv_std_logic_vector(56296, 16),
58361 => conv_std_logic_vector(56523, 16),
58362 => conv_std_logic_vector(56750, 16),
58363 => conv_std_logic_vector(56977, 16),
58364 => conv_std_logic_vector(57204, 16),
58365 => conv_std_logic_vector(57431, 16),
58366 => conv_std_logic_vector(57658, 16),
58367 => conv_std_logic_vector(57885, 16),
58368 => conv_std_logic_vector(0, 16),
58369 => conv_std_logic_vector(228, 16),
58370 => conv_std_logic_vector(456, 16),
58371 => conv_std_logic_vector(684, 16),
58372 => conv_std_logic_vector(912, 16),
58373 => conv_std_logic_vector(1140, 16),
58374 => conv_std_logic_vector(1368, 16),
58375 => conv_std_logic_vector(1596, 16),
58376 => conv_std_logic_vector(1824, 16),
58377 => conv_std_logic_vector(2052, 16),
58378 => conv_std_logic_vector(2280, 16),
58379 => conv_std_logic_vector(2508, 16),
58380 => conv_std_logic_vector(2736, 16),
58381 => conv_std_logic_vector(2964, 16),
58382 => conv_std_logic_vector(3192, 16),
58383 => conv_std_logic_vector(3420, 16),
58384 => conv_std_logic_vector(3648, 16),
58385 => conv_std_logic_vector(3876, 16),
58386 => conv_std_logic_vector(4104, 16),
58387 => conv_std_logic_vector(4332, 16),
58388 => conv_std_logic_vector(4560, 16),
58389 => conv_std_logic_vector(4788, 16),
58390 => conv_std_logic_vector(5016, 16),
58391 => conv_std_logic_vector(5244, 16),
58392 => conv_std_logic_vector(5472, 16),
58393 => conv_std_logic_vector(5700, 16),
58394 => conv_std_logic_vector(5928, 16),
58395 => conv_std_logic_vector(6156, 16),
58396 => conv_std_logic_vector(6384, 16),
58397 => conv_std_logic_vector(6612, 16),
58398 => conv_std_logic_vector(6840, 16),
58399 => conv_std_logic_vector(7068, 16),
58400 => conv_std_logic_vector(7296, 16),
58401 => conv_std_logic_vector(7524, 16),
58402 => conv_std_logic_vector(7752, 16),
58403 => conv_std_logic_vector(7980, 16),
58404 => conv_std_logic_vector(8208, 16),
58405 => conv_std_logic_vector(8436, 16),
58406 => conv_std_logic_vector(8664, 16),
58407 => conv_std_logic_vector(8892, 16),
58408 => conv_std_logic_vector(9120, 16),
58409 => conv_std_logic_vector(9348, 16),
58410 => conv_std_logic_vector(9576, 16),
58411 => conv_std_logic_vector(9804, 16),
58412 => conv_std_logic_vector(10032, 16),
58413 => conv_std_logic_vector(10260, 16),
58414 => conv_std_logic_vector(10488, 16),
58415 => conv_std_logic_vector(10716, 16),
58416 => conv_std_logic_vector(10944, 16),
58417 => conv_std_logic_vector(11172, 16),
58418 => conv_std_logic_vector(11400, 16),
58419 => conv_std_logic_vector(11628, 16),
58420 => conv_std_logic_vector(11856, 16),
58421 => conv_std_logic_vector(12084, 16),
58422 => conv_std_logic_vector(12312, 16),
58423 => conv_std_logic_vector(12540, 16),
58424 => conv_std_logic_vector(12768, 16),
58425 => conv_std_logic_vector(12996, 16),
58426 => conv_std_logic_vector(13224, 16),
58427 => conv_std_logic_vector(13452, 16),
58428 => conv_std_logic_vector(13680, 16),
58429 => conv_std_logic_vector(13908, 16),
58430 => conv_std_logic_vector(14136, 16),
58431 => conv_std_logic_vector(14364, 16),
58432 => conv_std_logic_vector(14592, 16),
58433 => conv_std_logic_vector(14820, 16),
58434 => conv_std_logic_vector(15048, 16),
58435 => conv_std_logic_vector(15276, 16),
58436 => conv_std_logic_vector(15504, 16),
58437 => conv_std_logic_vector(15732, 16),
58438 => conv_std_logic_vector(15960, 16),
58439 => conv_std_logic_vector(16188, 16),
58440 => conv_std_logic_vector(16416, 16),
58441 => conv_std_logic_vector(16644, 16),
58442 => conv_std_logic_vector(16872, 16),
58443 => conv_std_logic_vector(17100, 16),
58444 => conv_std_logic_vector(17328, 16),
58445 => conv_std_logic_vector(17556, 16),
58446 => conv_std_logic_vector(17784, 16),
58447 => conv_std_logic_vector(18012, 16),
58448 => conv_std_logic_vector(18240, 16),
58449 => conv_std_logic_vector(18468, 16),
58450 => conv_std_logic_vector(18696, 16),
58451 => conv_std_logic_vector(18924, 16),
58452 => conv_std_logic_vector(19152, 16),
58453 => conv_std_logic_vector(19380, 16),
58454 => conv_std_logic_vector(19608, 16),
58455 => conv_std_logic_vector(19836, 16),
58456 => conv_std_logic_vector(20064, 16),
58457 => conv_std_logic_vector(20292, 16),
58458 => conv_std_logic_vector(20520, 16),
58459 => conv_std_logic_vector(20748, 16),
58460 => conv_std_logic_vector(20976, 16),
58461 => conv_std_logic_vector(21204, 16),
58462 => conv_std_logic_vector(21432, 16),
58463 => conv_std_logic_vector(21660, 16),
58464 => conv_std_logic_vector(21888, 16),
58465 => conv_std_logic_vector(22116, 16),
58466 => conv_std_logic_vector(22344, 16),
58467 => conv_std_logic_vector(22572, 16),
58468 => conv_std_logic_vector(22800, 16),
58469 => conv_std_logic_vector(23028, 16),
58470 => conv_std_logic_vector(23256, 16),
58471 => conv_std_logic_vector(23484, 16),
58472 => conv_std_logic_vector(23712, 16),
58473 => conv_std_logic_vector(23940, 16),
58474 => conv_std_logic_vector(24168, 16),
58475 => conv_std_logic_vector(24396, 16),
58476 => conv_std_logic_vector(24624, 16),
58477 => conv_std_logic_vector(24852, 16),
58478 => conv_std_logic_vector(25080, 16),
58479 => conv_std_logic_vector(25308, 16),
58480 => conv_std_logic_vector(25536, 16),
58481 => conv_std_logic_vector(25764, 16),
58482 => conv_std_logic_vector(25992, 16),
58483 => conv_std_logic_vector(26220, 16),
58484 => conv_std_logic_vector(26448, 16),
58485 => conv_std_logic_vector(26676, 16),
58486 => conv_std_logic_vector(26904, 16),
58487 => conv_std_logic_vector(27132, 16),
58488 => conv_std_logic_vector(27360, 16),
58489 => conv_std_logic_vector(27588, 16),
58490 => conv_std_logic_vector(27816, 16),
58491 => conv_std_logic_vector(28044, 16),
58492 => conv_std_logic_vector(28272, 16),
58493 => conv_std_logic_vector(28500, 16),
58494 => conv_std_logic_vector(28728, 16),
58495 => conv_std_logic_vector(28956, 16),
58496 => conv_std_logic_vector(29184, 16),
58497 => conv_std_logic_vector(29412, 16),
58498 => conv_std_logic_vector(29640, 16),
58499 => conv_std_logic_vector(29868, 16),
58500 => conv_std_logic_vector(30096, 16),
58501 => conv_std_logic_vector(30324, 16),
58502 => conv_std_logic_vector(30552, 16),
58503 => conv_std_logic_vector(30780, 16),
58504 => conv_std_logic_vector(31008, 16),
58505 => conv_std_logic_vector(31236, 16),
58506 => conv_std_logic_vector(31464, 16),
58507 => conv_std_logic_vector(31692, 16),
58508 => conv_std_logic_vector(31920, 16),
58509 => conv_std_logic_vector(32148, 16),
58510 => conv_std_logic_vector(32376, 16),
58511 => conv_std_logic_vector(32604, 16),
58512 => conv_std_logic_vector(32832, 16),
58513 => conv_std_logic_vector(33060, 16),
58514 => conv_std_logic_vector(33288, 16),
58515 => conv_std_logic_vector(33516, 16),
58516 => conv_std_logic_vector(33744, 16),
58517 => conv_std_logic_vector(33972, 16),
58518 => conv_std_logic_vector(34200, 16),
58519 => conv_std_logic_vector(34428, 16),
58520 => conv_std_logic_vector(34656, 16),
58521 => conv_std_logic_vector(34884, 16),
58522 => conv_std_logic_vector(35112, 16),
58523 => conv_std_logic_vector(35340, 16),
58524 => conv_std_logic_vector(35568, 16),
58525 => conv_std_logic_vector(35796, 16),
58526 => conv_std_logic_vector(36024, 16),
58527 => conv_std_logic_vector(36252, 16),
58528 => conv_std_logic_vector(36480, 16),
58529 => conv_std_logic_vector(36708, 16),
58530 => conv_std_logic_vector(36936, 16),
58531 => conv_std_logic_vector(37164, 16),
58532 => conv_std_logic_vector(37392, 16),
58533 => conv_std_logic_vector(37620, 16),
58534 => conv_std_logic_vector(37848, 16),
58535 => conv_std_logic_vector(38076, 16),
58536 => conv_std_logic_vector(38304, 16),
58537 => conv_std_logic_vector(38532, 16),
58538 => conv_std_logic_vector(38760, 16),
58539 => conv_std_logic_vector(38988, 16),
58540 => conv_std_logic_vector(39216, 16),
58541 => conv_std_logic_vector(39444, 16),
58542 => conv_std_logic_vector(39672, 16),
58543 => conv_std_logic_vector(39900, 16),
58544 => conv_std_logic_vector(40128, 16),
58545 => conv_std_logic_vector(40356, 16),
58546 => conv_std_logic_vector(40584, 16),
58547 => conv_std_logic_vector(40812, 16),
58548 => conv_std_logic_vector(41040, 16),
58549 => conv_std_logic_vector(41268, 16),
58550 => conv_std_logic_vector(41496, 16),
58551 => conv_std_logic_vector(41724, 16),
58552 => conv_std_logic_vector(41952, 16),
58553 => conv_std_logic_vector(42180, 16),
58554 => conv_std_logic_vector(42408, 16),
58555 => conv_std_logic_vector(42636, 16),
58556 => conv_std_logic_vector(42864, 16),
58557 => conv_std_logic_vector(43092, 16),
58558 => conv_std_logic_vector(43320, 16),
58559 => conv_std_logic_vector(43548, 16),
58560 => conv_std_logic_vector(43776, 16),
58561 => conv_std_logic_vector(44004, 16),
58562 => conv_std_logic_vector(44232, 16),
58563 => conv_std_logic_vector(44460, 16),
58564 => conv_std_logic_vector(44688, 16),
58565 => conv_std_logic_vector(44916, 16),
58566 => conv_std_logic_vector(45144, 16),
58567 => conv_std_logic_vector(45372, 16),
58568 => conv_std_logic_vector(45600, 16),
58569 => conv_std_logic_vector(45828, 16),
58570 => conv_std_logic_vector(46056, 16),
58571 => conv_std_logic_vector(46284, 16),
58572 => conv_std_logic_vector(46512, 16),
58573 => conv_std_logic_vector(46740, 16),
58574 => conv_std_logic_vector(46968, 16),
58575 => conv_std_logic_vector(47196, 16),
58576 => conv_std_logic_vector(47424, 16),
58577 => conv_std_logic_vector(47652, 16),
58578 => conv_std_logic_vector(47880, 16),
58579 => conv_std_logic_vector(48108, 16),
58580 => conv_std_logic_vector(48336, 16),
58581 => conv_std_logic_vector(48564, 16),
58582 => conv_std_logic_vector(48792, 16),
58583 => conv_std_logic_vector(49020, 16),
58584 => conv_std_logic_vector(49248, 16),
58585 => conv_std_logic_vector(49476, 16),
58586 => conv_std_logic_vector(49704, 16),
58587 => conv_std_logic_vector(49932, 16),
58588 => conv_std_logic_vector(50160, 16),
58589 => conv_std_logic_vector(50388, 16),
58590 => conv_std_logic_vector(50616, 16),
58591 => conv_std_logic_vector(50844, 16),
58592 => conv_std_logic_vector(51072, 16),
58593 => conv_std_logic_vector(51300, 16),
58594 => conv_std_logic_vector(51528, 16),
58595 => conv_std_logic_vector(51756, 16),
58596 => conv_std_logic_vector(51984, 16),
58597 => conv_std_logic_vector(52212, 16),
58598 => conv_std_logic_vector(52440, 16),
58599 => conv_std_logic_vector(52668, 16),
58600 => conv_std_logic_vector(52896, 16),
58601 => conv_std_logic_vector(53124, 16),
58602 => conv_std_logic_vector(53352, 16),
58603 => conv_std_logic_vector(53580, 16),
58604 => conv_std_logic_vector(53808, 16),
58605 => conv_std_logic_vector(54036, 16),
58606 => conv_std_logic_vector(54264, 16),
58607 => conv_std_logic_vector(54492, 16),
58608 => conv_std_logic_vector(54720, 16),
58609 => conv_std_logic_vector(54948, 16),
58610 => conv_std_logic_vector(55176, 16),
58611 => conv_std_logic_vector(55404, 16),
58612 => conv_std_logic_vector(55632, 16),
58613 => conv_std_logic_vector(55860, 16),
58614 => conv_std_logic_vector(56088, 16),
58615 => conv_std_logic_vector(56316, 16),
58616 => conv_std_logic_vector(56544, 16),
58617 => conv_std_logic_vector(56772, 16),
58618 => conv_std_logic_vector(57000, 16),
58619 => conv_std_logic_vector(57228, 16),
58620 => conv_std_logic_vector(57456, 16),
58621 => conv_std_logic_vector(57684, 16),
58622 => conv_std_logic_vector(57912, 16),
58623 => conv_std_logic_vector(58140, 16),
58624 => conv_std_logic_vector(0, 16),
58625 => conv_std_logic_vector(229, 16),
58626 => conv_std_logic_vector(458, 16),
58627 => conv_std_logic_vector(687, 16),
58628 => conv_std_logic_vector(916, 16),
58629 => conv_std_logic_vector(1145, 16),
58630 => conv_std_logic_vector(1374, 16),
58631 => conv_std_logic_vector(1603, 16),
58632 => conv_std_logic_vector(1832, 16),
58633 => conv_std_logic_vector(2061, 16),
58634 => conv_std_logic_vector(2290, 16),
58635 => conv_std_logic_vector(2519, 16),
58636 => conv_std_logic_vector(2748, 16),
58637 => conv_std_logic_vector(2977, 16),
58638 => conv_std_logic_vector(3206, 16),
58639 => conv_std_logic_vector(3435, 16),
58640 => conv_std_logic_vector(3664, 16),
58641 => conv_std_logic_vector(3893, 16),
58642 => conv_std_logic_vector(4122, 16),
58643 => conv_std_logic_vector(4351, 16),
58644 => conv_std_logic_vector(4580, 16),
58645 => conv_std_logic_vector(4809, 16),
58646 => conv_std_logic_vector(5038, 16),
58647 => conv_std_logic_vector(5267, 16),
58648 => conv_std_logic_vector(5496, 16),
58649 => conv_std_logic_vector(5725, 16),
58650 => conv_std_logic_vector(5954, 16),
58651 => conv_std_logic_vector(6183, 16),
58652 => conv_std_logic_vector(6412, 16),
58653 => conv_std_logic_vector(6641, 16),
58654 => conv_std_logic_vector(6870, 16),
58655 => conv_std_logic_vector(7099, 16),
58656 => conv_std_logic_vector(7328, 16),
58657 => conv_std_logic_vector(7557, 16),
58658 => conv_std_logic_vector(7786, 16),
58659 => conv_std_logic_vector(8015, 16),
58660 => conv_std_logic_vector(8244, 16),
58661 => conv_std_logic_vector(8473, 16),
58662 => conv_std_logic_vector(8702, 16),
58663 => conv_std_logic_vector(8931, 16),
58664 => conv_std_logic_vector(9160, 16),
58665 => conv_std_logic_vector(9389, 16),
58666 => conv_std_logic_vector(9618, 16),
58667 => conv_std_logic_vector(9847, 16),
58668 => conv_std_logic_vector(10076, 16),
58669 => conv_std_logic_vector(10305, 16),
58670 => conv_std_logic_vector(10534, 16),
58671 => conv_std_logic_vector(10763, 16),
58672 => conv_std_logic_vector(10992, 16),
58673 => conv_std_logic_vector(11221, 16),
58674 => conv_std_logic_vector(11450, 16),
58675 => conv_std_logic_vector(11679, 16),
58676 => conv_std_logic_vector(11908, 16),
58677 => conv_std_logic_vector(12137, 16),
58678 => conv_std_logic_vector(12366, 16),
58679 => conv_std_logic_vector(12595, 16),
58680 => conv_std_logic_vector(12824, 16),
58681 => conv_std_logic_vector(13053, 16),
58682 => conv_std_logic_vector(13282, 16),
58683 => conv_std_logic_vector(13511, 16),
58684 => conv_std_logic_vector(13740, 16),
58685 => conv_std_logic_vector(13969, 16),
58686 => conv_std_logic_vector(14198, 16),
58687 => conv_std_logic_vector(14427, 16),
58688 => conv_std_logic_vector(14656, 16),
58689 => conv_std_logic_vector(14885, 16),
58690 => conv_std_logic_vector(15114, 16),
58691 => conv_std_logic_vector(15343, 16),
58692 => conv_std_logic_vector(15572, 16),
58693 => conv_std_logic_vector(15801, 16),
58694 => conv_std_logic_vector(16030, 16),
58695 => conv_std_logic_vector(16259, 16),
58696 => conv_std_logic_vector(16488, 16),
58697 => conv_std_logic_vector(16717, 16),
58698 => conv_std_logic_vector(16946, 16),
58699 => conv_std_logic_vector(17175, 16),
58700 => conv_std_logic_vector(17404, 16),
58701 => conv_std_logic_vector(17633, 16),
58702 => conv_std_logic_vector(17862, 16),
58703 => conv_std_logic_vector(18091, 16),
58704 => conv_std_logic_vector(18320, 16),
58705 => conv_std_logic_vector(18549, 16),
58706 => conv_std_logic_vector(18778, 16),
58707 => conv_std_logic_vector(19007, 16),
58708 => conv_std_logic_vector(19236, 16),
58709 => conv_std_logic_vector(19465, 16),
58710 => conv_std_logic_vector(19694, 16),
58711 => conv_std_logic_vector(19923, 16),
58712 => conv_std_logic_vector(20152, 16),
58713 => conv_std_logic_vector(20381, 16),
58714 => conv_std_logic_vector(20610, 16),
58715 => conv_std_logic_vector(20839, 16),
58716 => conv_std_logic_vector(21068, 16),
58717 => conv_std_logic_vector(21297, 16),
58718 => conv_std_logic_vector(21526, 16),
58719 => conv_std_logic_vector(21755, 16),
58720 => conv_std_logic_vector(21984, 16),
58721 => conv_std_logic_vector(22213, 16),
58722 => conv_std_logic_vector(22442, 16),
58723 => conv_std_logic_vector(22671, 16),
58724 => conv_std_logic_vector(22900, 16),
58725 => conv_std_logic_vector(23129, 16),
58726 => conv_std_logic_vector(23358, 16),
58727 => conv_std_logic_vector(23587, 16),
58728 => conv_std_logic_vector(23816, 16),
58729 => conv_std_logic_vector(24045, 16),
58730 => conv_std_logic_vector(24274, 16),
58731 => conv_std_logic_vector(24503, 16),
58732 => conv_std_logic_vector(24732, 16),
58733 => conv_std_logic_vector(24961, 16),
58734 => conv_std_logic_vector(25190, 16),
58735 => conv_std_logic_vector(25419, 16),
58736 => conv_std_logic_vector(25648, 16),
58737 => conv_std_logic_vector(25877, 16),
58738 => conv_std_logic_vector(26106, 16),
58739 => conv_std_logic_vector(26335, 16),
58740 => conv_std_logic_vector(26564, 16),
58741 => conv_std_logic_vector(26793, 16),
58742 => conv_std_logic_vector(27022, 16),
58743 => conv_std_logic_vector(27251, 16),
58744 => conv_std_logic_vector(27480, 16),
58745 => conv_std_logic_vector(27709, 16),
58746 => conv_std_logic_vector(27938, 16),
58747 => conv_std_logic_vector(28167, 16),
58748 => conv_std_logic_vector(28396, 16),
58749 => conv_std_logic_vector(28625, 16),
58750 => conv_std_logic_vector(28854, 16),
58751 => conv_std_logic_vector(29083, 16),
58752 => conv_std_logic_vector(29312, 16),
58753 => conv_std_logic_vector(29541, 16),
58754 => conv_std_logic_vector(29770, 16),
58755 => conv_std_logic_vector(29999, 16),
58756 => conv_std_logic_vector(30228, 16),
58757 => conv_std_logic_vector(30457, 16),
58758 => conv_std_logic_vector(30686, 16),
58759 => conv_std_logic_vector(30915, 16),
58760 => conv_std_logic_vector(31144, 16),
58761 => conv_std_logic_vector(31373, 16),
58762 => conv_std_logic_vector(31602, 16),
58763 => conv_std_logic_vector(31831, 16),
58764 => conv_std_logic_vector(32060, 16),
58765 => conv_std_logic_vector(32289, 16),
58766 => conv_std_logic_vector(32518, 16),
58767 => conv_std_logic_vector(32747, 16),
58768 => conv_std_logic_vector(32976, 16),
58769 => conv_std_logic_vector(33205, 16),
58770 => conv_std_logic_vector(33434, 16),
58771 => conv_std_logic_vector(33663, 16),
58772 => conv_std_logic_vector(33892, 16),
58773 => conv_std_logic_vector(34121, 16),
58774 => conv_std_logic_vector(34350, 16),
58775 => conv_std_logic_vector(34579, 16),
58776 => conv_std_logic_vector(34808, 16),
58777 => conv_std_logic_vector(35037, 16),
58778 => conv_std_logic_vector(35266, 16),
58779 => conv_std_logic_vector(35495, 16),
58780 => conv_std_logic_vector(35724, 16),
58781 => conv_std_logic_vector(35953, 16),
58782 => conv_std_logic_vector(36182, 16),
58783 => conv_std_logic_vector(36411, 16),
58784 => conv_std_logic_vector(36640, 16),
58785 => conv_std_logic_vector(36869, 16),
58786 => conv_std_logic_vector(37098, 16),
58787 => conv_std_logic_vector(37327, 16),
58788 => conv_std_logic_vector(37556, 16),
58789 => conv_std_logic_vector(37785, 16),
58790 => conv_std_logic_vector(38014, 16),
58791 => conv_std_logic_vector(38243, 16),
58792 => conv_std_logic_vector(38472, 16),
58793 => conv_std_logic_vector(38701, 16),
58794 => conv_std_logic_vector(38930, 16),
58795 => conv_std_logic_vector(39159, 16),
58796 => conv_std_logic_vector(39388, 16),
58797 => conv_std_logic_vector(39617, 16),
58798 => conv_std_logic_vector(39846, 16),
58799 => conv_std_logic_vector(40075, 16),
58800 => conv_std_logic_vector(40304, 16),
58801 => conv_std_logic_vector(40533, 16),
58802 => conv_std_logic_vector(40762, 16),
58803 => conv_std_logic_vector(40991, 16),
58804 => conv_std_logic_vector(41220, 16),
58805 => conv_std_logic_vector(41449, 16),
58806 => conv_std_logic_vector(41678, 16),
58807 => conv_std_logic_vector(41907, 16),
58808 => conv_std_logic_vector(42136, 16),
58809 => conv_std_logic_vector(42365, 16),
58810 => conv_std_logic_vector(42594, 16),
58811 => conv_std_logic_vector(42823, 16),
58812 => conv_std_logic_vector(43052, 16),
58813 => conv_std_logic_vector(43281, 16),
58814 => conv_std_logic_vector(43510, 16),
58815 => conv_std_logic_vector(43739, 16),
58816 => conv_std_logic_vector(43968, 16),
58817 => conv_std_logic_vector(44197, 16),
58818 => conv_std_logic_vector(44426, 16),
58819 => conv_std_logic_vector(44655, 16),
58820 => conv_std_logic_vector(44884, 16),
58821 => conv_std_logic_vector(45113, 16),
58822 => conv_std_logic_vector(45342, 16),
58823 => conv_std_logic_vector(45571, 16),
58824 => conv_std_logic_vector(45800, 16),
58825 => conv_std_logic_vector(46029, 16),
58826 => conv_std_logic_vector(46258, 16),
58827 => conv_std_logic_vector(46487, 16),
58828 => conv_std_logic_vector(46716, 16),
58829 => conv_std_logic_vector(46945, 16),
58830 => conv_std_logic_vector(47174, 16),
58831 => conv_std_logic_vector(47403, 16),
58832 => conv_std_logic_vector(47632, 16),
58833 => conv_std_logic_vector(47861, 16),
58834 => conv_std_logic_vector(48090, 16),
58835 => conv_std_logic_vector(48319, 16),
58836 => conv_std_logic_vector(48548, 16),
58837 => conv_std_logic_vector(48777, 16),
58838 => conv_std_logic_vector(49006, 16),
58839 => conv_std_logic_vector(49235, 16),
58840 => conv_std_logic_vector(49464, 16),
58841 => conv_std_logic_vector(49693, 16),
58842 => conv_std_logic_vector(49922, 16),
58843 => conv_std_logic_vector(50151, 16),
58844 => conv_std_logic_vector(50380, 16),
58845 => conv_std_logic_vector(50609, 16),
58846 => conv_std_logic_vector(50838, 16),
58847 => conv_std_logic_vector(51067, 16),
58848 => conv_std_logic_vector(51296, 16),
58849 => conv_std_logic_vector(51525, 16),
58850 => conv_std_logic_vector(51754, 16),
58851 => conv_std_logic_vector(51983, 16),
58852 => conv_std_logic_vector(52212, 16),
58853 => conv_std_logic_vector(52441, 16),
58854 => conv_std_logic_vector(52670, 16),
58855 => conv_std_logic_vector(52899, 16),
58856 => conv_std_logic_vector(53128, 16),
58857 => conv_std_logic_vector(53357, 16),
58858 => conv_std_logic_vector(53586, 16),
58859 => conv_std_logic_vector(53815, 16),
58860 => conv_std_logic_vector(54044, 16),
58861 => conv_std_logic_vector(54273, 16),
58862 => conv_std_logic_vector(54502, 16),
58863 => conv_std_logic_vector(54731, 16),
58864 => conv_std_logic_vector(54960, 16),
58865 => conv_std_logic_vector(55189, 16),
58866 => conv_std_logic_vector(55418, 16),
58867 => conv_std_logic_vector(55647, 16),
58868 => conv_std_logic_vector(55876, 16),
58869 => conv_std_logic_vector(56105, 16),
58870 => conv_std_logic_vector(56334, 16),
58871 => conv_std_logic_vector(56563, 16),
58872 => conv_std_logic_vector(56792, 16),
58873 => conv_std_logic_vector(57021, 16),
58874 => conv_std_logic_vector(57250, 16),
58875 => conv_std_logic_vector(57479, 16),
58876 => conv_std_logic_vector(57708, 16),
58877 => conv_std_logic_vector(57937, 16),
58878 => conv_std_logic_vector(58166, 16),
58879 => conv_std_logic_vector(58395, 16),
58880 => conv_std_logic_vector(0, 16),
58881 => conv_std_logic_vector(230, 16),
58882 => conv_std_logic_vector(460, 16),
58883 => conv_std_logic_vector(690, 16),
58884 => conv_std_logic_vector(920, 16),
58885 => conv_std_logic_vector(1150, 16),
58886 => conv_std_logic_vector(1380, 16),
58887 => conv_std_logic_vector(1610, 16),
58888 => conv_std_logic_vector(1840, 16),
58889 => conv_std_logic_vector(2070, 16),
58890 => conv_std_logic_vector(2300, 16),
58891 => conv_std_logic_vector(2530, 16),
58892 => conv_std_logic_vector(2760, 16),
58893 => conv_std_logic_vector(2990, 16),
58894 => conv_std_logic_vector(3220, 16),
58895 => conv_std_logic_vector(3450, 16),
58896 => conv_std_logic_vector(3680, 16),
58897 => conv_std_logic_vector(3910, 16),
58898 => conv_std_logic_vector(4140, 16),
58899 => conv_std_logic_vector(4370, 16),
58900 => conv_std_logic_vector(4600, 16),
58901 => conv_std_logic_vector(4830, 16),
58902 => conv_std_logic_vector(5060, 16),
58903 => conv_std_logic_vector(5290, 16),
58904 => conv_std_logic_vector(5520, 16),
58905 => conv_std_logic_vector(5750, 16),
58906 => conv_std_logic_vector(5980, 16),
58907 => conv_std_logic_vector(6210, 16),
58908 => conv_std_logic_vector(6440, 16),
58909 => conv_std_logic_vector(6670, 16),
58910 => conv_std_logic_vector(6900, 16),
58911 => conv_std_logic_vector(7130, 16),
58912 => conv_std_logic_vector(7360, 16),
58913 => conv_std_logic_vector(7590, 16),
58914 => conv_std_logic_vector(7820, 16),
58915 => conv_std_logic_vector(8050, 16),
58916 => conv_std_logic_vector(8280, 16),
58917 => conv_std_logic_vector(8510, 16),
58918 => conv_std_logic_vector(8740, 16),
58919 => conv_std_logic_vector(8970, 16),
58920 => conv_std_logic_vector(9200, 16),
58921 => conv_std_logic_vector(9430, 16),
58922 => conv_std_logic_vector(9660, 16),
58923 => conv_std_logic_vector(9890, 16),
58924 => conv_std_logic_vector(10120, 16),
58925 => conv_std_logic_vector(10350, 16),
58926 => conv_std_logic_vector(10580, 16),
58927 => conv_std_logic_vector(10810, 16),
58928 => conv_std_logic_vector(11040, 16),
58929 => conv_std_logic_vector(11270, 16),
58930 => conv_std_logic_vector(11500, 16),
58931 => conv_std_logic_vector(11730, 16),
58932 => conv_std_logic_vector(11960, 16),
58933 => conv_std_logic_vector(12190, 16),
58934 => conv_std_logic_vector(12420, 16),
58935 => conv_std_logic_vector(12650, 16),
58936 => conv_std_logic_vector(12880, 16),
58937 => conv_std_logic_vector(13110, 16),
58938 => conv_std_logic_vector(13340, 16),
58939 => conv_std_logic_vector(13570, 16),
58940 => conv_std_logic_vector(13800, 16),
58941 => conv_std_logic_vector(14030, 16),
58942 => conv_std_logic_vector(14260, 16),
58943 => conv_std_logic_vector(14490, 16),
58944 => conv_std_logic_vector(14720, 16),
58945 => conv_std_logic_vector(14950, 16),
58946 => conv_std_logic_vector(15180, 16),
58947 => conv_std_logic_vector(15410, 16),
58948 => conv_std_logic_vector(15640, 16),
58949 => conv_std_logic_vector(15870, 16),
58950 => conv_std_logic_vector(16100, 16),
58951 => conv_std_logic_vector(16330, 16),
58952 => conv_std_logic_vector(16560, 16),
58953 => conv_std_logic_vector(16790, 16),
58954 => conv_std_logic_vector(17020, 16),
58955 => conv_std_logic_vector(17250, 16),
58956 => conv_std_logic_vector(17480, 16),
58957 => conv_std_logic_vector(17710, 16),
58958 => conv_std_logic_vector(17940, 16),
58959 => conv_std_logic_vector(18170, 16),
58960 => conv_std_logic_vector(18400, 16),
58961 => conv_std_logic_vector(18630, 16),
58962 => conv_std_logic_vector(18860, 16),
58963 => conv_std_logic_vector(19090, 16),
58964 => conv_std_logic_vector(19320, 16),
58965 => conv_std_logic_vector(19550, 16),
58966 => conv_std_logic_vector(19780, 16),
58967 => conv_std_logic_vector(20010, 16),
58968 => conv_std_logic_vector(20240, 16),
58969 => conv_std_logic_vector(20470, 16),
58970 => conv_std_logic_vector(20700, 16),
58971 => conv_std_logic_vector(20930, 16),
58972 => conv_std_logic_vector(21160, 16),
58973 => conv_std_logic_vector(21390, 16),
58974 => conv_std_logic_vector(21620, 16),
58975 => conv_std_logic_vector(21850, 16),
58976 => conv_std_logic_vector(22080, 16),
58977 => conv_std_logic_vector(22310, 16),
58978 => conv_std_logic_vector(22540, 16),
58979 => conv_std_logic_vector(22770, 16),
58980 => conv_std_logic_vector(23000, 16),
58981 => conv_std_logic_vector(23230, 16),
58982 => conv_std_logic_vector(23460, 16),
58983 => conv_std_logic_vector(23690, 16),
58984 => conv_std_logic_vector(23920, 16),
58985 => conv_std_logic_vector(24150, 16),
58986 => conv_std_logic_vector(24380, 16),
58987 => conv_std_logic_vector(24610, 16),
58988 => conv_std_logic_vector(24840, 16),
58989 => conv_std_logic_vector(25070, 16),
58990 => conv_std_logic_vector(25300, 16),
58991 => conv_std_logic_vector(25530, 16),
58992 => conv_std_logic_vector(25760, 16),
58993 => conv_std_logic_vector(25990, 16),
58994 => conv_std_logic_vector(26220, 16),
58995 => conv_std_logic_vector(26450, 16),
58996 => conv_std_logic_vector(26680, 16),
58997 => conv_std_logic_vector(26910, 16),
58998 => conv_std_logic_vector(27140, 16),
58999 => conv_std_logic_vector(27370, 16),
59000 => conv_std_logic_vector(27600, 16),
59001 => conv_std_logic_vector(27830, 16),
59002 => conv_std_logic_vector(28060, 16),
59003 => conv_std_logic_vector(28290, 16),
59004 => conv_std_logic_vector(28520, 16),
59005 => conv_std_logic_vector(28750, 16),
59006 => conv_std_logic_vector(28980, 16),
59007 => conv_std_logic_vector(29210, 16),
59008 => conv_std_logic_vector(29440, 16),
59009 => conv_std_logic_vector(29670, 16),
59010 => conv_std_logic_vector(29900, 16),
59011 => conv_std_logic_vector(30130, 16),
59012 => conv_std_logic_vector(30360, 16),
59013 => conv_std_logic_vector(30590, 16),
59014 => conv_std_logic_vector(30820, 16),
59015 => conv_std_logic_vector(31050, 16),
59016 => conv_std_logic_vector(31280, 16),
59017 => conv_std_logic_vector(31510, 16),
59018 => conv_std_logic_vector(31740, 16),
59019 => conv_std_logic_vector(31970, 16),
59020 => conv_std_logic_vector(32200, 16),
59021 => conv_std_logic_vector(32430, 16),
59022 => conv_std_logic_vector(32660, 16),
59023 => conv_std_logic_vector(32890, 16),
59024 => conv_std_logic_vector(33120, 16),
59025 => conv_std_logic_vector(33350, 16),
59026 => conv_std_logic_vector(33580, 16),
59027 => conv_std_logic_vector(33810, 16),
59028 => conv_std_logic_vector(34040, 16),
59029 => conv_std_logic_vector(34270, 16),
59030 => conv_std_logic_vector(34500, 16),
59031 => conv_std_logic_vector(34730, 16),
59032 => conv_std_logic_vector(34960, 16),
59033 => conv_std_logic_vector(35190, 16),
59034 => conv_std_logic_vector(35420, 16),
59035 => conv_std_logic_vector(35650, 16),
59036 => conv_std_logic_vector(35880, 16),
59037 => conv_std_logic_vector(36110, 16),
59038 => conv_std_logic_vector(36340, 16),
59039 => conv_std_logic_vector(36570, 16),
59040 => conv_std_logic_vector(36800, 16),
59041 => conv_std_logic_vector(37030, 16),
59042 => conv_std_logic_vector(37260, 16),
59043 => conv_std_logic_vector(37490, 16),
59044 => conv_std_logic_vector(37720, 16),
59045 => conv_std_logic_vector(37950, 16),
59046 => conv_std_logic_vector(38180, 16),
59047 => conv_std_logic_vector(38410, 16),
59048 => conv_std_logic_vector(38640, 16),
59049 => conv_std_logic_vector(38870, 16),
59050 => conv_std_logic_vector(39100, 16),
59051 => conv_std_logic_vector(39330, 16),
59052 => conv_std_logic_vector(39560, 16),
59053 => conv_std_logic_vector(39790, 16),
59054 => conv_std_logic_vector(40020, 16),
59055 => conv_std_logic_vector(40250, 16),
59056 => conv_std_logic_vector(40480, 16),
59057 => conv_std_logic_vector(40710, 16),
59058 => conv_std_logic_vector(40940, 16),
59059 => conv_std_logic_vector(41170, 16),
59060 => conv_std_logic_vector(41400, 16),
59061 => conv_std_logic_vector(41630, 16),
59062 => conv_std_logic_vector(41860, 16),
59063 => conv_std_logic_vector(42090, 16),
59064 => conv_std_logic_vector(42320, 16),
59065 => conv_std_logic_vector(42550, 16),
59066 => conv_std_logic_vector(42780, 16),
59067 => conv_std_logic_vector(43010, 16),
59068 => conv_std_logic_vector(43240, 16),
59069 => conv_std_logic_vector(43470, 16),
59070 => conv_std_logic_vector(43700, 16),
59071 => conv_std_logic_vector(43930, 16),
59072 => conv_std_logic_vector(44160, 16),
59073 => conv_std_logic_vector(44390, 16),
59074 => conv_std_logic_vector(44620, 16),
59075 => conv_std_logic_vector(44850, 16),
59076 => conv_std_logic_vector(45080, 16),
59077 => conv_std_logic_vector(45310, 16),
59078 => conv_std_logic_vector(45540, 16),
59079 => conv_std_logic_vector(45770, 16),
59080 => conv_std_logic_vector(46000, 16),
59081 => conv_std_logic_vector(46230, 16),
59082 => conv_std_logic_vector(46460, 16),
59083 => conv_std_logic_vector(46690, 16),
59084 => conv_std_logic_vector(46920, 16),
59085 => conv_std_logic_vector(47150, 16),
59086 => conv_std_logic_vector(47380, 16),
59087 => conv_std_logic_vector(47610, 16),
59088 => conv_std_logic_vector(47840, 16),
59089 => conv_std_logic_vector(48070, 16),
59090 => conv_std_logic_vector(48300, 16),
59091 => conv_std_logic_vector(48530, 16),
59092 => conv_std_logic_vector(48760, 16),
59093 => conv_std_logic_vector(48990, 16),
59094 => conv_std_logic_vector(49220, 16),
59095 => conv_std_logic_vector(49450, 16),
59096 => conv_std_logic_vector(49680, 16),
59097 => conv_std_logic_vector(49910, 16),
59098 => conv_std_logic_vector(50140, 16),
59099 => conv_std_logic_vector(50370, 16),
59100 => conv_std_logic_vector(50600, 16),
59101 => conv_std_logic_vector(50830, 16),
59102 => conv_std_logic_vector(51060, 16),
59103 => conv_std_logic_vector(51290, 16),
59104 => conv_std_logic_vector(51520, 16),
59105 => conv_std_logic_vector(51750, 16),
59106 => conv_std_logic_vector(51980, 16),
59107 => conv_std_logic_vector(52210, 16),
59108 => conv_std_logic_vector(52440, 16),
59109 => conv_std_logic_vector(52670, 16),
59110 => conv_std_logic_vector(52900, 16),
59111 => conv_std_logic_vector(53130, 16),
59112 => conv_std_logic_vector(53360, 16),
59113 => conv_std_logic_vector(53590, 16),
59114 => conv_std_logic_vector(53820, 16),
59115 => conv_std_logic_vector(54050, 16),
59116 => conv_std_logic_vector(54280, 16),
59117 => conv_std_logic_vector(54510, 16),
59118 => conv_std_logic_vector(54740, 16),
59119 => conv_std_logic_vector(54970, 16),
59120 => conv_std_logic_vector(55200, 16),
59121 => conv_std_logic_vector(55430, 16),
59122 => conv_std_logic_vector(55660, 16),
59123 => conv_std_logic_vector(55890, 16),
59124 => conv_std_logic_vector(56120, 16),
59125 => conv_std_logic_vector(56350, 16),
59126 => conv_std_logic_vector(56580, 16),
59127 => conv_std_logic_vector(56810, 16),
59128 => conv_std_logic_vector(57040, 16),
59129 => conv_std_logic_vector(57270, 16),
59130 => conv_std_logic_vector(57500, 16),
59131 => conv_std_logic_vector(57730, 16),
59132 => conv_std_logic_vector(57960, 16),
59133 => conv_std_logic_vector(58190, 16),
59134 => conv_std_logic_vector(58420, 16),
59135 => conv_std_logic_vector(58650, 16),
59136 => conv_std_logic_vector(0, 16),
59137 => conv_std_logic_vector(231, 16),
59138 => conv_std_logic_vector(462, 16),
59139 => conv_std_logic_vector(693, 16),
59140 => conv_std_logic_vector(924, 16),
59141 => conv_std_logic_vector(1155, 16),
59142 => conv_std_logic_vector(1386, 16),
59143 => conv_std_logic_vector(1617, 16),
59144 => conv_std_logic_vector(1848, 16),
59145 => conv_std_logic_vector(2079, 16),
59146 => conv_std_logic_vector(2310, 16),
59147 => conv_std_logic_vector(2541, 16),
59148 => conv_std_logic_vector(2772, 16),
59149 => conv_std_logic_vector(3003, 16),
59150 => conv_std_logic_vector(3234, 16),
59151 => conv_std_logic_vector(3465, 16),
59152 => conv_std_logic_vector(3696, 16),
59153 => conv_std_logic_vector(3927, 16),
59154 => conv_std_logic_vector(4158, 16),
59155 => conv_std_logic_vector(4389, 16),
59156 => conv_std_logic_vector(4620, 16),
59157 => conv_std_logic_vector(4851, 16),
59158 => conv_std_logic_vector(5082, 16),
59159 => conv_std_logic_vector(5313, 16),
59160 => conv_std_logic_vector(5544, 16),
59161 => conv_std_logic_vector(5775, 16),
59162 => conv_std_logic_vector(6006, 16),
59163 => conv_std_logic_vector(6237, 16),
59164 => conv_std_logic_vector(6468, 16),
59165 => conv_std_logic_vector(6699, 16),
59166 => conv_std_logic_vector(6930, 16),
59167 => conv_std_logic_vector(7161, 16),
59168 => conv_std_logic_vector(7392, 16),
59169 => conv_std_logic_vector(7623, 16),
59170 => conv_std_logic_vector(7854, 16),
59171 => conv_std_logic_vector(8085, 16),
59172 => conv_std_logic_vector(8316, 16),
59173 => conv_std_logic_vector(8547, 16),
59174 => conv_std_logic_vector(8778, 16),
59175 => conv_std_logic_vector(9009, 16),
59176 => conv_std_logic_vector(9240, 16),
59177 => conv_std_logic_vector(9471, 16),
59178 => conv_std_logic_vector(9702, 16),
59179 => conv_std_logic_vector(9933, 16),
59180 => conv_std_logic_vector(10164, 16),
59181 => conv_std_logic_vector(10395, 16),
59182 => conv_std_logic_vector(10626, 16),
59183 => conv_std_logic_vector(10857, 16),
59184 => conv_std_logic_vector(11088, 16),
59185 => conv_std_logic_vector(11319, 16),
59186 => conv_std_logic_vector(11550, 16),
59187 => conv_std_logic_vector(11781, 16),
59188 => conv_std_logic_vector(12012, 16),
59189 => conv_std_logic_vector(12243, 16),
59190 => conv_std_logic_vector(12474, 16),
59191 => conv_std_logic_vector(12705, 16),
59192 => conv_std_logic_vector(12936, 16),
59193 => conv_std_logic_vector(13167, 16),
59194 => conv_std_logic_vector(13398, 16),
59195 => conv_std_logic_vector(13629, 16),
59196 => conv_std_logic_vector(13860, 16),
59197 => conv_std_logic_vector(14091, 16),
59198 => conv_std_logic_vector(14322, 16),
59199 => conv_std_logic_vector(14553, 16),
59200 => conv_std_logic_vector(14784, 16),
59201 => conv_std_logic_vector(15015, 16),
59202 => conv_std_logic_vector(15246, 16),
59203 => conv_std_logic_vector(15477, 16),
59204 => conv_std_logic_vector(15708, 16),
59205 => conv_std_logic_vector(15939, 16),
59206 => conv_std_logic_vector(16170, 16),
59207 => conv_std_logic_vector(16401, 16),
59208 => conv_std_logic_vector(16632, 16),
59209 => conv_std_logic_vector(16863, 16),
59210 => conv_std_logic_vector(17094, 16),
59211 => conv_std_logic_vector(17325, 16),
59212 => conv_std_logic_vector(17556, 16),
59213 => conv_std_logic_vector(17787, 16),
59214 => conv_std_logic_vector(18018, 16),
59215 => conv_std_logic_vector(18249, 16),
59216 => conv_std_logic_vector(18480, 16),
59217 => conv_std_logic_vector(18711, 16),
59218 => conv_std_logic_vector(18942, 16),
59219 => conv_std_logic_vector(19173, 16),
59220 => conv_std_logic_vector(19404, 16),
59221 => conv_std_logic_vector(19635, 16),
59222 => conv_std_logic_vector(19866, 16),
59223 => conv_std_logic_vector(20097, 16),
59224 => conv_std_logic_vector(20328, 16),
59225 => conv_std_logic_vector(20559, 16),
59226 => conv_std_logic_vector(20790, 16),
59227 => conv_std_logic_vector(21021, 16),
59228 => conv_std_logic_vector(21252, 16),
59229 => conv_std_logic_vector(21483, 16),
59230 => conv_std_logic_vector(21714, 16),
59231 => conv_std_logic_vector(21945, 16),
59232 => conv_std_logic_vector(22176, 16),
59233 => conv_std_logic_vector(22407, 16),
59234 => conv_std_logic_vector(22638, 16),
59235 => conv_std_logic_vector(22869, 16),
59236 => conv_std_logic_vector(23100, 16),
59237 => conv_std_logic_vector(23331, 16),
59238 => conv_std_logic_vector(23562, 16),
59239 => conv_std_logic_vector(23793, 16),
59240 => conv_std_logic_vector(24024, 16),
59241 => conv_std_logic_vector(24255, 16),
59242 => conv_std_logic_vector(24486, 16),
59243 => conv_std_logic_vector(24717, 16),
59244 => conv_std_logic_vector(24948, 16),
59245 => conv_std_logic_vector(25179, 16),
59246 => conv_std_logic_vector(25410, 16),
59247 => conv_std_logic_vector(25641, 16),
59248 => conv_std_logic_vector(25872, 16),
59249 => conv_std_logic_vector(26103, 16),
59250 => conv_std_logic_vector(26334, 16),
59251 => conv_std_logic_vector(26565, 16),
59252 => conv_std_logic_vector(26796, 16),
59253 => conv_std_logic_vector(27027, 16),
59254 => conv_std_logic_vector(27258, 16),
59255 => conv_std_logic_vector(27489, 16),
59256 => conv_std_logic_vector(27720, 16),
59257 => conv_std_logic_vector(27951, 16),
59258 => conv_std_logic_vector(28182, 16),
59259 => conv_std_logic_vector(28413, 16),
59260 => conv_std_logic_vector(28644, 16),
59261 => conv_std_logic_vector(28875, 16),
59262 => conv_std_logic_vector(29106, 16),
59263 => conv_std_logic_vector(29337, 16),
59264 => conv_std_logic_vector(29568, 16),
59265 => conv_std_logic_vector(29799, 16),
59266 => conv_std_logic_vector(30030, 16),
59267 => conv_std_logic_vector(30261, 16),
59268 => conv_std_logic_vector(30492, 16),
59269 => conv_std_logic_vector(30723, 16),
59270 => conv_std_logic_vector(30954, 16),
59271 => conv_std_logic_vector(31185, 16),
59272 => conv_std_logic_vector(31416, 16),
59273 => conv_std_logic_vector(31647, 16),
59274 => conv_std_logic_vector(31878, 16),
59275 => conv_std_logic_vector(32109, 16),
59276 => conv_std_logic_vector(32340, 16),
59277 => conv_std_logic_vector(32571, 16),
59278 => conv_std_logic_vector(32802, 16),
59279 => conv_std_logic_vector(33033, 16),
59280 => conv_std_logic_vector(33264, 16),
59281 => conv_std_logic_vector(33495, 16),
59282 => conv_std_logic_vector(33726, 16),
59283 => conv_std_logic_vector(33957, 16),
59284 => conv_std_logic_vector(34188, 16),
59285 => conv_std_logic_vector(34419, 16),
59286 => conv_std_logic_vector(34650, 16),
59287 => conv_std_logic_vector(34881, 16),
59288 => conv_std_logic_vector(35112, 16),
59289 => conv_std_logic_vector(35343, 16),
59290 => conv_std_logic_vector(35574, 16),
59291 => conv_std_logic_vector(35805, 16),
59292 => conv_std_logic_vector(36036, 16),
59293 => conv_std_logic_vector(36267, 16),
59294 => conv_std_logic_vector(36498, 16),
59295 => conv_std_logic_vector(36729, 16),
59296 => conv_std_logic_vector(36960, 16),
59297 => conv_std_logic_vector(37191, 16),
59298 => conv_std_logic_vector(37422, 16),
59299 => conv_std_logic_vector(37653, 16),
59300 => conv_std_logic_vector(37884, 16),
59301 => conv_std_logic_vector(38115, 16),
59302 => conv_std_logic_vector(38346, 16),
59303 => conv_std_logic_vector(38577, 16),
59304 => conv_std_logic_vector(38808, 16),
59305 => conv_std_logic_vector(39039, 16),
59306 => conv_std_logic_vector(39270, 16),
59307 => conv_std_logic_vector(39501, 16),
59308 => conv_std_logic_vector(39732, 16),
59309 => conv_std_logic_vector(39963, 16),
59310 => conv_std_logic_vector(40194, 16),
59311 => conv_std_logic_vector(40425, 16),
59312 => conv_std_logic_vector(40656, 16),
59313 => conv_std_logic_vector(40887, 16),
59314 => conv_std_logic_vector(41118, 16),
59315 => conv_std_logic_vector(41349, 16),
59316 => conv_std_logic_vector(41580, 16),
59317 => conv_std_logic_vector(41811, 16),
59318 => conv_std_logic_vector(42042, 16),
59319 => conv_std_logic_vector(42273, 16),
59320 => conv_std_logic_vector(42504, 16),
59321 => conv_std_logic_vector(42735, 16),
59322 => conv_std_logic_vector(42966, 16),
59323 => conv_std_logic_vector(43197, 16),
59324 => conv_std_logic_vector(43428, 16),
59325 => conv_std_logic_vector(43659, 16),
59326 => conv_std_logic_vector(43890, 16),
59327 => conv_std_logic_vector(44121, 16),
59328 => conv_std_logic_vector(44352, 16),
59329 => conv_std_logic_vector(44583, 16),
59330 => conv_std_logic_vector(44814, 16),
59331 => conv_std_logic_vector(45045, 16),
59332 => conv_std_logic_vector(45276, 16),
59333 => conv_std_logic_vector(45507, 16),
59334 => conv_std_logic_vector(45738, 16),
59335 => conv_std_logic_vector(45969, 16),
59336 => conv_std_logic_vector(46200, 16),
59337 => conv_std_logic_vector(46431, 16),
59338 => conv_std_logic_vector(46662, 16),
59339 => conv_std_logic_vector(46893, 16),
59340 => conv_std_logic_vector(47124, 16),
59341 => conv_std_logic_vector(47355, 16),
59342 => conv_std_logic_vector(47586, 16),
59343 => conv_std_logic_vector(47817, 16),
59344 => conv_std_logic_vector(48048, 16),
59345 => conv_std_logic_vector(48279, 16),
59346 => conv_std_logic_vector(48510, 16),
59347 => conv_std_logic_vector(48741, 16),
59348 => conv_std_logic_vector(48972, 16),
59349 => conv_std_logic_vector(49203, 16),
59350 => conv_std_logic_vector(49434, 16),
59351 => conv_std_logic_vector(49665, 16),
59352 => conv_std_logic_vector(49896, 16),
59353 => conv_std_logic_vector(50127, 16),
59354 => conv_std_logic_vector(50358, 16),
59355 => conv_std_logic_vector(50589, 16),
59356 => conv_std_logic_vector(50820, 16),
59357 => conv_std_logic_vector(51051, 16),
59358 => conv_std_logic_vector(51282, 16),
59359 => conv_std_logic_vector(51513, 16),
59360 => conv_std_logic_vector(51744, 16),
59361 => conv_std_logic_vector(51975, 16),
59362 => conv_std_logic_vector(52206, 16),
59363 => conv_std_logic_vector(52437, 16),
59364 => conv_std_logic_vector(52668, 16),
59365 => conv_std_logic_vector(52899, 16),
59366 => conv_std_logic_vector(53130, 16),
59367 => conv_std_logic_vector(53361, 16),
59368 => conv_std_logic_vector(53592, 16),
59369 => conv_std_logic_vector(53823, 16),
59370 => conv_std_logic_vector(54054, 16),
59371 => conv_std_logic_vector(54285, 16),
59372 => conv_std_logic_vector(54516, 16),
59373 => conv_std_logic_vector(54747, 16),
59374 => conv_std_logic_vector(54978, 16),
59375 => conv_std_logic_vector(55209, 16),
59376 => conv_std_logic_vector(55440, 16),
59377 => conv_std_logic_vector(55671, 16),
59378 => conv_std_logic_vector(55902, 16),
59379 => conv_std_logic_vector(56133, 16),
59380 => conv_std_logic_vector(56364, 16),
59381 => conv_std_logic_vector(56595, 16),
59382 => conv_std_logic_vector(56826, 16),
59383 => conv_std_logic_vector(57057, 16),
59384 => conv_std_logic_vector(57288, 16),
59385 => conv_std_logic_vector(57519, 16),
59386 => conv_std_logic_vector(57750, 16),
59387 => conv_std_logic_vector(57981, 16),
59388 => conv_std_logic_vector(58212, 16),
59389 => conv_std_logic_vector(58443, 16),
59390 => conv_std_logic_vector(58674, 16),
59391 => conv_std_logic_vector(58905, 16),
59392 => conv_std_logic_vector(0, 16),
59393 => conv_std_logic_vector(232, 16),
59394 => conv_std_logic_vector(464, 16),
59395 => conv_std_logic_vector(696, 16),
59396 => conv_std_logic_vector(928, 16),
59397 => conv_std_logic_vector(1160, 16),
59398 => conv_std_logic_vector(1392, 16),
59399 => conv_std_logic_vector(1624, 16),
59400 => conv_std_logic_vector(1856, 16),
59401 => conv_std_logic_vector(2088, 16),
59402 => conv_std_logic_vector(2320, 16),
59403 => conv_std_logic_vector(2552, 16),
59404 => conv_std_logic_vector(2784, 16),
59405 => conv_std_logic_vector(3016, 16),
59406 => conv_std_logic_vector(3248, 16),
59407 => conv_std_logic_vector(3480, 16),
59408 => conv_std_logic_vector(3712, 16),
59409 => conv_std_logic_vector(3944, 16),
59410 => conv_std_logic_vector(4176, 16),
59411 => conv_std_logic_vector(4408, 16),
59412 => conv_std_logic_vector(4640, 16),
59413 => conv_std_logic_vector(4872, 16),
59414 => conv_std_logic_vector(5104, 16),
59415 => conv_std_logic_vector(5336, 16),
59416 => conv_std_logic_vector(5568, 16),
59417 => conv_std_logic_vector(5800, 16),
59418 => conv_std_logic_vector(6032, 16),
59419 => conv_std_logic_vector(6264, 16),
59420 => conv_std_logic_vector(6496, 16),
59421 => conv_std_logic_vector(6728, 16),
59422 => conv_std_logic_vector(6960, 16),
59423 => conv_std_logic_vector(7192, 16),
59424 => conv_std_logic_vector(7424, 16),
59425 => conv_std_logic_vector(7656, 16),
59426 => conv_std_logic_vector(7888, 16),
59427 => conv_std_logic_vector(8120, 16),
59428 => conv_std_logic_vector(8352, 16),
59429 => conv_std_logic_vector(8584, 16),
59430 => conv_std_logic_vector(8816, 16),
59431 => conv_std_logic_vector(9048, 16),
59432 => conv_std_logic_vector(9280, 16),
59433 => conv_std_logic_vector(9512, 16),
59434 => conv_std_logic_vector(9744, 16),
59435 => conv_std_logic_vector(9976, 16),
59436 => conv_std_logic_vector(10208, 16),
59437 => conv_std_logic_vector(10440, 16),
59438 => conv_std_logic_vector(10672, 16),
59439 => conv_std_logic_vector(10904, 16),
59440 => conv_std_logic_vector(11136, 16),
59441 => conv_std_logic_vector(11368, 16),
59442 => conv_std_logic_vector(11600, 16),
59443 => conv_std_logic_vector(11832, 16),
59444 => conv_std_logic_vector(12064, 16),
59445 => conv_std_logic_vector(12296, 16),
59446 => conv_std_logic_vector(12528, 16),
59447 => conv_std_logic_vector(12760, 16),
59448 => conv_std_logic_vector(12992, 16),
59449 => conv_std_logic_vector(13224, 16),
59450 => conv_std_logic_vector(13456, 16),
59451 => conv_std_logic_vector(13688, 16),
59452 => conv_std_logic_vector(13920, 16),
59453 => conv_std_logic_vector(14152, 16),
59454 => conv_std_logic_vector(14384, 16),
59455 => conv_std_logic_vector(14616, 16),
59456 => conv_std_logic_vector(14848, 16),
59457 => conv_std_logic_vector(15080, 16),
59458 => conv_std_logic_vector(15312, 16),
59459 => conv_std_logic_vector(15544, 16),
59460 => conv_std_logic_vector(15776, 16),
59461 => conv_std_logic_vector(16008, 16),
59462 => conv_std_logic_vector(16240, 16),
59463 => conv_std_logic_vector(16472, 16),
59464 => conv_std_logic_vector(16704, 16),
59465 => conv_std_logic_vector(16936, 16),
59466 => conv_std_logic_vector(17168, 16),
59467 => conv_std_logic_vector(17400, 16),
59468 => conv_std_logic_vector(17632, 16),
59469 => conv_std_logic_vector(17864, 16),
59470 => conv_std_logic_vector(18096, 16),
59471 => conv_std_logic_vector(18328, 16),
59472 => conv_std_logic_vector(18560, 16),
59473 => conv_std_logic_vector(18792, 16),
59474 => conv_std_logic_vector(19024, 16),
59475 => conv_std_logic_vector(19256, 16),
59476 => conv_std_logic_vector(19488, 16),
59477 => conv_std_logic_vector(19720, 16),
59478 => conv_std_logic_vector(19952, 16),
59479 => conv_std_logic_vector(20184, 16),
59480 => conv_std_logic_vector(20416, 16),
59481 => conv_std_logic_vector(20648, 16),
59482 => conv_std_logic_vector(20880, 16),
59483 => conv_std_logic_vector(21112, 16),
59484 => conv_std_logic_vector(21344, 16),
59485 => conv_std_logic_vector(21576, 16),
59486 => conv_std_logic_vector(21808, 16),
59487 => conv_std_logic_vector(22040, 16),
59488 => conv_std_logic_vector(22272, 16),
59489 => conv_std_logic_vector(22504, 16),
59490 => conv_std_logic_vector(22736, 16),
59491 => conv_std_logic_vector(22968, 16),
59492 => conv_std_logic_vector(23200, 16),
59493 => conv_std_logic_vector(23432, 16),
59494 => conv_std_logic_vector(23664, 16),
59495 => conv_std_logic_vector(23896, 16),
59496 => conv_std_logic_vector(24128, 16),
59497 => conv_std_logic_vector(24360, 16),
59498 => conv_std_logic_vector(24592, 16),
59499 => conv_std_logic_vector(24824, 16),
59500 => conv_std_logic_vector(25056, 16),
59501 => conv_std_logic_vector(25288, 16),
59502 => conv_std_logic_vector(25520, 16),
59503 => conv_std_logic_vector(25752, 16),
59504 => conv_std_logic_vector(25984, 16),
59505 => conv_std_logic_vector(26216, 16),
59506 => conv_std_logic_vector(26448, 16),
59507 => conv_std_logic_vector(26680, 16),
59508 => conv_std_logic_vector(26912, 16),
59509 => conv_std_logic_vector(27144, 16),
59510 => conv_std_logic_vector(27376, 16),
59511 => conv_std_logic_vector(27608, 16),
59512 => conv_std_logic_vector(27840, 16),
59513 => conv_std_logic_vector(28072, 16),
59514 => conv_std_logic_vector(28304, 16),
59515 => conv_std_logic_vector(28536, 16),
59516 => conv_std_logic_vector(28768, 16),
59517 => conv_std_logic_vector(29000, 16),
59518 => conv_std_logic_vector(29232, 16),
59519 => conv_std_logic_vector(29464, 16),
59520 => conv_std_logic_vector(29696, 16),
59521 => conv_std_logic_vector(29928, 16),
59522 => conv_std_logic_vector(30160, 16),
59523 => conv_std_logic_vector(30392, 16),
59524 => conv_std_logic_vector(30624, 16),
59525 => conv_std_logic_vector(30856, 16),
59526 => conv_std_logic_vector(31088, 16),
59527 => conv_std_logic_vector(31320, 16),
59528 => conv_std_logic_vector(31552, 16),
59529 => conv_std_logic_vector(31784, 16),
59530 => conv_std_logic_vector(32016, 16),
59531 => conv_std_logic_vector(32248, 16),
59532 => conv_std_logic_vector(32480, 16),
59533 => conv_std_logic_vector(32712, 16),
59534 => conv_std_logic_vector(32944, 16),
59535 => conv_std_logic_vector(33176, 16),
59536 => conv_std_logic_vector(33408, 16),
59537 => conv_std_logic_vector(33640, 16),
59538 => conv_std_logic_vector(33872, 16),
59539 => conv_std_logic_vector(34104, 16),
59540 => conv_std_logic_vector(34336, 16),
59541 => conv_std_logic_vector(34568, 16),
59542 => conv_std_logic_vector(34800, 16),
59543 => conv_std_logic_vector(35032, 16),
59544 => conv_std_logic_vector(35264, 16),
59545 => conv_std_logic_vector(35496, 16),
59546 => conv_std_logic_vector(35728, 16),
59547 => conv_std_logic_vector(35960, 16),
59548 => conv_std_logic_vector(36192, 16),
59549 => conv_std_logic_vector(36424, 16),
59550 => conv_std_logic_vector(36656, 16),
59551 => conv_std_logic_vector(36888, 16),
59552 => conv_std_logic_vector(37120, 16),
59553 => conv_std_logic_vector(37352, 16),
59554 => conv_std_logic_vector(37584, 16),
59555 => conv_std_logic_vector(37816, 16),
59556 => conv_std_logic_vector(38048, 16),
59557 => conv_std_logic_vector(38280, 16),
59558 => conv_std_logic_vector(38512, 16),
59559 => conv_std_logic_vector(38744, 16),
59560 => conv_std_logic_vector(38976, 16),
59561 => conv_std_logic_vector(39208, 16),
59562 => conv_std_logic_vector(39440, 16),
59563 => conv_std_logic_vector(39672, 16),
59564 => conv_std_logic_vector(39904, 16),
59565 => conv_std_logic_vector(40136, 16),
59566 => conv_std_logic_vector(40368, 16),
59567 => conv_std_logic_vector(40600, 16),
59568 => conv_std_logic_vector(40832, 16),
59569 => conv_std_logic_vector(41064, 16),
59570 => conv_std_logic_vector(41296, 16),
59571 => conv_std_logic_vector(41528, 16),
59572 => conv_std_logic_vector(41760, 16),
59573 => conv_std_logic_vector(41992, 16),
59574 => conv_std_logic_vector(42224, 16),
59575 => conv_std_logic_vector(42456, 16),
59576 => conv_std_logic_vector(42688, 16),
59577 => conv_std_logic_vector(42920, 16),
59578 => conv_std_logic_vector(43152, 16),
59579 => conv_std_logic_vector(43384, 16),
59580 => conv_std_logic_vector(43616, 16),
59581 => conv_std_logic_vector(43848, 16),
59582 => conv_std_logic_vector(44080, 16),
59583 => conv_std_logic_vector(44312, 16),
59584 => conv_std_logic_vector(44544, 16),
59585 => conv_std_logic_vector(44776, 16),
59586 => conv_std_logic_vector(45008, 16),
59587 => conv_std_logic_vector(45240, 16),
59588 => conv_std_logic_vector(45472, 16),
59589 => conv_std_logic_vector(45704, 16),
59590 => conv_std_logic_vector(45936, 16),
59591 => conv_std_logic_vector(46168, 16),
59592 => conv_std_logic_vector(46400, 16),
59593 => conv_std_logic_vector(46632, 16),
59594 => conv_std_logic_vector(46864, 16),
59595 => conv_std_logic_vector(47096, 16),
59596 => conv_std_logic_vector(47328, 16),
59597 => conv_std_logic_vector(47560, 16),
59598 => conv_std_logic_vector(47792, 16),
59599 => conv_std_logic_vector(48024, 16),
59600 => conv_std_logic_vector(48256, 16),
59601 => conv_std_logic_vector(48488, 16),
59602 => conv_std_logic_vector(48720, 16),
59603 => conv_std_logic_vector(48952, 16),
59604 => conv_std_logic_vector(49184, 16),
59605 => conv_std_logic_vector(49416, 16),
59606 => conv_std_logic_vector(49648, 16),
59607 => conv_std_logic_vector(49880, 16),
59608 => conv_std_logic_vector(50112, 16),
59609 => conv_std_logic_vector(50344, 16),
59610 => conv_std_logic_vector(50576, 16),
59611 => conv_std_logic_vector(50808, 16),
59612 => conv_std_logic_vector(51040, 16),
59613 => conv_std_logic_vector(51272, 16),
59614 => conv_std_logic_vector(51504, 16),
59615 => conv_std_logic_vector(51736, 16),
59616 => conv_std_logic_vector(51968, 16),
59617 => conv_std_logic_vector(52200, 16),
59618 => conv_std_logic_vector(52432, 16),
59619 => conv_std_logic_vector(52664, 16),
59620 => conv_std_logic_vector(52896, 16),
59621 => conv_std_logic_vector(53128, 16),
59622 => conv_std_logic_vector(53360, 16),
59623 => conv_std_logic_vector(53592, 16),
59624 => conv_std_logic_vector(53824, 16),
59625 => conv_std_logic_vector(54056, 16),
59626 => conv_std_logic_vector(54288, 16),
59627 => conv_std_logic_vector(54520, 16),
59628 => conv_std_logic_vector(54752, 16),
59629 => conv_std_logic_vector(54984, 16),
59630 => conv_std_logic_vector(55216, 16),
59631 => conv_std_logic_vector(55448, 16),
59632 => conv_std_logic_vector(55680, 16),
59633 => conv_std_logic_vector(55912, 16),
59634 => conv_std_logic_vector(56144, 16),
59635 => conv_std_logic_vector(56376, 16),
59636 => conv_std_logic_vector(56608, 16),
59637 => conv_std_logic_vector(56840, 16),
59638 => conv_std_logic_vector(57072, 16),
59639 => conv_std_logic_vector(57304, 16),
59640 => conv_std_logic_vector(57536, 16),
59641 => conv_std_logic_vector(57768, 16),
59642 => conv_std_logic_vector(58000, 16),
59643 => conv_std_logic_vector(58232, 16),
59644 => conv_std_logic_vector(58464, 16),
59645 => conv_std_logic_vector(58696, 16),
59646 => conv_std_logic_vector(58928, 16),
59647 => conv_std_logic_vector(59160, 16),
59648 => conv_std_logic_vector(0, 16),
59649 => conv_std_logic_vector(233, 16),
59650 => conv_std_logic_vector(466, 16),
59651 => conv_std_logic_vector(699, 16),
59652 => conv_std_logic_vector(932, 16),
59653 => conv_std_logic_vector(1165, 16),
59654 => conv_std_logic_vector(1398, 16),
59655 => conv_std_logic_vector(1631, 16),
59656 => conv_std_logic_vector(1864, 16),
59657 => conv_std_logic_vector(2097, 16),
59658 => conv_std_logic_vector(2330, 16),
59659 => conv_std_logic_vector(2563, 16),
59660 => conv_std_logic_vector(2796, 16),
59661 => conv_std_logic_vector(3029, 16),
59662 => conv_std_logic_vector(3262, 16),
59663 => conv_std_logic_vector(3495, 16),
59664 => conv_std_logic_vector(3728, 16),
59665 => conv_std_logic_vector(3961, 16),
59666 => conv_std_logic_vector(4194, 16),
59667 => conv_std_logic_vector(4427, 16),
59668 => conv_std_logic_vector(4660, 16),
59669 => conv_std_logic_vector(4893, 16),
59670 => conv_std_logic_vector(5126, 16),
59671 => conv_std_logic_vector(5359, 16),
59672 => conv_std_logic_vector(5592, 16),
59673 => conv_std_logic_vector(5825, 16),
59674 => conv_std_logic_vector(6058, 16),
59675 => conv_std_logic_vector(6291, 16),
59676 => conv_std_logic_vector(6524, 16),
59677 => conv_std_logic_vector(6757, 16),
59678 => conv_std_logic_vector(6990, 16),
59679 => conv_std_logic_vector(7223, 16),
59680 => conv_std_logic_vector(7456, 16),
59681 => conv_std_logic_vector(7689, 16),
59682 => conv_std_logic_vector(7922, 16),
59683 => conv_std_logic_vector(8155, 16),
59684 => conv_std_logic_vector(8388, 16),
59685 => conv_std_logic_vector(8621, 16),
59686 => conv_std_logic_vector(8854, 16),
59687 => conv_std_logic_vector(9087, 16),
59688 => conv_std_logic_vector(9320, 16),
59689 => conv_std_logic_vector(9553, 16),
59690 => conv_std_logic_vector(9786, 16),
59691 => conv_std_logic_vector(10019, 16),
59692 => conv_std_logic_vector(10252, 16),
59693 => conv_std_logic_vector(10485, 16),
59694 => conv_std_logic_vector(10718, 16),
59695 => conv_std_logic_vector(10951, 16),
59696 => conv_std_logic_vector(11184, 16),
59697 => conv_std_logic_vector(11417, 16),
59698 => conv_std_logic_vector(11650, 16),
59699 => conv_std_logic_vector(11883, 16),
59700 => conv_std_logic_vector(12116, 16),
59701 => conv_std_logic_vector(12349, 16),
59702 => conv_std_logic_vector(12582, 16),
59703 => conv_std_logic_vector(12815, 16),
59704 => conv_std_logic_vector(13048, 16),
59705 => conv_std_logic_vector(13281, 16),
59706 => conv_std_logic_vector(13514, 16),
59707 => conv_std_logic_vector(13747, 16),
59708 => conv_std_logic_vector(13980, 16),
59709 => conv_std_logic_vector(14213, 16),
59710 => conv_std_logic_vector(14446, 16),
59711 => conv_std_logic_vector(14679, 16),
59712 => conv_std_logic_vector(14912, 16),
59713 => conv_std_logic_vector(15145, 16),
59714 => conv_std_logic_vector(15378, 16),
59715 => conv_std_logic_vector(15611, 16),
59716 => conv_std_logic_vector(15844, 16),
59717 => conv_std_logic_vector(16077, 16),
59718 => conv_std_logic_vector(16310, 16),
59719 => conv_std_logic_vector(16543, 16),
59720 => conv_std_logic_vector(16776, 16),
59721 => conv_std_logic_vector(17009, 16),
59722 => conv_std_logic_vector(17242, 16),
59723 => conv_std_logic_vector(17475, 16),
59724 => conv_std_logic_vector(17708, 16),
59725 => conv_std_logic_vector(17941, 16),
59726 => conv_std_logic_vector(18174, 16),
59727 => conv_std_logic_vector(18407, 16),
59728 => conv_std_logic_vector(18640, 16),
59729 => conv_std_logic_vector(18873, 16),
59730 => conv_std_logic_vector(19106, 16),
59731 => conv_std_logic_vector(19339, 16),
59732 => conv_std_logic_vector(19572, 16),
59733 => conv_std_logic_vector(19805, 16),
59734 => conv_std_logic_vector(20038, 16),
59735 => conv_std_logic_vector(20271, 16),
59736 => conv_std_logic_vector(20504, 16),
59737 => conv_std_logic_vector(20737, 16),
59738 => conv_std_logic_vector(20970, 16),
59739 => conv_std_logic_vector(21203, 16),
59740 => conv_std_logic_vector(21436, 16),
59741 => conv_std_logic_vector(21669, 16),
59742 => conv_std_logic_vector(21902, 16),
59743 => conv_std_logic_vector(22135, 16),
59744 => conv_std_logic_vector(22368, 16),
59745 => conv_std_logic_vector(22601, 16),
59746 => conv_std_logic_vector(22834, 16),
59747 => conv_std_logic_vector(23067, 16),
59748 => conv_std_logic_vector(23300, 16),
59749 => conv_std_logic_vector(23533, 16),
59750 => conv_std_logic_vector(23766, 16),
59751 => conv_std_logic_vector(23999, 16),
59752 => conv_std_logic_vector(24232, 16),
59753 => conv_std_logic_vector(24465, 16),
59754 => conv_std_logic_vector(24698, 16),
59755 => conv_std_logic_vector(24931, 16),
59756 => conv_std_logic_vector(25164, 16),
59757 => conv_std_logic_vector(25397, 16),
59758 => conv_std_logic_vector(25630, 16),
59759 => conv_std_logic_vector(25863, 16),
59760 => conv_std_logic_vector(26096, 16),
59761 => conv_std_logic_vector(26329, 16),
59762 => conv_std_logic_vector(26562, 16),
59763 => conv_std_logic_vector(26795, 16),
59764 => conv_std_logic_vector(27028, 16),
59765 => conv_std_logic_vector(27261, 16),
59766 => conv_std_logic_vector(27494, 16),
59767 => conv_std_logic_vector(27727, 16),
59768 => conv_std_logic_vector(27960, 16),
59769 => conv_std_logic_vector(28193, 16),
59770 => conv_std_logic_vector(28426, 16),
59771 => conv_std_logic_vector(28659, 16),
59772 => conv_std_logic_vector(28892, 16),
59773 => conv_std_logic_vector(29125, 16),
59774 => conv_std_logic_vector(29358, 16),
59775 => conv_std_logic_vector(29591, 16),
59776 => conv_std_logic_vector(29824, 16),
59777 => conv_std_logic_vector(30057, 16),
59778 => conv_std_logic_vector(30290, 16),
59779 => conv_std_logic_vector(30523, 16),
59780 => conv_std_logic_vector(30756, 16),
59781 => conv_std_logic_vector(30989, 16),
59782 => conv_std_logic_vector(31222, 16),
59783 => conv_std_logic_vector(31455, 16),
59784 => conv_std_logic_vector(31688, 16),
59785 => conv_std_logic_vector(31921, 16),
59786 => conv_std_logic_vector(32154, 16),
59787 => conv_std_logic_vector(32387, 16),
59788 => conv_std_logic_vector(32620, 16),
59789 => conv_std_logic_vector(32853, 16),
59790 => conv_std_logic_vector(33086, 16),
59791 => conv_std_logic_vector(33319, 16),
59792 => conv_std_logic_vector(33552, 16),
59793 => conv_std_logic_vector(33785, 16),
59794 => conv_std_logic_vector(34018, 16),
59795 => conv_std_logic_vector(34251, 16),
59796 => conv_std_logic_vector(34484, 16),
59797 => conv_std_logic_vector(34717, 16),
59798 => conv_std_logic_vector(34950, 16),
59799 => conv_std_logic_vector(35183, 16),
59800 => conv_std_logic_vector(35416, 16),
59801 => conv_std_logic_vector(35649, 16),
59802 => conv_std_logic_vector(35882, 16),
59803 => conv_std_logic_vector(36115, 16),
59804 => conv_std_logic_vector(36348, 16),
59805 => conv_std_logic_vector(36581, 16),
59806 => conv_std_logic_vector(36814, 16),
59807 => conv_std_logic_vector(37047, 16),
59808 => conv_std_logic_vector(37280, 16),
59809 => conv_std_logic_vector(37513, 16),
59810 => conv_std_logic_vector(37746, 16),
59811 => conv_std_logic_vector(37979, 16),
59812 => conv_std_logic_vector(38212, 16),
59813 => conv_std_logic_vector(38445, 16),
59814 => conv_std_logic_vector(38678, 16),
59815 => conv_std_logic_vector(38911, 16),
59816 => conv_std_logic_vector(39144, 16),
59817 => conv_std_logic_vector(39377, 16),
59818 => conv_std_logic_vector(39610, 16),
59819 => conv_std_logic_vector(39843, 16),
59820 => conv_std_logic_vector(40076, 16),
59821 => conv_std_logic_vector(40309, 16),
59822 => conv_std_logic_vector(40542, 16),
59823 => conv_std_logic_vector(40775, 16),
59824 => conv_std_logic_vector(41008, 16),
59825 => conv_std_logic_vector(41241, 16),
59826 => conv_std_logic_vector(41474, 16),
59827 => conv_std_logic_vector(41707, 16),
59828 => conv_std_logic_vector(41940, 16),
59829 => conv_std_logic_vector(42173, 16),
59830 => conv_std_logic_vector(42406, 16),
59831 => conv_std_logic_vector(42639, 16),
59832 => conv_std_logic_vector(42872, 16),
59833 => conv_std_logic_vector(43105, 16),
59834 => conv_std_logic_vector(43338, 16),
59835 => conv_std_logic_vector(43571, 16),
59836 => conv_std_logic_vector(43804, 16),
59837 => conv_std_logic_vector(44037, 16),
59838 => conv_std_logic_vector(44270, 16),
59839 => conv_std_logic_vector(44503, 16),
59840 => conv_std_logic_vector(44736, 16),
59841 => conv_std_logic_vector(44969, 16),
59842 => conv_std_logic_vector(45202, 16),
59843 => conv_std_logic_vector(45435, 16),
59844 => conv_std_logic_vector(45668, 16),
59845 => conv_std_logic_vector(45901, 16),
59846 => conv_std_logic_vector(46134, 16),
59847 => conv_std_logic_vector(46367, 16),
59848 => conv_std_logic_vector(46600, 16),
59849 => conv_std_logic_vector(46833, 16),
59850 => conv_std_logic_vector(47066, 16),
59851 => conv_std_logic_vector(47299, 16),
59852 => conv_std_logic_vector(47532, 16),
59853 => conv_std_logic_vector(47765, 16),
59854 => conv_std_logic_vector(47998, 16),
59855 => conv_std_logic_vector(48231, 16),
59856 => conv_std_logic_vector(48464, 16),
59857 => conv_std_logic_vector(48697, 16),
59858 => conv_std_logic_vector(48930, 16),
59859 => conv_std_logic_vector(49163, 16),
59860 => conv_std_logic_vector(49396, 16),
59861 => conv_std_logic_vector(49629, 16),
59862 => conv_std_logic_vector(49862, 16),
59863 => conv_std_logic_vector(50095, 16),
59864 => conv_std_logic_vector(50328, 16),
59865 => conv_std_logic_vector(50561, 16),
59866 => conv_std_logic_vector(50794, 16),
59867 => conv_std_logic_vector(51027, 16),
59868 => conv_std_logic_vector(51260, 16),
59869 => conv_std_logic_vector(51493, 16),
59870 => conv_std_logic_vector(51726, 16),
59871 => conv_std_logic_vector(51959, 16),
59872 => conv_std_logic_vector(52192, 16),
59873 => conv_std_logic_vector(52425, 16),
59874 => conv_std_logic_vector(52658, 16),
59875 => conv_std_logic_vector(52891, 16),
59876 => conv_std_logic_vector(53124, 16),
59877 => conv_std_logic_vector(53357, 16),
59878 => conv_std_logic_vector(53590, 16),
59879 => conv_std_logic_vector(53823, 16),
59880 => conv_std_logic_vector(54056, 16),
59881 => conv_std_logic_vector(54289, 16),
59882 => conv_std_logic_vector(54522, 16),
59883 => conv_std_logic_vector(54755, 16),
59884 => conv_std_logic_vector(54988, 16),
59885 => conv_std_logic_vector(55221, 16),
59886 => conv_std_logic_vector(55454, 16),
59887 => conv_std_logic_vector(55687, 16),
59888 => conv_std_logic_vector(55920, 16),
59889 => conv_std_logic_vector(56153, 16),
59890 => conv_std_logic_vector(56386, 16),
59891 => conv_std_logic_vector(56619, 16),
59892 => conv_std_logic_vector(56852, 16),
59893 => conv_std_logic_vector(57085, 16),
59894 => conv_std_logic_vector(57318, 16),
59895 => conv_std_logic_vector(57551, 16),
59896 => conv_std_logic_vector(57784, 16),
59897 => conv_std_logic_vector(58017, 16),
59898 => conv_std_logic_vector(58250, 16),
59899 => conv_std_logic_vector(58483, 16),
59900 => conv_std_logic_vector(58716, 16),
59901 => conv_std_logic_vector(58949, 16),
59902 => conv_std_logic_vector(59182, 16),
59903 => conv_std_logic_vector(59415, 16),
59904 => conv_std_logic_vector(0, 16),
59905 => conv_std_logic_vector(234, 16),
59906 => conv_std_logic_vector(468, 16),
59907 => conv_std_logic_vector(702, 16),
59908 => conv_std_logic_vector(936, 16),
59909 => conv_std_logic_vector(1170, 16),
59910 => conv_std_logic_vector(1404, 16),
59911 => conv_std_logic_vector(1638, 16),
59912 => conv_std_logic_vector(1872, 16),
59913 => conv_std_logic_vector(2106, 16),
59914 => conv_std_logic_vector(2340, 16),
59915 => conv_std_logic_vector(2574, 16),
59916 => conv_std_logic_vector(2808, 16),
59917 => conv_std_logic_vector(3042, 16),
59918 => conv_std_logic_vector(3276, 16),
59919 => conv_std_logic_vector(3510, 16),
59920 => conv_std_logic_vector(3744, 16),
59921 => conv_std_logic_vector(3978, 16),
59922 => conv_std_logic_vector(4212, 16),
59923 => conv_std_logic_vector(4446, 16),
59924 => conv_std_logic_vector(4680, 16),
59925 => conv_std_logic_vector(4914, 16),
59926 => conv_std_logic_vector(5148, 16),
59927 => conv_std_logic_vector(5382, 16),
59928 => conv_std_logic_vector(5616, 16),
59929 => conv_std_logic_vector(5850, 16),
59930 => conv_std_logic_vector(6084, 16),
59931 => conv_std_logic_vector(6318, 16),
59932 => conv_std_logic_vector(6552, 16),
59933 => conv_std_logic_vector(6786, 16),
59934 => conv_std_logic_vector(7020, 16),
59935 => conv_std_logic_vector(7254, 16),
59936 => conv_std_logic_vector(7488, 16),
59937 => conv_std_logic_vector(7722, 16),
59938 => conv_std_logic_vector(7956, 16),
59939 => conv_std_logic_vector(8190, 16),
59940 => conv_std_logic_vector(8424, 16),
59941 => conv_std_logic_vector(8658, 16),
59942 => conv_std_logic_vector(8892, 16),
59943 => conv_std_logic_vector(9126, 16),
59944 => conv_std_logic_vector(9360, 16),
59945 => conv_std_logic_vector(9594, 16),
59946 => conv_std_logic_vector(9828, 16),
59947 => conv_std_logic_vector(10062, 16),
59948 => conv_std_logic_vector(10296, 16),
59949 => conv_std_logic_vector(10530, 16),
59950 => conv_std_logic_vector(10764, 16),
59951 => conv_std_logic_vector(10998, 16),
59952 => conv_std_logic_vector(11232, 16),
59953 => conv_std_logic_vector(11466, 16),
59954 => conv_std_logic_vector(11700, 16),
59955 => conv_std_logic_vector(11934, 16),
59956 => conv_std_logic_vector(12168, 16),
59957 => conv_std_logic_vector(12402, 16),
59958 => conv_std_logic_vector(12636, 16),
59959 => conv_std_logic_vector(12870, 16),
59960 => conv_std_logic_vector(13104, 16),
59961 => conv_std_logic_vector(13338, 16),
59962 => conv_std_logic_vector(13572, 16),
59963 => conv_std_logic_vector(13806, 16),
59964 => conv_std_logic_vector(14040, 16),
59965 => conv_std_logic_vector(14274, 16),
59966 => conv_std_logic_vector(14508, 16),
59967 => conv_std_logic_vector(14742, 16),
59968 => conv_std_logic_vector(14976, 16),
59969 => conv_std_logic_vector(15210, 16),
59970 => conv_std_logic_vector(15444, 16),
59971 => conv_std_logic_vector(15678, 16),
59972 => conv_std_logic_vector(15912, 16),
59973 => conv_std_logic_vector(16146, 16),
59974 => conv_std_logic_vector(16380, 16),
59975 => conv_std_logic_vector(16614, 16),
59976 => conv_std_logic_vector(16848, 16),
59977 => conv_std_logic_vector(17082, 16),
59978 => conv_std_logic_vector(17316, 16),
59979 => conv_std_logic_vector(17550, 16),
59980 => conv_std_logic_vector(17784, 16),
59981 => conv_std_logic_vector(18018, 16),
59982 => conv_std_logic_vector(18252, 16),
59983 => conv_std_logic_vector(18486, 16),
59984 => conv_std_logic_vector(18720, 16),
59985 => conv_std_logic_vector(18954, 16),
59986 => conv_std_logic_vector(19188, 16),
59987 => conv_std_logic_vector(19422, 16),
59988 => conv_std_logic_vector(19656, 16),
59989 => conv_std_logic_vector(19890, 16),
59990 => conv_std_logic_vector(20124, 16),
59991 => conv_std_logic_vector(20358, 16),
59992 => conv_std_logic_vector(20592, 16),
59993 => conv_std_logic_vector(20826, 16),
59994 => conv_std_logic_vector(21060, 16),
59995 => conv_std_logic_vector(21294, 16),
59996 => conv_std_logic_vector(21528, 16),
59997 => conv_std_logic_vector(21762, 16),
59998 => conv_std_logic_vector(21996, 16),
59999 => conv_std_logic_vector(22230, 16),
60000 => conv_std_logic_vector(22464, 16),
60001 => conv_std_logic_vector(22698, 16),
60002 => conv_std_logic_vector(22932, 16),
60003 => conv_std_logic_vector(23166, 16),
60004 => conv_std_logic_vector(23400, 16),
60005 => conv_std_logic_vector(23634, 16),
60006 => conv_std_logic_vector(23868, 16),
60007 => conv_std_logic_vector(24102, 16),
60008 => conv_std_logic_vector(24336, 16),
60009 => conv_std_logic_vector(24570, 16),
60010 => conv_std_logic_vector(24804, 16),
60011 => conv_std_logic_vector(25038, 16),
60012 => conv_std_logic_vector(25272, 16),
60013 => conv_std_logic_vector(25506, 16),
60014 => conv_std_logic_vector(25740, 16),
60015 => conv_std_logic_vector(25974, 16),
60016 => conv_std_logic_vector(26208, 16),
60017 => conv_std_logic_vector(26442, 16),
60018 => conv_std_logic_vector(26676, 16),
60019 => conv_std_logic_vector(26910, 16),
60020 => conv_std_logic_vector(27144, 16),
60021 => conv_std_logic_vector(27378, 16),
60022 => conv_std_logic_vector(27612, 16),
60023 => conv_std_logic_vector(27846, 16),
60024 => conv_std_logic_vector(28080, 16),
60025 => conv_std_logic_vector(28314, 16),
60026 => conv_std_logic_vector(28548, 16),
60027 => conv_std_logic_vector(28782, 16),
60028 => conv_std_logic_vector(29016, 16),
60029 => conv_std_logic_vector(29250, 16),
60030 => conv_std_logic_vector(29484, 16),
60031 => conv_std_logic_vector(29718, 16),
60032 => conv_std_logic_vector(29952, 16),
60033 => conv_std_logic_vector(30186, 16),
60034 => conv_std_logic_vector(30420, 16),
60035 => conv_std_logic_vector(30654, 16),
60036 => conv_std_logic_vector(30888, 16),
60037 => conv_std_logic_vector(31122, 16),
60038 => conv_std_logic_vector(31356, 16),
60039 => conv_std_logic_vector(31590, 16),
60040 => conv_std_logic_vector(31824, 16),
60041 => conv_std_logic_vector(32058, 16),
60042 => conv_std_logic_vector(32292, 16),
60043 => conv_std_logic_vector(32526, 16),
60044 => conv_std_logic_vector(32760, 16),
60045 => conv_std_logic_vector(32994, 16),
60046 => conv_std_logic_vector(33228, 16),
60047 => conv_std_logic_vector(33462, 16),
60048 => conv_std_logic_vector(33696, 16),
60049 => conv_std_logic_vector(33930, 16),
60050 => conv_std_logic_vector(34164, 16),
60051 => conv_std_logic_vector(34398, 16),
60052 => conv_std_logic_vector(34632, 16),
60053 => conv_std_logic_vector(34866, 16),
60054 => conv_std_logic_vector(35100, 16),
60055 => conv_std_logic_vector(35334, 16),
60056 => conv_std_logic_vector(35568, 16),
60057 => conv_std_logic_vector(35802, 16),
60058 => conv_std_logic_vector(36036, 16),
60059 => conv_std_logic_vector(36270, 16),
60060 => conv_std_logic_vector(36504, 16),
60061 => conv_std_logic_vector(36738, 16),
60062 => conv_std_logic_vector(36972, 16),
60063 => conv_std_logic_vector(37206, 16),
60064 => conv_std_logic_vector(37440, 16),
60065 => conv_std_logic_vector(37674, 16),
60066 => conv_std_logic_vector(37908, 16),
60067 => conv_std_logic_vector(38142, 16),
60068 => conv_std_logic_vector(38376, 16),
60069 => conv_std_logic_vector(38610, 16),
60070 => conv_std_logic_vector(38844, 16),
60071 => conv_std_logic_vector(39078, 16),
60072 => conv_std_logic_vector(39312, 16),
60073 => conv_std_logic_vector(39546, 16),
60074 => conv_std_logic_vector(39780, 16),
60075 => conv_std_logic_vector(40014, 16),
60076 => conv_std_logic_vector(40248, 16),
60077 => conv_std_logic_vector(40482, 16),
60078 => conv_std_logic_vector(40716, 16),
60079 => conv_std_logic_vector(40950, 16),
60080 => conv_std_logic_vector(41184, 16),
60081 => conv_std_logic_vector(41418, 16),
60082 => conv_std_logic_vector(41652, 16),
60083 => conv_std_logic_vector(41886, 16),
60084 => conv_std_logic_vector(42120, 16),
60085 => conv_std_logic_vector(42354, 16),
60086 => conv_std_logic_vector(42588, 16),
60087 => conv_std_logic_vector(42822, 16),
60088 => conv_std_logic_vector(43056, 16),
60089 => conv_std_logic_vector(43290, 16),
60090 => conv_std_logic_vector(43524, 16),
60091 => conv_std_logic_vector(43758, 16),
60092 => conv_std_logic_vector(43992, 16),
60093 => conv_std_logic_vector(44226, 16),
60094 => conv_std_logic_vector(44460, 16),
60095 => conv_std_logic_vector(44694, 16),
60096 => conv_std_logic_vector(44928, 16),
60097 => conv_std_logic_vector(45162, 16),
60098 => conv_std_logic_vector(45396, 16),
60099 => conv_std_logic_vector(45630, 16),
60100 => conv_std_logic_vector(45864, 16),
60101 => conv_std_logic_vector(46098, 16),
60102 => conv_std_logic_vector(46332, 16),
60103 => conv_std_logic_vector(46566, 16),
60104 => conv_std_logic_vector(46800, 16),
60105 => conv_std_logic_vector(47034, 16),
60106 => conv_std_logic_vector(47268, 16),
60107 => conv_std_logic_vector(47502, 16),
60108 => conv_std_logic_vector(47736, 16),
60109 => conv_std_logic_vector(47970, 16),
60110 => conv_std_logic_vector(48204, 16),
60111 => conv_std_logic_vector(48438, 16),
60112 => conv_std_logic_vector(48672, 16),
60113 => conv_std_logic_vector(48906, 16),
60114 => conv_std_logic_vector(49140, 16),
60115 => conv_std_logic_vector(49374, 16),
60116 => conv_std_logic_vector(49608, 16),
60117 => conv_std_logic_vector(49842, 16),
60118 => conv_std_logic_vector(50076, 16),
60119 => conv_std_logic_vector(50310, 16),
60120 => conv_std_logic_vector(50544, 16),
60121 => conv_std_logic_vector(50778, 16),
60122 => conv_std_logic_vector(51012, 16),
60123 => conv_std_logic_vector(51246, 16),
60124 => conv_std_logic_vector(51480, 16),
60125 => conv_std_logic_vector(51714, 16),
60126 => conv_std_logic_vector(51948, 16),
60127 => conv_std_logic_vector(52182, 16),
60128 => conv_std_logic_vector(52416, 16),
60129 => conv_std_logic_vector(52650, 16),
60130 => conv_std_logic_vector(52884, 16),
60131 => conv_std_logic_vector(53118, 16),
60132 => conv_std_logic_vector(53352, 16),
60133 => conv_std_logic_vector(53586, 16),
60134 => conv_std_logic_vector(53820, 16),
60135 => conv_std_logic_vector(54054, 16),
60136 => conv_std_logic_vector(54288, 16),
60137 => conv_std_logic_vector(54522, 16),
60138 => conv_std_logic_vector(54756, 16),
60139 => conv_std_logic_vector(54990, 16),
60140 => conv_std_logic_vector(55224, 16),
60141 => conv_std_logic_vector(55458, 16),
60142 => conv_std_logic_vector(55692, 16),
60143 => conv_std_logic_vector(55926, 16),
60144 => conv_std_logic_vector(56160, 16),
60145 => conv_std_logic_vector(56394, 16),
60146 => conv_std_logic_vector(56628, 16),
60147 => conv_std_logic_vector(56862, 16),
60148 => conv_std_logic_vector(57096, 16),
60149 => conv_std_logic_vector(57330, 16),
60150 => conv_std_logic_vector(57564, 16),
60151 => conv_std_logic_vector(57798, 16),
60152 => conv_std_logic_vector(58032, 16),
60153 => conv_std_logic_vector(58266, 16),
60154 => conv_std_logic_vector(58500, 16),
60155 => conv_std_logic_vector(58734, 16),
60156 => conv_std_logic_vector(58968, 16),
60157 => conv_std_logic_vector(59202, 16),
60158 => conv_std_logic_vector(59436, 16),
60159 => conv_std_logic_vector(59670, 16),
60160 => conv_std_logic_vector(0, 16),
60161 => conv_std_logic_vector(235, 16),
60162 => conv_std_logic_vector(470, 16),
60163 => conv_std_logic_vector(705, 16),
60164 => conv_std_logic_vector(940, 16),
60165 => conv_std_logic_vector(1175, 16),
60166 => conv_std_logic_vector(1410, 16),
60167 => conv_std_logic_vector(1645, 16),
60168 => conv_std_logic_vector(1880, 16),
60169 => conv_std_logic_vector(2115, 16),
60170 => conv_std_logic_vector(2350, 16),
60171 => conv_std_logic_vector(2585, 16),
60172 => conv_std_logic_vector(2820, 16),
60173 => conv_std_logic_vector(3055, 16),
60174 => conv_std_logic_vector(3290, 16),
60175 => conv_std_logic_vector(3525, 16),
60176 => conv_std_logic_vector(3760, 16),
60177 => conv_std_logic_vector(3995, 16),
60178 => conv_std_logic_vector(4230, 16),
60179 => conv_std_logic_vector(4465, 16),
60180 => conv_std_logic_vector(4700, 16),
60181 => conv_std_logic_vector(4935, 16),
60182 => conv_std_logic_vector(5170, 16),
60183 => conv_std_logic_vector(5405, 16),
60184 => conv_std_logic_vector(5640, 16),
60185 => conv_std_logic_vector(5875, 16),
60186 => conv_std_logic_vector(6110, 16),
60187 => conv_std_logic_vector(6345, 16),
60188 => conv_std_logic_vector(6580, 16),
60189 => conv_std_logic_vector(6815, 16),
60190 => conv_std_logic_vector(7050, 16),
60191 => conv_std_logic_vector(7285, 16),
60192 => conv_std_logic_vector(7520, 16),
60193 => conv_std_logic_vector(7755, 16),
60194 => conv_std_logic_vector(7990, 16),
60195 => conv_std_logic_vector(8225, 16),
60196 => conv_std_logic_vector(8460, 16),
60197 => conv_std_logic_vector(8695, 16),
60198 => conv_std_logic_vector(8930, 16),
60199 => conv_std_logic_vector(9165, 16),
60200 => conv_std_logic_vector(9400, 16),
60201 => conv_std_logic_vector(9635, 16),
60202 => conv_std_logic_vector(9870, 16),
60203 => conv_std_logic_vector(10105, 16),
60204 => conv_std_logic_vector(10340, 16),
60205 => conv_std_logic_vector(10575, 16),
60206 => conv_std_logic_vector(10810, 16),
60207 => conv_std_logic_vector(11045, 16),
60208 => conv_std_logic_vector(11280, 16),
60209 => conv_std_logic_vector(11515, 16),
60210 => conv_std_logic_vector(11750, 16),
60211 => conv_std_logic_vector(11985, 16),
60212 => conv_std_logic_vector(12220, 16),
60213 => conv_std_logic_vector(12455, 16),
60214 => conv_std_logic_vector(12690, 16),
60215 => conv_std_logic_vector(12925, 16),
60216 => conv_std_logic_vector(13160, 16),
60217 => conv_std_logic_vector(13395, 16),
60218 => conv_std_logic_vector(13630, 16),
60219 => conv_std_logic_vector(13865, 16),
60220 => conv_std_logic_vector(14100, 16),
60221 => conv_std_logic_vector(14335, 16),
60222 => conv_std_logic_vector(14570, 16),
60223 => conv_std_logic_vector(14805, 16),
60224 => conv_std_logic_vector(15040, 16),
60225 => conv_std_logic_vector(15275, 16),
60226 => conv_std_logic_vector(15510, 16),
60227 => conv_std_logic_vector(15745, 16),
60228 => conv_std_logic_vector(15980, 16),
60229 => conv_std_logic_vector(16215, 16),
60230 => conv_std_logic_vector(16450, 16),
60231 => conv_std_logic_vector(16685, 16),
60232 => conv_std_logic_vector(16920, 16),
60233 => conv_std_logic_vector(17155, 16),
60234 => conv_std_logic_vector(17390, 16),
60235 => conv_std_logic_vector(17625, 16),
60236 => conv_std_logic_vector(17860, 16),
60237 => conv_std_logic_vector(18095, 16),
60238 => conv_std_logic_vector(18330, 16),
60239 => conv_std_logic_vector(18565, 16),
60240 => conv_std_logic_vector(18800, 16),
60241 => conv_std_logic_vector(19035, 16),
60242 => conv_std_logic_vector(19270, 16),
60243 => conv_std_logic_vector(19505, 16),
60244 => conv_std_logic_vector(19740, 16),
60245 => conv_std_logic_vector(19975, 16),
60246 => conv_std_logic_vector(20210, 16),
60247 => conv_std_logic_vector(20445, 16),
60248 => conv_std_logic_vector(20680, 16),
60249 => conv_std_logic_vector(20915, 16),
60250 => conv_std_logic_vector(21150, 16),
60251 => conv_std_logic_vector(21385, 16),
60252 => conv_std_logic_vector(21620, 16),
60253 => conv_std_logic_vector(21855, 16),
60254 => conv_std_logic_vector(22090, 16),
60255 => conv_std_logic_vector(22325, 16),
60256 => conv_std_logic_vector(22560, 16),
60257 => conv_std_logic_vector(22795, 16),
60258 => conv_std_logic_vector(23030, 16),
60259 => conv_std_logic_vector(23265, 16),
60260 => conv_std_logic_vector(23500, 16),
60261 => conv_std_logic_vector(23735, 16),
60262 => conv_std_logic_vector(23970, 16),
60263 => conv_std_logic_vector(24205, 16),
60264 => conv_std_logic_vector(24440, 16),
60265 => conv_std_logic_vector(24675, 16),
60266 => conv_std_logic_vector(24910, 16),
60267 => conv_std_logic_vector(25145, 16),
60268 => conv_std_logic_vector(25380, 16),
60269 => conv_std_logic_vector(25615, 16),
60270 => conv_std_logic_vector(25850, 16),
60271 => conv_std_logic_vector(26085, 16),
60272 => conv_std_logic_vector(26320, 16),
60273 => conv_std_logic_vector(26555, 16),
60274 => conv_std_logic_vector(26790, 16),
60275 => conv_std_logic_vector(27025, 16),
60276 => conv_std_logic_vector(27260, 16),
60277 => conv_std_logic_vector(27495, 16),
60278 => conv_std_logic_vector(27730, 16),
60279 => conv_std_logic_vector(27965, 16),
60280 => conv_std_logic_vector(28200, 16),
60281 => conv_std_logic_vector(28435, 16),
60282 => conv_std_logic_vector(28670, 16),
60283 => conv_std_logic_vector(28905, 16),
60284 => conv_std_logic_vector(29140, 16),
60285 => conv_std_logic_vector(29375, 16),
60286 => conv_std_logic_vector(29610, 16),
60287 => conv_std_logic_vector(29845, 16),
60288 => conv_std_logic_vector(30080, 16),
60289 => conv_std_logic_vector(30315, 16),
60290 => conv_std_logic_vector(30550, 16),
60291 => conv_std_logic_vector(30785, 16),
60292 => conv_std_logic_vector(31020, 16),
60293 => conv_std_logic_vector(31255, 16),
60294 => conv_std_logic_vector(31490, 16),
60295 => conv_std_logic_vector(31725, 16),
60296 => conv_std_logic_vector(31960, 16),
60297 => conv_std_logic_vector(32195, 16),
60298 => conv_std_logic_vector(32430, 16),
60299 => conv_std_logic_vector(32665, 16),
60300 => conv_std_logic_vector(32900, 16),
60301 => conv_std_logic_vector(33135, 16),
60302 => conv_std_logic_vector(33370, 16),
60303 => conv_std_logic_vector(33605, 16),
60304 => conv_std_logic_vector(33840, 16),
60305 => conv_std_logic_vector(34075, 16),
60306 => conv_std_logic_vector(34310, 16),
60307 => conv_std_logic_vector(34545, 16),
60308 => conv_std_logic_vector(34780, 16),
60309 => conv_std_logic_vector(35015, 16),
60310 => conv_std_logic_vector(35250, 16),
60311 => conv_std_logic_vector(35485, 16),
60312 => conv_std_logic_vector(35720, 16),
60313 => conv_std_logic_vector(35955, 16),
60314 => conv_std_logic_vector(36190, 16),
60315 => conv_std_logic_vector(36425, 16),
60316 => conv_std_logic_vector(36660, 16),
60317 => conv_std_logic_vector(36895, 16),
60318 => conv_std_logic_vector(37130, 16),
60319 => conv_std_logic_vector(37365, 16),
60320 => conv_std_logic_vector(37600, 16),
60321 => conv_std_logic_vector(37835, 16),
60322 => conv_std_logic_vector(38070, 16),
60323 => conv_std_logic_vector(38305, 16),
60324 => conv_std_logic_vector(38540, 16),
60325 => conv_std_logic_vector(38775, 16),
60326 => conv_std_logic_vector(39010, 16),
60327 => conv_std_logic_vector(39245, 16),
60328 => conv_std_logic_vector(39480, 16),
60329 => conv_std_logic_vector(39715, 16),
60330 => conv_std_logic_vector(39950, 16),
60331 => conv_std_logic_vector(40185, 16),
60332 => conv_std_logic_vector(40420, 16),
60333 => conv_std_logic_vector(40655, 16),
60334 => conv_std_logic_vector(40890, 16),
60335 => conv_std_logic_vector(41125, 16),
60336 => conv_std_logic_vector(41360, 16),
60337 => conv_std_logic_vector(41595, 16),
60338 => conv_std_logic_vector(41830, 16),
60339 => conv_std_logic_vector(42065, 16),
60340 => conv_std_logic_vector(42300, 16),
60341 => conv_std_logic_vector(42535, 16),
60342 => conv_std_logic_vector(42770, 16),
60343 => conv_std_logic_vector(43005, 16),
60344 => conv_std_logic_vector(43240, 16),
60345 => conv_std_logic_vector(43475, 16),
60346 => conv_std_logic_vector(43710, 16),
60347 => conv_std_logic_vector(43945, 16),
60348 => conv_std_logic_vector(44180, 16),
60349 => conv_std_logic_vector(44415, 16),
60350 => conv_std_logic_vector(44650, 16),
60351 => conv_std_logic_vector(44885, 16),
60352 => conv_std_logic_vector(45120, 16),
60353 => conv_std_logic_vector(45355, 16),
60354 => conv_std_logic_vector(45590, 16),
60355 => conv_std_logic_vector(45825, 16),
60356 => conv_std_logic_vector(46060, 16),
60357 => conv_std_logic_vector(46295, 16),
60358 => conv_std_logic_vector(46530, 16),
60359 => conv_std_logic_vector(46765, 16),
60360 => conv_std_logic_vector(47000, 16),
60361 => conv_std_logic_vector(47235, 16),
60362 => conv_std_logic_vector(47470, 16),
60363 => conv_std_logic_vector(47705, 16),
60364 => conv_std_logic_vector(47940, 16),
60365 => conv_std_logic_vector(48175, 16),
60366 => conv_std_logic_vector(48410, 16),
60367 => conv_std_logic_vector(48645, 16),
60368 => conv_std_logic_vector(48880, 16),
60369 => conv_std_logic_vector(49115, 16),
60370 => conv_std_logic_vector(49350, 16),
60371 => conv_std_logic_vector(49585, 16),
60372 => conv_std_logic_vector(49820, 16),
60373 => conv_std_logic_vector(50055, 16),
60374 => conv_std_logic_vector(50290, 16),
60375 => conv_std_logic_vector(50525, 16),
60376 => conv_std_logic_vector(50760, 16),
60377 => conv_std_logic_vector(50995, 16),
60378 => conv_std_logic_vector(51230, 16),
60379 => conv_std_logic_vector(51465, 16),
60380 => conv_std_logic_vector(51700, 16),
60381 => conv_std_logic_vector(51935, 16),
60382 => conv_std_logic_vector(52170, 16),
60383 => conv_std_logic_vector(52405, 16),
60384 => conv_std_logic_vector(52640, 16),
60385 => conv_std_logic_vector(52875, 16),
60386 => conv_std_logic_vector(53110, 16),
60387 => conv_std_logic_vector(53345, 16),
60388 => conv_std_logic_vector(53580, 16),
60389 => conv_std_logic_vector(53815, 16),
60390 => conv_std_logic_vector(54050, 16),
60391 => conv_std_logic_vector(54285, 16),
60392 => conv_std_logic_vector(54520, 16),
60393 => conv_std_logic_vector(54755, 16),
60394 => conv_std_logic_vector(54990, 16),
60395 => conv_std_logic_vector(55225, 16),
60396 => conv_std_logic_vector(55460, 16),
60397 => conv_std_logic_vector(55695, 16),
60398 => conv_std_logic_vector(55930, 16),
60399 => conv_std_logic_vector(56165, 16),
60400 => conv_std_logic_vector(56400, 16),
60401 => conv_std_logic_vector(56635, 16),
60402 => conv_std_logic_vector(56870, 16),
60403 => conv_std_logic_vector(57105, 16),
60404 => conv_std_logic_vector(57340, 16),
60405 => conv_std_logic_vector(57575, 16),
60406 => conv_std_logic_vector(57810, 16),
60407 => conv_std_logic_vector(58045, 16),
60408 => conv_std_logic_vector(58280, 16),
60409 => conv_std_logic_vector(58515, 16),
60410 => conv_std_logic_vector(58750, 16),
60411 => conv_std_logic_vector(58985, 16),
60412 => conv_std_logic_vector(59220, 16),
60413 => conv_std_logic_vector(59455, 16),
60414 => conv_std_logic_vector(59690, 16),
60415 => conv_std_logic_vector(59925, 16),
60416 => conv_std_logic_vector(0, 16),
60417 => conv_std_logic_vector(236, 16),
60418 => conv_std_logic_vector(472, 16),
60419 => conv_std_logic_vector(708, 16),
60420 => conv_std_logic_vector(944, 16),
60421 => conv_std_logic_vector(1180, 16),
60422 => conv_std_logic_vector(1416, 16),
60423 => conv_std_logic_vector(1652, 16),
60424 => conv_std_logic_vector(1888, 16),
60425 => conv_std_logic_vector(2124, 16),
60426 => conv_std_logic_vector(2360, 16),
60427 => conv_std_logic_vector(2596, 16),
60428 => conv_std_logic_vector(2832, 16),
60429 => conv_std_logic_vector(3068, 16),
60430 => conv_std_logic_vector(3304, 16),
60431 => conv_std_logic_vector(3540, 16),
60432 => conv_std_logic_vector(3776, 16),
60433 => conv_std_logic_vector(4012, 16),
60434 => conv_std_logic_vector(4248, 16),
60435 => conv_std_logic_vector(4484, 16),
60436 => conv_std_logic_vector(4720, 16),
60437 => conv_std_logic_vector(4956, 16),
60438 => conv_std_logic_vector(5192, 16),
60439 => conv_std_logic_vector(5428, 16),
60440 => conv_std_logic_vector(5664, 16),
60441 => conv_std_logic_vector(5900, 16),
60442 => conv_std_logic_vector(6136, 16),
60443 => conv_std_logic_vector(6372, 16),
60444 => conv_std_logic_vector(6608, 16),
60445 => conv_std_logic_vector(6844, 16),
60446 => conv_std_logic_vector(7080, 16),
60447 => conv_std_logic_vector(7316, 16),
60448 => conv_std_logic_vector(7552, 16),
60449 => conv_std_logic_vector(7788, 16),
60450 => conv_std_logic_vector(8024, 16),
60451 => conv_std_logic_vector(8260, 16),
60452 => conv_std_logic_vector(8496, 16),
60453 => conv_std_logic_vector(8732, 16),
60454 => conv_std_logic_vector(8968, 16),
60455 => conv_std_logic_vector(9204, 16),
60456 => conv_std_logic_vector(9440, 16),
60457 => conv_std_logic_vector(9676, 16),
60458 => conv_std_logic_vector(9912, 16),
60459 => conv_std_logic_vector(10148, 16),
60460 => conv_std_logic_vector(10384, 16),
60461 => conv_std_logic_vector(10620, 16),
60462 => conv_std_logic_vector(10856, 16),
60463 => conv_std_logic_vector(11092, 16),
60464 => conv_std_logic_vector(11328, 16),
60465 => conv_std_logic_vector(11564, 16),
60466 => conv_std_logic_vector(11800, 16),
60467 => conv_std_logic_vector(12036, 16),
60468 => conv_std_logic_vector(12272, 16),
60469 => conv_std_logic_vector(12508, 16),
60470 => conv_std_logic_vector(12744, 16),
60471 => conv_std_logic_vector(12980, 16),
60472 => conv_std_logic_vector(13216, 16),
60473 => conv_std_logic_vector(13452, 16),
60474 => conv_std_logic_vector(13688, 16),
60475 => conv_std_logic_vector(13924, 16),
60476 => conv_std_logic_vector(14160, 16),
60477 => conv_std_logic_vector(14396, 16),
60478 => conv_std_logic_vector(14632, 16),
60479 => conv_std_logic_vector(14868, 16),
60480 => conv_std_logic_vector(15104, 16),
60481 => conv_std_logic_vector(15340, 16),
60482 => conv_std_logic_vector(15576, 16),
60483 => conv_std_logic_vector(15812, 16),
60484 => conv_std_logic_vector(16048, 16),
60485 => conv_std_logic_vector(16284, 16),
60486 => conv_std_logic_vector(16520, 16),
60487 => conv_std_logic_vector(16756, 16),
60488 => conv_std_logic_vector(16992, 16),
60489 => conv_std_logic_vector(17228, 16),
60490 => conv_std_logic_vector(17464, 16),
60491 => conv_std_logic_vector(17700, 16),
60492 => conv_std_logic_vector(17936, 16),
60493 => conv_std_logic_vector(18172, 16),
60494 => conv_std_logic_vector(18408, 16),
60495 => conv_std_logic_vector(18644, 16),
60496 => conv_std_logic_vector(18880, 16),
60497 => conv_std_logic_vector(19116, 16),
60498 => conv_std_logic_vector(19352, 16),
60499 => conv_std_logic_vector(19588, 16),
60500 => conv_std_logic_vector(19824, 16),
60501 => conv_std_logic_vector(20060, 16),
60502 => conv_std_logic_vector(20296, 16),
60503 => conv_std_logic_vector(20532, 16),
60504 => conv_std_logic_vector(20768, 16),
60505 => conv_std_logic_vector(21004, 16),
60506 => conv_std_logic_vector(21240, 16),
60507 => conv_std_logic_vector(21476, 16),
60508 => conv_std_logic_vector(21712, 16),
60509 => conv_std_logic_vector(21948, 16),
60510 => conv_std_logic_vector(22184, 16),
60511 => conv_std_logic_vector(22420, 16),
60512 => conv_std_logic_vector(22656, 16),
60513 => conv_std_logic_vector(22892, 16),
60514 => conv_std_logic_vector(23128, 16),
60515 => conv_std_logic_vector(23364, 16),
60516 => conv_std_logic_vector(23600, 16),
60517 => conv_std_logic_vector(23836, 16),
60518 => conv_std_logic_vector(24072, 16),
60519 => conv_std_logic_vector(24308, 16),
60520 => conv_std_logic_vector(24544, 16),
60521 => conv_std_logic_vector(24780, 16),
60522 => conv_std_logic_vector(25016, 16),
60523 => conv_std_logic_vector(25252, 16),
60524 => conv_std_logic_vector(25488, 16),
60525 => conv_std_logic_vector(25724, 16),
60526 => conv_std_logic_vector(25960, 16),
60527 => conv_std_logic_vector(26196, 16),
60528 => conv_std_logic_vector(26432, 16),
60529 => conv_std_logic_vector(26668, 16),
60530 => conv_std_logic_vector(26904, 16),
60531 => conv_std_logic_vector(27140, 16),
60532 => conv_std_logic_vector(27376, 16),
60533 => conv_std_logic_vector(27612, 16),
60534 => conv_std_logic_vector(27848, 16),
60535 => conv_std_logic_vector(28084, 16),
60536 => conv_std_logic_vector(28320, 16),
60537 => conv_std_logic_vector(28556, 16),
60538 => conv_std_logic_vector(28792, 16),
60539 => conv_std_logic_vector(29028, 16),
60540 => conv_std_logic_vector(29264, 16),
60541 => conv_std_logic_vector(29500, 16),
60542 => conv_std_logic_vector(29736, 16),
60543 => conv_std_logic_vector(29972, 16),
60544 => conv_std_logic_vector(30208, 16),
60545 => conv_std_logic_vector(30444, 16),
60546 => conv_std_logic_vector(30680, 16),
60547 => conv_std_logic_vector(30916, 16),
60548 => conv_std_logic_vector(31152, 16),
60549 => conv_std_logic_vector(31388, 16),
60550 => conv_std_logic_vector(31624, 16),
60551 => conv_std_logic_vector(31860, 16),
60552 => conv_std_logic_vector(32096, 16),
60553 => conv_std_logic_vector(32332, 16),
60554 => conv_std_logic_vector(32568, 16),
60555 => conv_std_logic_vector(32804, 16),
60556 => conv_std_logic_vector(33040, 16),
60557 => conv_std_logic_vector(33276, 16),
60558 => conv_std_logic_vector(33512, 16),
60559 => conv_std_logic_vector(33748, 16),
60560 => conv_std_logic_vector(33984, 16),
60561 => conv_std_logic_vector(34220, 16),
60562 => conv_std_logic_vector(34456, 16),
60563 => conv_std_logic_vector(34692, 16),
60564 => conv_std_logic_vector(34928, 16),
60565 => conv_std_logic_vector(35164, 16),
60566 => conv_std_logic_vector(35400, 16),
60567 => conv_std_logic_vector(35636, 16),
60568 => conv_std_logic_vector(35872, 16),
60569 => conv_std_logic_vector(36108, 16),
60570 => conv_std_logic_vector(36344, 16),
60571 => conv_std_logic_vector(36580, 16),
60572 => conv_std_logic_vector(36816, 16),
60573 => conv_std_logic_vector(37052, 16),
60574 => conv_std_logic_vector(37288, 16),
60575 => conv_std_logic_vector(37524, 16),
60576 => conv_std_logic_vector(37760, 16),
60577 => conv_std_logic_vector(37996, 16),
60578 => conv_std_logic_vector(38232, 16),
60579 => conv_std_logic_vector(38468, 16),
60580 => conv_std_logic_vector(38704, 16),
60581 => conv_std_logic_vector(38940, 16),
60582 => conv_std_logic_vector(39176, 16),
60583 => conv_std_logic_vector(39412, 16),
60584 => conv_std_logic_vector(39648, 16),
60585 => conv_std_logic_vector(39884, 16),
60586 => conv_std_logic_vector(40120, 16),
60587 => conv_std_logic_vector(40356, 16),
60588 => conv_std_logic_vector(40592, 16),
60589 => conv_std_logic_vector(40828, 16),
60590 => conv_std_logic_vector(41064, 16),
60591 => conv_std_logic_vector(41300, 16),
60592 => conv_std_logic_vector(41536, 16),
60593 => conv_std_logic_vector(41772, 16),
60594 => conv_std_logic_vector(42008, 16),
60595 => conv_std_logic_vector(42244, 16),
60596 => conv_std_logic_vector(42480, 16),
60597 => conv_std_logic_vector(42716, 16),
60598 => conv_std_logic_vector(42952, 16),
60599 => conv_std_logic_vector(43188, 16),
60600 => conv_std_logic_vector(43424, 16),
60601 => conv_std_logic_vector(43660, 16),
60602 => conv_std_logic_vector(43896, 16),
60603 => conv_std_logic_vector(44132, 16),
60604 => conv_std_logic_vector(44368, 16),
60605 => conv_std_logic_vector(44604, 16),
60606 => conv_std_logic_vector(44840, 16),
60607 => conv_std_logic_vector(45076, 16),
60608 => conv_std_logic_vector(45312, 16),
60609 => conv_std_logic_vector(45548, 16),
60610 => conv_std_logic_vector(45784, 16),
60611 => conv_std_logic_vector(46020, 16),
60612 => conv_std_logic_vector(46256, 16),
60613 => conv_std_logic_vector(46492, 16),
60614 => conv_std_logic_vector(46728, 16),
60615 => conv_std_logic_vector(46964, 16),
60616 => conv_std_logic_vector(47200, 16),
60617 => conv_std_logic_vector(47436, 16),
60618 => conv_std_logic_vector(47672, 16),
60619 => conv_std_logic_vector(47908, 16),
60620 => conv_std_logic_vector(48144, 16),
60621 => conv_std_logic_vector(48380, 16),
60622 => conv_std_logic_vector(48616, 16),
60623 => conv_std_logic_vector(48852, 16),
60624 => conv_std_logic_vector(49088, 16),
60625 => conv_std_logic_vector(49324, 16),
60626 => conv_std_logic_vector(49560, 16),
60627 => conv_std_logic_vector(49796, 16),
60628 => conv_std_logic_vector(50032, 16),
60629 => conv_std_logic_vector(50268, 16),
60630 => conv_std_logic_vector(50504, 16),
60631 => conv_std_logic_vector(50740, 16),
60632 => conv_std_logic_vector(50976, 16),
60633 => conv_std_logic_vector(51212, 16),
60634 => conv_std_logic_vector(51448, 16),
60635 => conv_std_logic_vector(51684, 16),
60636 => conv_std_logic_vector(51920, 16),
60637 => conv_std_logic_vector(52156, 16),
60638 => conv_std_logic_vector(52392, 16),
60639 => conv_std_logic_vector(52628, 16),
60640 => conv_std_logic_vector(52864, 16),
60641 => conv_std_logic_vector(53100, 16),
60642 => conv_std_logic_vector(53336, 16),
60643 => conv_std_logic_vector(53572, 16),
60644 => conv_std_logic_vector(53808, 16),
60645 => conv_std_logic_vector(54044, 16),
60646 => conv_std_logic_vector(54280, 16),
60647 => conv_std_logic_vector(54516, 16),
60648 => conv_std_logic_vector(54752, 16),
60649 => conv_std_logic_vector(54988, 16),
60650 => conv_std_logic_vector(55224, 16),
60651 => conv_std_logic_vector(55460, 16),
60652 => conv_std_logic_vector(55696, 16),
60653 => conv_std_logic_vector(55932, 16),
60654 => conv_std_logic_vector(56168, 16),
60655 => conv_std_logic_vector(56404, 16),
60656 => conv_std_logic_vector(56640, 16),
60657 => conv_std_logic_vector(56876, 16),
60658 => conv_std_logic_vector(57112, 16),
60659 => conv_std_logic_vector(57348, 16),
60660 => conv_std_logic_vector(57584, 16),
60661 => conv_std_logic_vector(57820, 16),
60662 => conv_std_logic_vector(58056, 16),
60663 => conv_std_logic_vector(58292, 16),
60664 => conv_std_logic_vector(58528, 16),
60665 => conv_std_logic_vector(58764, 16),
60666 => conv_std_logic_vector(59000, 16),
60667 => conv_std_logic_vector(59236, 16),
60668 => conv_std_logic_vector(59472, 16),
60669 => conv_std_logic_vector(59708, 16),
60670 => conv_std_logic_vector(59944, 16),
60671 => conv_std_logic_vector(60180, 16),
60672 => conv_std_logic_vector(0, 16),
60673 => conv_std_logic_vector(237, 16),
60674 => conv_std_logic_vector(474, 16),
60675 => conv_std_logic_vector(711, 16),
60676 => conv_std_logic_vector(948, 16),
60677 => conv_std_logic_vector(1185, 16),
60678 => conv_std_logic_vector(1422, 16),
60679 => conv_std_logic_vector(1659, 16),
60680 => conv_std_logic_vector(1896, 16),
60681 => conv_std_logic_vector(2133, 16),
60682 => conv_std_logic_vector(2370, 16),
60683 => conv_std_logic_vector(2607, 16),
60684 => conv_std_logic_vector(2844, 16),
60685 => conv_std_logic_vector(3081, 16),
60686 => conv_std_logic_vector(3318, 16),
60687 => conv_std_logic_vector(3555, 16),
60688 => conv_std_logic_vector(3792, 16),
60689 => conv_std_logic_vector(4029, 16),
60690 => conv_std_logic_vector(4266, 16),
60691 => conv_std_logic_vector(4503, 16),
60692 => conv_std_logic_vector(4740, 16),
60693 => conv_std_logic_vector(4977, 16),
60694 => conv_std_logic_vector(5214, 16),
60695 => conv_std_logic_vector(5451, 16),
60696 => conv_std_logic_vector(5688, 16),
60697 => conv_std_logic_vector(5925, 16),
60698 => conv_std_logic_vector(6162, 16),
60699 => conv_std_logic_vector(6399, 16),
60700 => conv_std_logic_vector(6636, 16),
60701 => conv_std_logic_vector(6873, 16),
60702 => conv_std_logic_vector(7110, 16),
60703 => conv_std_logic_vector(7347, 16),
60704 => conv_std_logic_vector(7584, 16),
60705 => conv_std_logic_vector(7821, 16),
60706 => conv_std_logic_vector(8058, 16),
60707 => conv_std_logic_vector(8295, 16),
60708 => conv_std_logic_vector(8532, 16),
60709 => conv_std_logic_vector(8769, 16),
60710 => conv_std_logic_vector(9006, 16),
60711 => conv_std_logic_vector(9243, 16),
60712 => conv_std_logic_vector(9480, 16),
60713 => conv_std_logic_vector(9717, 16),
60714 => conv_std_logic_vector(9954, 16),
60715 => conv_std_logic_vector(10191, 16),
60716 => conv_std_logic_vector(10428, 16),
60717 => conv_std_logic_vector(10665, 16),
60718 => conv_std_logic_vector(10902, 16),
60719 => conv_std_logic_vector(11139, 16),
60720 => conv_std_logic_vector(11376, 16),
60721 => conv_std_logic_vector(11613, 16),
60722 => conv_std_logic_vector(11850, 16),
60723 => conv_std_logic_vector(12087, 16),
60724 => conv_std_logic_vector(12324, 16),
60725 => conv_std_logic_vector(12561, 16),
60726 => conv_std_logic_vector(12798, 16),
60727 => conv_std_logic_vector(13035, 16),
60728 => conv_std_logic_vector(13272, 16),
60729 => conv_std_logic_vector(13509, 16),
60730 => conv_std_logic_vector(13746, 16),
60731 => conv_std_logic_vector(13983, 16),
60732 => conv_std_logic_vector(14220, 16),
60733 => conv_std_logic_vector(14457, 16),
60734 => conv_std_logic_vector(14694, 16),
60735 => conv_std_logic_vector(14931, 16),
60736 => conv_std_logic_vector(15168, 16),
60737 => conv_std_logic_vector(15405, 16),
60738 => conv_std_logic_vector(15642, 16),
60739 => conv_std_logic_vector(15879, 16),
60740 => conv_std_logic_vector(16116, 16),
60741 => conv_std_logic_vector(16353, 16),
60742 => conv_std_logic_vector(16590, 16),
60743 => conv_std_logic_vector(16827, 16),
60744 => conv_std_logic_vector(17064, 16),
60745 => conv_std_logic_vector(17301, 16),
60746 => conv_std_logic_vector(17538, 16),
60747 => conv_std_logic_vector(17775, 16),
60748 => conv_std_logic_vector(18012, 16),
60749 => conv_std_logic_vector(18249, 16),
60750 => conv_std_logic_vector(18486, 16),
60751 => conv_std_logic_vector(18723, 16),
60752 => conv_std_logic_vector(18960, 16),
60753 => conv_std_logic_vector(19197, 16),
60754 => conv_std_logic_vector(19434, 16),
60755 => conv_std_logic_vector(19671, 16),
60756 => conv_std_logic_vector(19908, 16),
60757 => conv_std_logic_vector(20145, 16),
60758 => conv_std_logic_vector(20382, 16),
60759 => conv_std_logic_vector(20619, 16),
60760 => conv_std_logic_vector(20856, 16),
60761 => conv_std_logic_vector(21093, 16),
60762 => conv_std_logic_vector(21330, 16),
60763 => conv_std_logic_vector(21567, 16),
60764 => conv_std_logic_vector(21804, 16),
60765 => conv_std_logic_vector(22041, 16),
60766 => conv_std_logic_vector(22278, 16),
60767 => conv_std_logic_vector(22515, 16),
60768 => conv_std_logic_vector(22752, 16),
60769 => conv_std_logic_vector(22989, 16),
60770 => conv_std_logic_vector(23226, 16),
60771 => conv_std_logic_vector(23463, 16),
60772 => conv_std_logic_vector(23700, 16),
60773 => conv_std_logic_vector(23937, 16),
60774 => conv_std_logic_vector(24174, 16),
60775 => conv_std_logic_vector(24411, 16),
60776 => conv_std_logic_vector(24648, 16),
60777 => conv_std_logic_vector(24885, 16),
60778 => conv_std_logic_vector(25122, 16),
60779 => conv_std_logic_vector(25359, 16),
60780 => conv_std_logic_vector(25596, 16),
60781 => conv_std_logic_vector(25833, 16),
60782 => conv_std_logic_vector(26070, 16),
60783 => conv_std_logic_vector(26307, 16),
60784 => conv_std_logic_vector(26544, 16),
60785 => conv_std_logic_vector(26781, 16),
60786 => conv_std_logic_vector(27018, 16),
60787 => conv_std_logic_vector(27255, 16),
60788 => conv_std_logic_vector(27492, 16),
60789 => conv_std_logic_vector(27729, 16),
60790 => conv_std_logic_vector(27966, 16),
60791 => conv_std_logic_vector(28203, 16),
60792 => conv_std_logic_vector(28440, 16),
60793 => conv_std_logic_vector(28677, 16),
60794 => conv_std_logic_vector(28914, 16),
60795 => conv_std_logic_vector(29151, 16),
60796 => conv_std_logic_vector(29388, 16),
60797 => conv_std_logic_vector(29625, 16),
60798 => conv_std_logic_vector(29862, 16),
60799 => conv_std_logic_vector(30099, 16),
60800 => conv_std_logic_vector(30336, 16),
60801 => conv_std_logic_vector(30573, 16),
60802 => conv_std_logic_vector(30810, 16),
60803 => conv_std_logic_vector(31047, 16),
60804 => conv_std_logic_vector(31284, 16),
60805 => conv_std_logic_vector(31521, 16),
60806 => conv_std_logic_vector(31758, 16),
60807 => conv_std_logic_vector(31995, 16),
60808 => conv_std_logic_vector(32232, 16),
60809 => conv_std_logic_vector(32469, 16),
60810 => conv_std_logic_vector(32706, 16),
60811 => conv_std_logic_vector(32943, 16),
60812 => conv_std_logic_vector(33180, 16),
60813 => conv_std_logic_vector(33417, 16),
60814 => conv_std_logic_vector(33654, 16),
60815 => conv_std_logic_vector(33891, 16),
60816 => conv_std_logic_vector(34128, 16),
60817 => conv_std_logic_vector(34365, 16),
60818 => conv_std_logic_vector(34602, 16),
60819 => conv_std_logic_vector(34839, 16),
60820 => conv_std_logic_vector(35076, 16),
60821 => conv_std_logic_vector(35313, 16),
60822 => conv_std_logic_vector(35550, 16),
60823 => conv_std_logic_vector(35787, 16),
60824 => conv_std_logic_vector(36024, 16),
60825 => conv_std_logic_vector(36261, 16),
60826 => conv_std_logic_vector(36498, 16),
60827 => conv_std_logic_vector(36735, 16),
60828 => conv_std_logic_vector(36972, 16),
60829 => conv_std_logic_vector(37209, 16),
60830 => conv_std_logic_vector(37446, 16),
60831 => conv_std_logic_vector(37683, 16),
60832 => conv_std_logic_vector(37920, 16),
60833 => conv_std_logic_vector(38157, 16),
60834 => conv_std_logic_vector(38394, 16),
60835 => conv_std_logic_vector(38631, 16),
60836 => conv_std_logic_vector(38868, 16),
60837 => conv_std_logic_vector(39105, 16),
60838 => conv_std_logic_vector(39342, 16),
60839 => conv_std_logic_vector(39579, 16),
60840 => conv_std_logic_vector(39816, 16),
60841 => conv_std_logic_vector(40053, 16),
60842 => conv_std_logic_vector(40290, 16),
60843 => conv_std_logic_vector(40527, 16),
60844 => conv_std_logic_vector(40764, 16),
60845 => conv_std_logic_vector(41001, 16),
60846 => conv_std_logic_vector(41238, 16),
60847 => conv_std_logic_vector(41475, 16),
60848 => conv_std_logic_vector(41712, 16),
60849 => conv_std_logic_vector(41949, 16),
60850 => conv_std_logic_vector(42186, 16),
60851 => conv_std_logic_vector(42423, 16),
60852 => conv_std_logic_vector(42660, 16),
60853 => conv_std_logic_vector(42897, 16),
60854 => conv_std_logic_vector(43134, 16),
60855 => conv_std_logic_vector(43371, 16),
60856 => conv_std_logic_vector(43608, 16),
60857 => conv_std_logic_vector(43845, 16),
60858 => conv_std_logic_vector(44082, 16),
60859 => conv_std_logic_vector(44319, 16),
60860 => conv_std_logic_vector(44556, 16),
60861 => conv_std_logic_vector(44793, 16),
60862 => conv_std_logic_vector(45030, 16),
60863 => conv_std_logic_vector(45267, 16),
60864 => conv_std_logic_vector(45504, 16),
60865 => conv_std_logic_vector(45741, 16),
60866 => conv_std_logic_vector(45978, 16),
60867 => conv_std_logic_vector(46215, 16),
60868 => conv_std_logic_vector(46452, 16),
60869 => conv_std_logic_vector(46689, 16),
60870 => conv_std_logic_vector(46926, 16),
60871 => conv_std_logic_vector(47163, 16),
60872 => conv_std_logic_vector(47400, 16),
60873 => conv_std_logic_vector(47637, 16),
60874 => conv_std_logic_vector(47874, 16),
60875 => conv_std_logic_vector(48111, 16),
60876 => conv_std_logic_vector(48348, 16),
60877 => conv_std_logic_vector(48585, 16),
60878 => conv_std_logic_vector(48822, 16),
60879 => conv_std_logic_vector(49059, 16),
60880 => conv_std_logic_vector(49296, 16),
60881 => conv_std_logic_vector(49533, 16),
60882 => conv_std_logic_vector(49770, 16),
60883 => conv_std_logic_vector(50007, 16),
60884 => conv_std_logic_vector(50244, 16),
60885 => conv_std_logic_vector(50481, 16),
60886 => conv_std_logic_vector(50718, 16),
60887 => conv_std_logic_vector(50955, 16),
60888 => conv_std_logic_vector(51192, 16),
60889 => conv_std_logic_vector(51429, 16),
60890 => conv_std_logic_vector(51666, 16),
60891 => conv_std_logic_vector(51903, 16),
60892 => conv_std_logic_vector(52140, 16),
60893 => conv_std_logic_vector(52377, 16),
60894 => conv_std_logic_vector(52614, 16),
60895 => conv_std_logic_vector(52851, 16),
60896 => conv_std_logic_vector(53088, 16),
60897 => conv_std_logic_vector(53325, 16),
60898 => conv_std_logic_vector(53562, 16),
60899 => conv_std_logic_vector(53799, 16),
60900 => conv_std_logic_vector(54036, 16),
60901 => conv_std_logic_vector(54273, 16),
60902 => conv_std_logic_vector(54510, 16),
60903 => conv_std_logic_vector(54747, 16),
60904 => conv_std_logic_vector(54984, 16),
60905 => conv_std_logic_vector(55221, 16),
60906 => conv_std_logic_vector(55458, 16),
60907 => conv_std_logic_vector(55695, 16),
60908 => conv_std_logic_vector(55932, 16),
60909 => conv_std_logic_vector(56169, 16),
60910 => conv_std_logic_vector(56406, 16),
60911 => conv_std_logic_vector(56643, 16),
60912 => conv_std_logic_vector(56880, 16),
60913 => conv_std_logic_vector(57117, 16),
60914 => conv_std_logic_vector(57354, 16),
60915 => conv_std_logic_vector(57591, 16),
60916 => conv_std_logic_vector(57828, 16),
60917 => conv_std_logic_vector(58065, 16),
60918 => conv_std_logic_vector(58302, 16),
60919 => conv_std_logic_vector(58539, 16),
60920 => conv_std_logic_vector(58776, 16),
60921 => conv_std_logic_vector(59013, 16),
60922 => conv_std_logic_vector(59250, 16),
60923 => conv_std_logic_vector(59487, 16),
60924 => conv_std_logic_vector(59724, 16),
60925 => conv_std_logic_vector(59961, 16),
60926 => conv_std_logic_vector(60198, 16),
60927 => conv_std_logic_vector(60435, 16),
60928 => conv_std_logic_vector(0, 16),
60929 => conv_std_logic_vector(238, 16),
60930 => conv_std_logic_vector(476, 16),
60931 => conv_std_logic_vector(714, 16),
60932 => conv_std_logic_vector(952, 16),
60933 => conv_std_logic_vector(1190, 16),
60934 => conv_std_logic_vector(1428, 16),
60935 => conv_std_logic_vector(1666, 16),
60936 => conv_std_logic_vector(1904, 16),
60937 => conv_std_logic_vector(2142, 16),
60938 => conv_std_logic_vector(2380, 16),
60939 => conv_std_logic_vector(2618, 16),
60940 => conv_std_logic_vector(2856, 16),
60941 => conv_std_logic_vector(3094, 16),
60942 => conv_std_logic_vector(3332, 16),
60943 => conv_std_logic_vector(3570, 16),
60944 => conv_std_logic_vector(3808, 16),
60945 => conv_std_logic_vector(4046, 16),
60946 => conv_std_logic_vector(4284, 16),
60947 => conv_std_logic_vector(4522, 16),
60948 => conv_std_logic_vector(4760, 16),
60949 => conv_std_logic_vector(4998, 16),
60950 => conv_std_logic_vector(5236, 16),
60951 => conv_std_logic_vector(5474, 16),
60952 => conv_std_logic_vector(5712, 16),
60953 => conv_std_logic_vector(5950, 16),
60954 => conv_std_logic_vector(6188, 16),
60955 => conv_std_logic_vector(6426, 16),
60956 => conv_std_logic_vector(6664, 16),
60957 => conv_std_logic_vector(6902, 16),
60958 => conv_std_logic_vector(7140, 16),
60959 => conv_std_logic_vector(7378, 16),
60960 => conv_std_logic_vector(7616, 16),
60961 => conv_std_logic_vector(7854, 16),
60962 => conv_std_logic_vector(8092, 16),
60963 => conv_std_logic_vector(8330, 16),
60964 => conv_std_logic_vector(8568, 16),
60965 => conv_std_logic_vector(8806, 16),
60966 => conv_std_logic_vector(9044, 16),
60967 => conv_std_logic_vector(9282, 16),
60968 => conv_std_logic_vector(9520, 16),
60969 => conv_std_logic_vector(9758, 16),
60970 => conv_std_logic_vector(9996, 16),
60971 => conv_std_logic_vector(10234, 16),
60972 => conv_std_logic_vector(10472, 16),
60973 => conv_std_logic_vector(10710, 16),
60974 => conv_std_logic_vector(10948, 16),
60975 => conv_std_logic_vector(11186, 16),
60976 => conv_std_logic_vector(11424, 16),
60977 => conv_std_logic_vector(11662, 16),
60978 => conv_std_logic_vector(11900, 16),
60979 => conv_std_logic_vector(12138, 16),
60980 => conv_std_logic_vector(12376, 16),
60981 => conv_std_logic_vector(12614, 16),
60982 => conv_std_logic_vector(12852, 16),
60983 => conv_std_logic_vector(13090, 16),
60984 => conv_std_logic_vector(13328, 16),
60985 => conv_std_logic_vector(13566, 16),
60986 => conv_std_logic_vector(13804, 16),
60987 => conv_std_logic_vector(14042, 16),
60988 => conv_std_logic_vector(14280, 16),
60989 => conv_std_logic_vector(14518, 16),
60990 => conv_std_logic_vector(14756, 16),
60991 => conv_std_logic_vector(14994, 16),
60992 => conv_std_logic_vector(15232, 16),
60993 => conv_std_logic_vector(15470, 16),
60994 => conv_std_logic_vector(15708, 16),
60995 => conv_std_logic_vector(15946, 16),
60996 => conv_std_logic_vector(16184, 16),
60997 => conv_std_logic_vector(16422, 16),
60998 => conv_std_logic_vector(16660, 16),
60999 => conv_std_logic_vector(16898, 16),
61000 => conv_std_logic_vector(17136, 16),
61001 => conv_std_logic_vector(17374, 16),
61002 => conv_std_logic_vector(17612, 16),
61003 => conv_std_logic_vector(17850, 16),
61004 => conv_std_logic_vector(18088, 16),
61005 => conv_std_logic_vector(18326, 16),
61006 => conv_std_logic_vector(18564, 16),
61007 => conv_std_logic_vector(18802, 16),
61008 => conv_std_logic_vector(19040, 16),
61009 => conv_std_logic_vector(19278, 16),
61010 => conv_std_logic_vector(19516, 16),
61011 => conv_std_logic_vector(19754, 16),
61012 => conv_std_logic_vector(19992, 16),
61013 => conv_std_logic_vector(20230, 16),
61014 => conv_std_logic_vector(20468, 16),
61015 => conv_std_logic_vector(20706, 16),
61016 => conv_std_logic_vector(20944, 16),
61017 => conv_std_logic_vector(21182, 16),
61018 => conv_std_logic_vector(21420, 16),
61019 => conv_std_logic_vector(21658, 16),
61020 => conv_std_logic_vector(21896, 16),
61021 => conv_std_logic_vector(22134, 16),
61022 => conv_std_logic_vector(22372, 16),
61023 => conv_std_logic_vector(22610, 16),
61024 => conv_std_logic_vector(22848, 16),
61025 => conv_std_logic_vector(23086, 16),
61026 => conv_std_logic_vector(23324, 16),
61027 => conv_std_logic_vector(23562, 16),
61028 => conv_std_logic_vector(23800, 16),
61029 => conv_std_logic_vector(24038, 16),
61030 => conv_std_logic_vector(24276, 16),
61031 => conv_std_logic_vector(24514, 16),
61032 => conv_std_logic_vector(24752, 16),
61033 => conv_std_logic_vector(24990, 16),
61034 => conv_std_logic_vector(25228, 16),
61035 => conv_std_logic_vector(25466, 16),
61036 => conv_std_logic_vector(25704, 16),
61037 => conv_std_logic_vector(25942, 16),
61038 => conv_std_logic_vector(26180, 16),
61039 => conv_std_logic_vector(26418, 16),
61040 => conv_std_logic_vector(26656, 16),
61041 => conv_std_logic_vector(26894, 16),
61042 => conv_std_logic_vector(27132, 16),
61043 => conv_std_logic_vector(27370, 16),
61044 => conv_std_logic_vector(27608, 16),
61045 => conv_std_logic_vector(27846, 16),
61046 => conv_std_logic_vector(28084, 16),
61047 => conv_std_logic_vector(28322, 16),
61048 => conv_std_logic_vector(28560, 16),
61049 => conv_std_logic_vector(28798, 16),
61050 => conv_std_logic_vector(29036, 16),
61051 => conv_std_logic_vector(29274, 16),
61052 => conv_std_logic_vector(29512, 16),
61053 => conv_std_logic_vector(29750, 16),
61054 => conv_std_logic_vector(29988, 16),
61055 => conv_std_logic_vector(30226, 16),
61056 => conv_std_logic_vector(30464, 16),
61057 => conv_std_logic_vector(30702, 16),
61058 => conv_std_logic_vector(30940, 16),
61059 => conv_std_logic_vector(31178, 16),
61060 => conv_std_logic_vector(31416, 16),
61061 => conv_std_logic_vector(31654, 16),
61062 => conv_std_logic_vector(31892, 16),
61063 => conv_std_logic_vector(32130, 16),
61064 => conv_std_logic_vector(32368, 16),
61065 => conv_std_logic_vector(32606, 16),
61066 => conv_std_logic_vector(32844, 16),
61067 => conv_std_logic_vector(33082, 16),
61068 => conv_std_logic_vector(33320, 16),
61069 => conv_std_logic_vector(33558, 16),
61070 => conv_std_logic_vector(33796, 16),
61071 => conv_std_logic_vector(34034, 16),
61072 => conv_std_logic_vector(34272, 16),
61073 => conv_std_logic_vector(34510, 16),
61074 => conv_std_logic_vector(34748, 16),
61075 => conv_std_logic_vector(34986, 16),
61076 => conv_std_logic_vector(35224, 16),
61077 => conv_std_logic_vector(35462, 16),
61078 => conv_std_logic_vector(35700, 16),
61079 => conv_std_logic_vector(35938, 16),
61080 => conv_std_logic_vector(36176, 16),
61081 => conv_std_logic_vector(36414, 16),
61082 => conv_std_logic_vector(36652, 16),
61083 => conv_std_logic_vector(36890, 16),
61084 => conv_std_logic_vector(37128, 16),
61085 => conv_std_logic_vector(37366, 16),
61086 => conv_std_logic_vector(37604, 16),
61087 => conv_std_logic_vector(37842, 16),
61088 => conv_std_logic_vector(38080, 16),
61089 => conv_std_logic_vector(38318, 16),
61090 => conv_std_logic_vector(38556, 16),
61091 => conv_std_logic_vector(38794, 16),
61092 => conv_std_logic_vector(39032, 16),
61093 => conv_std_logic_vector(39270, 16),
61094 => conv_std_logic_vector(39508, 16),
61095 => conv_std_logic_vector(39746, 16),
61096 => conv_std_logic_vector(39984, 16),
61097 => conv_std_logic_vector(40222, 16),
61098 => conv_std_logic_vector(40460, 16),
61099 => conv_std_logic_vector(40698, 16),
61100 => conv_std_logic_vector(40936, 16),
61101 => conv_std_logic_vector(41174, 16),
61102 => conv_std_logic_vector(41412, 16),
61103 => conv_std_logic_vector(41650, 16),
61104 => conv_std_logic_vector(41888, 16),
61105 => conv_std_logic_vector(42126, 16),
61106 => conv_std_logic_vector(42364, 16),
61107 => conv_std_logic_vector(42602, 16),
61108 => conv_std_logic_vector(42840, 16),
61109 => conv_std_logic_vector(43078, 16),
61110 => conv_std_logic_vector(43316, 16),
61111 => conv_std_logic_vector(43554, 16),
61112 => conv_std_logic_vector(43792, 16),
61113 => conv_std_logic_vector(44030, 16),
61114 => conv_std_logic_vector(44268, 16),
61115 => conv_std_logic_vector(44506, 16),
61116 => conv_std_logic_vector(44744, 16),
61117 => conv_std_logic_vector(44982, 16),
61118 => conv_std_logic_vector(45220, 16),
61119 => conv_std_logic_vector(45458, 16),
61120 => conv_std_logic_vector(45696, 16),
61121 => conv_std_logic_vector(45934, 16),
61122 => conv_std_logic_vector(46172, 16),
61123 => conv_std_logic_vector(46410, 16),
61124 => conv_std_logic_vector(46648, 16),
61125 => conv_std_logic_vector(46886, 16),
61126 => conv_std_logic_vector(47124, 16),
61127 => conv_std_logic_vector(47362, 16),
61128 => conv_std_logic_vector(47600, 16),
61129 => conv_std_logic_vector(47838, 16),
61130 => conv_std_logic_vector(48076, 16),
61131 => conv_std_logic_vector(48314, 16),
61132 => conv_std_logic_vector(48552, 16),
61133 => conv_std_logic_vector(48790, 16),
61134 => conv_std_logic_vector(49028, 16),
61135 => conv_std_logic_vector(49266, 16),
61136 => conv_std_logic_vector(49504, 16),
61137 => conv_std_logic_vector(49742, 16),
61138 => conv_std_logic_vector(49980, 16),
61139 => conv_std_logic_vector(50218, 16),
61140 => conv_std_logic_vector(50456, 16),
61141 => conv_std_logic_vector(50694, 16),
61142 => conv_std_logic_vector(50932, 16),
61143 => conv_std_logic_vector(51170, 16),
61144 => conv_std_logic_vector(51408, 16),
61145 => conv_std_logic_vector(51646, 16),
61146 => conv_std_logic_vector(51884, 16),
61147 => conv_std_logic_vector(52122, 16),
61148 => conv_std_logic_vector(52360, 16),
61149 => conv_std_logic_vector(52598, 16),
61150 => conv_std_logic_vector(52836, 16),
61151 => conv_std_logic_vector(53074, 16),
61152 => conv_std_logic_vector(53312, 16),
61153 => conv_std_logic_vector(53550, 16),
61154 => conv_std_logic_vector(53788, 16),
61155 => conv_std_logic_vector(54026, 16),
61156 => conv_std_logic_vector(54264, 16),
61157 => conv_std_logic_vector(54502, 16),
61158 => conv_std_logic_vector(54740, 16),
61159 => conv_std_logic_vector(54978, 16),
61160 => conv_std_logic_vector(55216, 16),
61161 => conv_std_logic_vector(55454, 16),
61162 => conv_std_logic_vector(55692, 16),
61163 => conv_std_logic_vector(55930, 16),
61164 => conv_std_logic_vector(56168, 16),
61165 => conv_std_logic_vector(56406, 16),
61166 => conv_std_logic_vector(56644, 16),
61167 => conv_std_logic_vector(56882, 16),
61168 => conv_std_logic_vector(57120, 16),
61169 => conv_std_logic_vector(57358, 16),
61170 => conv_std_logic_vector(57596, 16),
61171 => conv_std_logic_vector(57834, 16),
61172 => conv_std_logic_vector(58072, 16),
61173 => conv_std_logic_vector(58310, 16),
61174 => conv_std_logic_vector(58548, 16),
61175 => conv_std_logic_vector(58786, 16),
61176 => conv_std_logic_vector(59024, 16),
61177 => conv_std_logic_vector(59262, 16),
61178 => conv_std_logic_vector(59500, 16),
61179 => conv_std_logic_vector(59738, 16),
61180 => conv_std_logic_vector(59976, 16),
61181 => conv_std_logic_vector(60214, 16),
61182 => conv_std_logic_vector(60452, 16),
61183 => conv_std_logic_vector(60690, 16),
61184 => conv_std_logic_vector(0, 16),
61185 => conv_std_logic_vector(239, 16),
61186 => conv_std_logic_vector(478, 16),
61187 => conv_std_logic_vector(717, 16),
61188 => conv_std_logic_vector(956, 16),
61189 => conv_std_logic_vector(1195, 16),
61190 => conv_std_logic_vector(1434, 16),
61191 => conv_std_logic_vector(1673, 16),
61192 => conv_std_logic_vector(1912, 16),
61193 => conv_std_logic_vector(2151, 16),
61194 => conv_std_logic_vector(2390, 16),
61195 => conv_std_logic_vector(2629, 16),
61196 => conv_std_logic_vector(2868, 16),
61197 => conv_std_logic_vector(3107, 16),
61198 => conv_std_logic_vector(3346, 16),
61199 => conv_std_logic_vector(3585, 16),
61200 => conv_std_logic_vector(3824, 16),
61201 => conv_std_logic_vector(4063, 16),
61202 => conv_std_logic_vector(4302, 16),
61203 => conv_std_logic_vector(4541, 16),
61204 => conv_std_logic_vector(4780, 16),
61205 => conv_std_logic_vector(5019, 16),
61206 => conv_std_logic_vector(5258, 16),
61207 => conv_std_logic_vector(5497, 16),
61208 => conv_std_logic_vector(5736, 16),
61209 => conv_std_logic_vector(5975, 16),
61210 => conv_std_logic_vector(6214, 16),
61211 => conv_std_logic_vector(6453, 16),
61212 => conv_std_logic_vector(6692, 16),
61213 => conv_std_logic_vector(6931, 16),
61214 => conv_std_logic_vector(7170, 16),
61215 => conv_std_logic_vector(7409, 16),
61216 => conv_std_logic_vector(7648, 16),
61217 => conv_std_logic_vector(7887, 16),
61218 => conv_std_logic_vector(8126, 16),
61219 => conv_std_logic_vector(8365, 16),
61220 => conv_std_logic_vector(8604, 16),
61221 => conv_std_logic_vector(8843, 16),
61222 => conv_std_logic_vector(9082, 16),
61223 => conv_std_logic_vector(9321, 16),
61224 => conv_std_logic_vector(9560, 16),
61225 => conv_std_logic_vector(9799, 16),
61226 => conv_std_logic_vector(10038, 16),
61227 => conv_std_logic_vector(10277, 16),
61228 => conv_std_logic_vector(10516, 16),
61229 => conv_std_logic_vector(10755, 16),
61230 => conv_std_logic_vector(10994, 16),
61231 => conv_std_logic_vector(11233, 16),
61232 => conv_std_logic_vector(11472, 16),
61233 => conv_std_logic_vector(11711, 16),
61234 => conv_std_logic_vector(11950, 16),
61235 => conv_std_logic_vector(12189, 16),
61236 => conv_std_logic_vector(12428, 16),
61237 => conv_std_logic_vector(12667, 16),
61238 => conv_std_logic_vector(12906, 16),
61239 => conv_std_logic_vector(13145, 16),
61240 => conv_std_logic_vector(13384, 16),
61241 => conv_std_logic_vector(13623, 16),
61242 => conv_std_logic_vector(13862, 16),
61243 => conv_std_logic_vector(14101, 16),
61244 => conv_std_logic_vector(14340, 16),
61245 => conv_std_logic_vector(14579, 16),
61246 => conv_std_logic_vector(14818, 16),
61247 => conv_std_logic_vector(15057, 16),
61248 => conv_std_logic_vector(15296, 16),
61249 => conv_std_logic_vector(15535, 16),
61250 => conv_std_logic_vector(15774, 16),
61251 => conv_std_logic_vector(16013, 16),
61252 => conv_std_logic_vector(16252, 16),
61253 => conv_std_logic_vector(16491, 16),
61254 => conv_std_logic_vector(16730, 16),
61255 => conv_std_logic_vector(16969, 16),
61256 => conv_std_logic_vector(17208, 16),
61257 => conv_std_logic_vector(17447, 16),
61258 => conv_std_logic_vector(17686, 16),
61259 => conv_std_logic_vector(17925, 16),
61260 => conv_std_logic_vector(18164, 16),
61261 => conv_std_logic_vector(18403, 16),
61262 => conv_std_logic_vector(18642, 16),
61263 => conv_std_logic_vector(18881, 16),
61264 => conv_std_logic_vector(19120, 16),
61265 => conv_std_logic_vector(19359, 16),
61266 => conv_std_logic_vector(19598, 16),
61267 => conv_std_logic_vector(19837, 16),
61268 => conv_std_logic_vector(20076, 16),
61269 => conv_std_logic_vector(20315, 16),
61270 => conv_std_logic_vector(20554, 16),
61271 => conv_std_logic_vector(20793, 16),
61272 => conv_std_logic_vector(21032, 16),
61273 => conv_std_logic_vector(21271, 16),
61274 => conv_std_logic_vector(21510, 16),
61275 => conv_std_logic_vector(21749, 16),
61276 => conv_std_logic_vector(21988, 16),
61277 => conv_std_logic_vector(22227, 16),
61278 => conv_std_logic_vector(22466, 16),
61279 => conv_std_logic_vector(22705, 16),
61280 => conv_std_logic_vector(22944, 16),
61281 => conv_std_logic_vector(23183, 16),
61282 => conv_std_logic_vector(23422, 16),
61283 => conv_std_logic_vector(23661, 16),
61284 => conv_std_logic_vector(23900, 16),
61285 => conv_std_logic_vector(24139, 16),
61286 => conv_std_logic_vector(24378, 16),
61287 => conv_std_logic_vector(24617, 16),
61288 => conv_std_logic_vector(24856, 16),
61289 => conv_std_logic_vector(25095, 16),
61290 => conv_std_logic_vector(25334, 16),
61291 => conv_std_logic_vector(25573, 16),
61292 => conv_std_logic_vector(25812, 16),
61293 => conv_std_logic_vector(26051, 16),
61294 => conv_std_logic_vector(26290, 16),
61295 => conv_std_logic_vector(26529, 16),
61296 => conv_std_logic_vector(26768, 16),
61297 => conv_std_logic_vector(27007, 16),
61298 => conv_std_logic_vector(27246, 16),
61299 => conv_std_logic_vector(27485, 16),
61300 => conv_std_logic_vector(27724, 16),
61301 => conv_std_logic_vector(27963, 16),
61302 => conv_std_logic_vector(28202, 16),
61303 => conv_std_logic_vector(28441, 16),
61304 => conv_std_logic_vector(28680, 16),
61305 => conv_std_logic_vector(28919, 16),
61306 => conv_std_logic_vector(29158, 16),
61307 => conv_std_logic_vector(29397, 16),
61308 => conv_std_logic_vector(29636, 16),
61309 => conv_std_logic_vector(29875, 16),
61310 => conv_std_logic_vector(30114, 16),
61311 => conv_std_logic_vector(30353, 16),
61312 => conv_std_logic_vector(30592, 16),
61313 => conv_std_logic_vector(30831, 16),
61314 => conv_std_logic_vector(31070, 16),
61315 => conv_std_logic_vector(31309, 16),
61316 => conv_std_logic_vector(31548, 16),
61317 => conv_std_logic_vector(31787, 16),
61318 => conv_std_logic_vector(32026, 16),
61319 => conv_std_logic_vector(32265, 16),
61320 => conv_std_logic_vector(32504, 16),
61321 => conv_std_logic_vector(32743, 16),
61322 => conv_std_logic_vector(32982, 16),
61323 => conv_std_logic_vector(33221, 16),
61324 => conv_std_logic_vector(33460, 16),
61325 => conv_std_logic_vector(33699, 16),
61326 => conv_std_logic_vector(33938, 16),
61327 => conv_std_logic_vector(34177, 16),
61328 => conv_std_logic_vector(34416, 16),
61329 => conv_std_logic_vector(34655, 16),
61330 => conv_std_logic_vector(34894, 16),
61331 => conv_std_logic_vector(35133, 16),
61332 => conv_std_logic_vector(35372, 16),
61333 => conv_std_logic_vector(35611, 16),
61334 => conv_std_logic_vector(35850, 16),
61335 => conv_std_logic_vector(36089, 16),
61336 => conv_std_logic_vector(36328, 16),
61337 => conv_std_logic_vector(36567, 16),
61338 => conv_std_logic_vector(36806, 16),
61339 => conv_std_logic_vector(37045, 16),
61340 => conv_std_logic_vector(37284, 16),
61341 => conv_std_logic_vector(37523, 16),
61342 => conv_std_logic_vector(37762, 16),
61343 => conv_std_logic_vector(38001, 16),
61344 => conv_std_logic_vector(38240, 16),
61345 => conv_std_logic_vector(38479, 16),
61346 => conv_std_logic_vector(38718, 16),
61347 => conv_std_logic_vector(38957, 16),
61348 => conv_std_logic_vector(39196, 16),
61349 => conv_std_logic_vector(39435, 16),
61350 => conv_std_logic_vector(39674, 16),
61351 => conv_std_logic_vector(39913, 16),
61352 => conv_std_logic_vector(40152, 16),
61353 => conv_std_logic_vector(40391, 16),
61354 => conv_std_logic_vector(40630, 16),
61355 => conv_std_logic_vector(40869, 16),
61356 => conv_std_logic_vector(41108, 16),
61357 => conv_std_logic_vector(41347, 16),
61358 => conv_std_logic_vector(41586, 16),
61359 => conv_std_logic_vector(41825, 16),
61360 => conv_std_logic_vector(42064, 16),
61361 => conv_std_logic_vector(42303, 16),
61362 => conv_std_logic_vector(42542, 16),
61363 => conv_std_logic_vector(42781, 16),
61364 => conv_std_logic_vector(43020, 16),
61365 => conv_std_logic_vector(43259, 16),
61366 => conv_std_logic_vector(43498, 16),
61367 => conv_std_logic_vector(43737, 16),
61368 => conv_std_logic_vector(43976, 16),
61369 => conv_std_logic_vector(44215, 16),
61370 => conv_std_logic_vector(44454, 16),
61371 => conv_std_logic_vector(44693, 16),
61372 => conv_std_logic_vector(44932, 16),
61373 => conv_std_logic_vector(45171, 16),
61374 => conv_std_logic_vector(45410, 16),
61375 => conv_std_logic_vector(45649, 16),
61376 => conv_std_logic_vector(45888, 16),
61377 => conv_std_logic_vector(46127, 16),
61378 => conv_std_logic_vector(46366, 16),
61379 => conv_std_logic_vector(46605, 16),
61380 => conv_std_logic_vector(46844, 16),
61381 => conv_std_logic_vector(47083, 16),
61382 => conv_std_logic_vector(47322, 16),
61383 => conv_std_logic_vector(47561, 16),
61384 => conv_std_logic_vector(47800, 16),
61385 => conv_std_logic_vector(48039, 16),
61386 => conv_std_logic_vector(48278, 16),
61387 => conv_std_logic_vector(48517, 16),
61388 => conv_std_logic_vector(48756, 16),
61389 => conv_std_logic_vector(48995, 16),
61390 => conv_std_logic_vector(49234, 16),
61391 => conv_std_logic_vector(49473, 16),
61392 => conv_std_logic_vector(49712, 16),
61393 => conv_std_logic_vector(49951, 16),
61394 => conv_std_logic_vector(50190, 16),
61395 => conv_std_logic_vector(50429, 16),
61396 => conv_std_logic_vector(50668, 16),
61397 => conv_std_logic_vector(50907, 16),
61398 => conv_std_logic_vector(51146, 16),
61399 => conv_std_logic_vector(51385, 16),
61400 => conv_std_logic_vector(51624, 16),
61401 => conv_std_logic_vector(51863, 16),
61402 => conv_std_logic_vector(52102, 16),
61403 => conv_std_logic_vector(52341, 16),
61404 => conv_std_logic_vector(52580, 16),
61405 => conv_std_logic_vector(52819, 16),
61406 => conv_std_logic_vector(53058, 16),
61407 => conv_std_logic_vector(53297, 16),
61408 => conv_std_logic_vector(53536, 16),
61409 => conv_std_logic_vector(53775, 16),
61410 => conv_std_logic_vector(54014, 16),
61411 => conv_std_logic_vector(54253, 16),
61412 => conv_std_logic_vector(54492, 16),
61413 => conv_std_logic_vector(54731, 16),
61414 => conv_std_logic_vector(54970, 16),
61415 => conv_std_logic_vector(55209, 16),
61416 => conv_std_logic_vector(55448, 16),
61417 => conv_std_logic_vector(55687, 16),
61418 => conv_std_logic_vector(55926, 16),
61419 => conv_std_logic_vector(56165, 16),
61420 => conv_std_logic_vector(56404, 16),
61421 => conv_std_logic_vector(56643, 16),
61422 => conv_std_logic_vector(56882, 16),
61423 => conv_std_logic_vector(57121, 16),
61424 => conv_std_logic_vector(57360, 16),
61425 => conv_std_logic_vector(57599, 16),
61426 => conv_std_logic_vector(57838, 16),
61427 => conv_std_logic_vector(58077, 16),
61428 => conv_std_logic_vector(58316, 16),
61429 => conv_std_logic_vector(58555, 16),
61430 => conv_std_logic_vector(58794, 16),
61431 => conv_std_logic_vector(59033, 16),
61432 => conv_std_logic_vector(59272, 16),
61433 => conv_std_logic_vector(59511, 16),
61434 => conv_std_logic_vector(59750, 16),
61435 => conv_std_logic_vector(59989, 16),
61436 => conv_std_logic_vector(60228, 16),
61437 => conv_std_logic_vector(60467, 16),
61438 => conv_std_logic_vector(60706, 16),
61439 => conv_std_logic_vector(60945, 16),
61440 => conv_std_logic_vector(0, 16),
61441 => conv_std_logic_vector(240, 16),
61442 => conv_std_logic_vector(480, 16),
61443 => conv_std_logic_vector(720, 16),
61444 => conv_std_logic_vector(960, 16),
61445 => conv_std_logic_vector(1200, 16),
61446 => conv_std_logic_vector(1440, 16),
61447 => conv_std_logic_vector(1680, 16),
61448 => conv_std_logic_vector(1920, 16),
61449 => conv_std_logic_vector(2160, 16),
61450 => conv_std_logic_vector(2400, 16),
61451 => conv_std_logic_vector(2640, 16),
61452 => conv_std_logic_vector(2880, 16),
61453 => conv_std_logic_vector(3120, 16),
61454 => conv_std_logic_vector(3360, 16),
61455 => conv_std_logic_vector(3600, 16),
61456 => conv_std_logic_vector(3840, 16),
61457 => conv_std_logic_vector(4080, 16),
61458 => conv_std_logic_vector(4320, 16),
61459 => conv_std_logic_vector(4560, 16),
61460 => conv_std_logic_vector(4800, 16),
61461 => conv_std_logic_vector(5040, 16),
61462 => conv_std_logic_vector(5280, 16),
61463 => conv_std_logic_vector(5520, 16),
61464 => conv_std_logic_vector(5760, 16),
61465 => conv_std_logic_vector(6000, 16),
61466 => conv_std_logic_vector(6240, 16),
61467 => conv_std_logic_vector(6480, 16),
61468 => conv_std_logic_vector(6720, 16),
61469 => conv_std_logic_vector(6960, 16),
61470 => conv_std_logic_vector(7200, 16),
61471 => conv_std_logic_vector(7440, 16),
61472 => conv_std_logic_vector(7680, 16),
61473 => conv_std_logic_vector(7920, 16),
61474 => conv_std_logic_vector(8160, 16),
61475 => conv_std_logic_vector(8400, 16),
61476 => conv_std_logic_vector(8640, 16),
61477 => conv_std_logic_vector(8880, 16),
61478 => conv_std_logic_vector(9120, 16),
61479 => conv_std_logic_vector(9360, 16),
61480 => conv_std_logic_vector(9600, 16),
61481 => conv_std_logic_vector(9840, 16),
61482 => conv_std_logic_vector(10080, 16),
61483 => conv_std_logic_vector(10320, 16),
61484 => conv_std_logic_vector(10560, 16),
61485 => conv_std_logic_vector(10800, 16),
61486 => conv_std_logic_vector(11040, 16),
61487 => conv_std_logic_vector(11280, 16),
61488 => conv_std_logic_vector(11520, 16),
61489 => conv_std_logic_vector(11760, 16),
61490 => conv_std_logic_vector(12000, 16),
61491 => conv_std_logic_vector(12240, 16),
61492 => conv_std_logic_vector(12480, 16),
61493 => conv_std_logic_vector(12720, 16),
61494 => conv_std_logic_vector(12960, 16),
61495 => conv_std_logic_vector(13200, 16),
61496 => conv_std_logic_vector(13440, 16),
61497 => conv_std_logic_vector(13680, 16),
61498 => conv_std_logic_vector(13920, 16),
61499 => conv_std_logic_vector(14160, 16),
61500 => conv_std_logic_vector(14400, 16),
61501 => conv_std_logic_vector(14640, 16),
61502 => conv_std_logic_vector(14880, 16),
61503 => conv_std_logic_vector(15120, 16),
61504 => conv_std_logic_vector(15360, 16),
61505 => conv_std_logic_vector(15600, 16),
61506 => conv_std_logic_vector(15840, 16),
61507 => conv_std_logic_vector(16080, 16),
61508 => conv_std_logic_vector(16320, 16),
61509 => conv_std_logic_vector(16560, 16),
61510 => conv_std_logic_vector(16800, 16),
61511 => conv_std_logic_vector(17040, 16),
61512 => conv_std_logic_vector(17280, 16),
61513 => conv_std_logic_vector(17520, 16),
61514 => conv_std_logic_vector(17760, 16),
61515 => conv_std_logic_vector(18000, 16),
61516 => conv_std_logic_vector(18240, 16),
61517 => conv_std_logic_vector(18480, 16),
61518 => conv_std_logic_vector(18720, 16),
61519 => conv_std_logic_vector(18960, 16),
61520 => conv_std_logic_vector(19200, 16),
61521 => conv_std_logic_vector(19440, 16),
61522 => conv_std_logic_vector(19680, 16),
61523 => conv_std_logic_vector(19920, 16),
61524 => conv_std_logic_vector(20160, 16),
61525 => conv_std_logic_vector(20400, 16),
61526 => conv_std_logic_vector(20640, 16),
61527 => conv_std_logic_vector(20880, 16),
61528 => conv_std_logic_vector(21120, 16),
61529 => conv_std_logic_vector(21360, 16),
61530 => conv_std_logic_vector(21600, 16),
61531 => conv_std_logic_vector(21840, 16),
61532 => conv_std_logic_vector(22080, 16),
61533 => conv_std_logic_vector(22320, 16),
61534 => conv_std_logic_vector(22560, 16),
61535 => conv_std_logic_vector(22800, 16),
61536 => conv_std_logic_vector(23040, 16),
61537 => conv_std_logic_vector(23280, 16),
61538 => conv_std_logic_vector(23520, 16),
61539 => conv_std_logic_vector(23760, 16),
61540 => conv_std_logic_vector(24000, 16),
61541 => conv_std_logic_vector(24240, 16),
61542 => conv_std_logic_vector(24480, 16),
61543 => conv_std_logic_vector(24720, 16),
61544 => conv_std_logic_vector(24960, 16),
61545 => conv_std_logic_vector(25200, 16),
61546 => conv_std_logic_vector(25440, 16),
61547 => conv_std_logic_vector(25680, 16),
61548 => conv_std_logic_vector(25920, 16),
61549 => conv_std_logic_vector(26160, 16),
61550 => conv_std_logic_vector(26400, 16),
61551 => conv_std_logic_vector(26640, 16),
61552 => conv_std_logic_vector(26880, 16),
61553 => conv_std_logic_vector(27120, 16),
61554 => conv_std_logic_vector(27360, 16),
61555 => conv_std_logic_vector(27600, 16),
61556 => conv_std_logic_vector(27840, 16),
61557 => conv_std_logic_vector(28080, 16),
61558 => conv_std_logic_vector(28320, 16),
61559 => conv_std_logic_vector(28560, 16),
61560 => conv_std_logic_vector(28800, 16),
61561 => conv_std_logic_vector(29040, 16),
61562 => conv_std_logic_vector(29280, 16),
61563 => conv_std_logic_vector(29520, 16),
61564 => conv_std_logic_vector(29760, 16),
61565 => conv_std_logic_vector(30000, 16),
61566 => conv_std_logic_vector(30240, 16),
61567 => conv_std_logic_vector(30480, 16),
61568 => conv_std_logic_vector(30720, 16),
61569 => conv_std_logic_vector(30960, 16),
61570 => conv_std_logic_vector(31200, 16),
61571 => conv_std_logic_vector(31440, 16),
61572 => conv_std_logic_vector(31680, 16),
61573 => conv_std_logic_vector(31920, 16),
61574 => conv_std_logic_vector(32160, 16),
61575 => conv_std_logic_vector(32400, 16),
61576 => conv_std_logic_vector(32640, 16),
61577 => conv_std_logic_vector(32880, 16),
61578 => conv_std_logic_vector(33120, 16),
61579 => conv_std_logic_vector(33360, 16),
61580 => conv_std_logic_vector(33600, 16),
61581 => conv_std_logic_vector(33840, 16),
61582 => conv_std_logic_vector(34080, 16),
61583 => conv_std_logic_vector(34320, 16),
61584 => conv_std_logic_vector(34560, 16),
61585 => conv_std_logic_vector(34800, 16),
61586 => conv_std_logic_vector(35040, 16),
61587 => conv_std_logic_vector(35280, 16),
61588 => conv_std_logic_vector(35520, 16),
61589 => conv_std_logic_vector(35760, 16),
61590 => conv_std_logic_vector(36000, 16),
61591 => conv_std_logic_vector(36240, 16),
61592 => conv_std_logic_vector(36480, 16),
61593 => conv_std_logic_vector(36720, 16),
61594 => conv_std_logic_vector(36960, 16),
61595 => conv_std_logic_vector(37200, 16),
61596 => conv_std_logic_vector(37440, 16),
61597 => conv_std_logic_vector(37680, 16),
61598 => conv_std_logic_vector(37920, 16),
61599 => conv_std_logic_vector(38160, 16),
61600 => conv_std_logic_vector(38400, 16),
61601 => conv_std_logic_vector(38640, 16),
61602 => conv_std_logic_vector(38880, 16),
61603 => conv_std_logic_vector(39120, 16),
61604 => conv_std_logic_vector(39360, 16),
61605 => conv_std_logic_vector(39600, 16),
61606 => conv_std_logic_vector(39840, 16),
61607 => conv_std_logic_vector(40080, 16),
61608 => conv_std_logic_vector(40320, 16),
61609 => conv_std_logic_vector(40560, 16),
61610 => conv_std_logic_vector(40800, 16),
61611 => conv_std_logic_vector(41040, 16),
61612 => conv_std_logic_vector(41280, 16),
61613 => conv_std_logic_vector(41520, 16),
61614 => conv_std_logic_vector(41760, 16),
61615 => conv_std_logic_vector(42000, 16),
61616 => conv_std_logic_vector(42240, 16),
61617 => conv_std_logic_vector(42480, 16),
61618 => conv_std_logic_vector(42720, 16),
61619 => conv_std_logic_vector(42960, 16),
61620 => conv_std_logic_vector(43200, 16),
61621 => conv_std_logic_vector(43440, 16),
61622 => conv_std_logic_vector(43680, 16),
61623 => conv_std_logic_vector(43920, 16),
61624 => conv_std_logic_vector(44160, 16),
61625 => conv_std_logic_vector(44400, 16),
61626 => conv_std_logic_vector(44640, 16),
61627 => conv_std_logic_vector(44880, 16),
61628 => conv_std_logic_vector(45120, 16),
61629 => conv_std_logic_vector(45360, 16),
61630 => conv_std_logic_vector(45600, 16),
61631 => conv_std_logic_vector(45840, 16),
61632 => conv_std_logic_vector(46080, 16),
61633 => conv_std_logic_vector(46320, 16),
61634 => conv_std_logic_vector(46560, 16),
61635 => conv_std_logic_vector(46800, 16),
61636 => conv_std_logic_vector(47040, 16),
61637 => conv_std_logic_vector(47280, 16),
61638 => conv_std_logic_vector(47520, 16),
61639 => conv_std_logic_vector(47760, 16),
61640 => conv_std_logic_vector(48000, 16),
61641 => conv_std_logic_vector(48240, 16),
61642 => conv_std_logic_vector(48480, 16),
61643 => conv_std_logic_vector(48720, 16),
61644 => conv_std_logic_vector(48960, 16),
61645 => conv_std_logic_vector(49200, 16),
61646 => conv_std_logic_vector(49440, 16),
61647 => conv_std_logic_vector(49680, 16),
61648 => conv_std_logic_vector(49920, 16),
61649 => conv_std_logic_vector(50160, 16),
61650 => conv_std_logic_vector(50400, 16),
61651 => conv_std_logic_vector(50640, 16),
61652 => conv_std_logic_vector(50880, 16),
61653 => conv_std_logic_vector(51120, 16),
61654 => conv_std_logic_vector(51360, 16),
61655 => conv_std_logic_vector(51600, 16),
61656 => conv_std_logic_vector(51840, 16),
61657 => conv_std_logic_vector(52080, 16),
61658 => conv_std_logic_vector(52320, 16),
61659 => conv_std_logic_vector(52560, 16),
61660 => conv_std_logic_vector(52800, 16),
61661 => conv_std_logic_vector(53040, 16),
61662 => conv_std_logic_vector(53280, 16),
61663 => conv_std_logic_vector(53520, 16),
61664 => conv_std_logic_vector(53760, 16),
61665 => conv_std_logic_vector(54000, 16),
61666 => conv_std_logic_vector(54240, 16),
61667 => conv_std_logic_vector(54480, 16),
61668 => conv_std_logic_vector(54720, 16),
61669 => conv_std_logic_vector(54960, 16),
61670 => conv_std_logic_vector(55200, 16),
61671 => conv_std_logic_vector(55440, 16),
61672 => conv_std_logic_vector(55680, 16),
61673 => conv_std_logic_vector(55920, 16),
61674 => conv_std_logic_vector(56160, 16),
61675 => conv_std_logic_vector(56400, 16),
61676 => conv_std_logic_vector(56640, 16),
61677 => conv_std_logic_vector(56880, 16),
61678 => conv_std_logic_vector(57120, 16),
61679 => conv_std_logic_vector(57360, 16),
61680 => conv_std_logic_vector(57600, 16),
61681 => conv_std_logic_vector(57840, 16),
61682 => conv_std_logic_vector(58080, 16),
61683 => conv_std_logic_vector(58320, 16),
61684 => conv_std_logic_vector(58560, 16),
61685 => conv_std_logic_vector(58800, 16),
61686 => conv_std_logic_vector(59040, 16),
61687 => conv_std_logic_vector(59280, 16),
61688 => conv_std_logic_vector(59520, 16),
61689 => conv_std_logic_vector(59760, 16),
61690 => conv_std_logic_vector(60000, 16),
61691 => conv_std_logic_vector(60240, 16),
61692 => conv_std_logic_vector(60480, 16),
61693 => conv_std_logic_vector(60720, 16),
61694 => conv_std_logic_vector(60960, 16),
61695 => conv_std_logic_vector(61200, 16),
61696 => conv_std_logic_vector(0, 16),
61697 => conv_std_logic_vector(241, 16),
61698 => conv_std_logic_vector(482, 16),
61699 => conv_std_logic_vector(723, 16),
61700 => conv_std_logic_vector(964, 16),
61701 => conv_std_logic_vector(1205, 16),
61702 => conv_std_logic_vector(1446, 16),
61703 => conv_std_logic_vector(1687, 16),
61704 => conv_std_logic_vector(1928, 16),
61705 => conv_std_logic_vector(2169, 16),
61706 => conv_std_logic_vector(2410, 16),
61707 => conv_std_logic_vector(2651, 16),
61708 => conv_std_logic_vector(2892, 16),
61709 => conv_std_logic_vector(3133, 16),
61710 => conv_std_logic_vector(3374, 16),
61711 => conv_std_logic_vector(3615, 16),
61712 => conv_std_logic_vector(3856, 16),
61713 => conv_std_logic_vector(4097, 16),
61714 => conv_std_logic_vector(4338, 16),
61715 => conv_std_logic_vector(4579, 16),
61716 => conv_std_logic_vector(4820, 16),
61717 => conv_std_logic_vector(5061, 16),
61718 => conv_std_logic_vector(5302, 16),
61719 => conv_std_logic_vector(5543, 16),
61720 => conv_std_logic_vector(5784, 16),
61721 => conv_std_logic_vector(6025, 16),
61722 => conv_std_logic_vector(6266, 16),
61723 => conv_std_logic_vector(6507, 16),
61724 => conv_std_logic_vector(6748, 16),
61725 => conv_std_logic_vector(6989, 16),
61726 => conv_std_logic_vector(7230, 16),
61727 => conv_std_logic_vector(7471, 16),
61728 => conv_std_logic_vector(7712, 16),
61729 => conv_std_logic_vector(7953, 16),
61730 => conv_std_logic_vector(8194, 16),
61731 => conv_std_logic_vector(8435, 16),
61732 => conv_std_logic_vector(8676, 16),
61733 => conv_std_logic_vector(8917, 16),
61734 => conv_std_logic_vector(9158, 16),
61735 => conv_std_logic_vector(9399, 16),
61736 => conv_std_logic_vector(9640, 16),
61737 => conv_std_logic_vector(9881, 16),
61738 => conv_std_logic_vector(10122, 16),
61739 => conv_std_logic_vector(10363, 16),
61740 => conv_std_logic_vector(10604, 16),
61741 => conv_std_logic_vector(10845, 16),
61742 => conv_std_logic_vector(11086, 16),
61743 => conv_std_logic_vector(11327, 16),
61744 => conv_std_logic_vector(11568, 16),
61745 => conv_std_logic_vector(11809, 16),
61746 => conv_std_logic_vector(12050, 16),
61747 => conv_std_logic_vector(12291, 16),
61748 => conv_std_logic_vector(12532, 16),
61749 => conv_std_logic_vector(12773, 16),
61750 => conv_std_logic_vector(13014, 16),
61751 => conv_std_logic_vector(13255, 16),
61752 => conv_std_logic_vector(13496, 16),
61753 => conv_std_logic_vector(13737, 16),
61754 => conv_std_logic_vector(13978, 16),
61755 => conv_std_logic_vector(14219, 16),
61756 => conv_std_logic_vector(14460, 16),
61757 => conv_std_logic_vector(14701, 16),
61758 => conv_std_logic_vector(14942, 16),
61759 => conv_std_logic_vector(15183, 16),
61760 => conv_std_logic_vector(15424, 16),
61761 => conv_std_logic_vector(15665, 16),
61762 => conv_std_logic_vector(15906, 16),
61763 => conv_std_logic_vector(16147, 16),
61764 => conv_std_logic_vector(16388, 16),
61765 => conv_std_logic_vector(16629, 16),
61766 => conv_std_logic_vector(16870, 16),
61767 => conv_std_logic_vector(17111, 16),
61768 => conv_std_logic_vector(17352, 16),
61769 => conv_std_logic_vector(17593, 16),
61770 => conv_std_logic_vector(17834, 16),
61771 => conv_std_logic_vector(18075, 16),
61772 => conv_std_logic_vector(18316, 16),
61773 => conv_std_logic_vector(18557, 16),
61774 => conv_std_logic_vector(18798, 16),
61775 => conv_std_logic_vector(19039, 16),
61776 => conv_std_logic_vector(19280, 16),
61777 => conv_std_logic_vector(19521, 16),
61778 => conv_std_logic_vector(19762, 16),
61779 => conv_std_logic_vector(20003, 16),
61780 => conv_std_logic_vector(20244, 16),
61781 => conv_std_logic_vector(20485, 16),
61782 => conv_std_logic_vector(20726, 16),
61783 => conv_std_logic_vector(20967, 16),
61784 => conv_std_logic_vector(21208, 16),
61785 => conv_std_logic_vector(21449, 16),
61786 => conv_std_logic_vector(21690, 16),
61787 => conv_std_logic_vector(21931, 16),
61788 => conv_std_logic_vector(22172, 16),
61789 => conv_std_logic_vector(22413, 16),
61790 => conv_std_logic_vector(22654, 16),
61791 => conv_std_logic_vector(22895, 16),
61792 => conv_std_logic_vector(23136, 16),
61793 => conv_std_logic_vector(23377, 16),
61794 => conv_std_logic_vector(23618, 16),
61795 => conv_std_logic_vector(23859, 16),
61796 => conv_std_logic_vector(24100, 16),
61797 => conv_std_logic_vector(24341, 16),
61798 => conv_std_logic_vector(24582, 16),
61799 => conv_std_logic_vector(24823, 16),
61800 => conv_std_logic_vector(25064, 16),
61801 => conv_std_logic_vector(25305, 16),
61802 => conv_std_logic_vector(25546, 16),
61803 => conv_std_logic_vector(25787, 16),
61804 => conv_std_logic_vector(26028, 16),
61805 => conv_std_logic_vector(26269, 16),
61806 => conv_std_logic_vector(26510, 16),
61807 => conv_std_logic_vector(26751, 16),
61808 => conv_std_logic_vector(26992, 16),
61809 => conv_std_logic_vector(27233, 16),
61810 => conv_std_logic_vector(27474, 16),
61811 => conv_std_logic_vector(27715, 16),
61812 => conv_std_logic_vector(27956, 16),
61813 => conv_std_logic_vector(28197, 16),
61814 => conv_std_logic_vector(28438, 16),
61815 => conv_std_logic_vector(28679, 16),
61816 => conv_std_logic_vector(28920, 16),
61817 => conv_std_logic_vector(29161, 16),
61818 => conv_std_logic_vector(29402, 16),
61819 => conv_std_logic_vector(29643, 16),
61820 => conv_std_logic_vector(29884, 16),
61821 => conv_std_logic_vector(30125, 16),
61822 => conv_std_logic_vector(30366, 16),
61823 => conv_std_logic_vector(30607, 16),
61824 => conv_std_logic_vector(30848, 16),
61825 => conv_std_logic_vector(31089, 16),
61826 => conv_std_logic_vector(31330, 16),
61827 => conv_std_logic_vector(31571, 16),
61828 => conv_std_logic_vector(31812, 16),
61829 => conv_std_logic_vector(32053, 16),
61830 => conv_std_logic_vector(32294, 16),
61831 => conv_std_logic_vector(32535, 16),
61832 => conv_std_logic_vector(32776, 16),
61833 => conv_std_logic_vector(33017, 16),
61834 => conv_std_logic_vector(33258, 16),
61835 => conv_std_logic_vector(33499, 16),
61836 => conv_std_logic_vector(33740, 16),
61837 => conv_std_logic_vector(33981, 16),
61838 => conv_std_logic_vector(34222, 16),
61839 => conv_std_logic_vector(34463, 16),
61840 => conv_std_logic_vector(34704, 16),
61841 => conv_std_logic_vector(34945, 16),
61842 => conv_std_logic_vector(35186, 16),
61843 => conv_std_logic_vector(35427, 16),
61844 => conv_std_logic_vector(35668, 16),
61845 => conv_std_logic_vector(35909, 16),
61846 => conv_std_logic_vector(36150, 16),
61847 => conv_std_logic_vector(36391, 16),
61848 => conv_std_logic_vector(36632, 16),
61849 => conv_std_logic_vector(36873, 16),
61850 => conv_std_logic_vector(37114, 16),
61851 => conv_std_logic_vector(37355, 16),
61852 => conv_std_logic_vector(37596, 16),
61853 => conv_std_logic_vector(37837, 16),
61854 => conv_std_logic_vector(38078, 16),
61855 => conv_std_logic_vector(38319, 16),
61856 => conv_std_logic_vector(38560, 16),
61857 => conv_std_logic_vector(38801, 16),
61858 => conv_std_logic_vector(39042, 16),
61859 => conv_std_logic_vector(39283, 16),
61860 => conv_std_logic_vector(39524, 16),
61861 => conv_std_logic_vector(39765, 16),
61862 => conv_std_logic_vector(40006, 16),
61863 => conv_std_logic_vector(40247, 16),
61864 => conv_std_logic_vector(40488, 16),
61865 => conv_std_logic_vector(40729, 16),
61866 => conv_std_logic_vector(40970, 16),
61867 => conv_std_logic_vector(41211, 16),
61868 => conv_std_logic_vector(41452, 16),
61869 => conv_std_logic_vector(41693, 16),
61870 => conv_std_logic_vector(41934, 16),
61871 => conv_std_logic_vector(42175, 16),
61872 => conv_std_logic_vector(42416, 16),
61873 => conv_std_logic_vector(42657, 16),
61874 => conv_std_logic_vector(42898, 16),
61875 => conv_std_logic_vector(43139, 16),
61876 => conv_std_logic_vector(43380, 16),
61877 => conv_std_logic_vector(43621, 16),
61878 => conv_std_logic_vector(43862, 16),
61879 => conv_std_logic_vector(44103, 16),
61880 => conv_std_logic_vector(44344, 16),
61881 => conv_std_logic_vector(44585, 16),
61882 => conv_std_logic_vector(44826, 16),
61883 => conv_std_logic_vector(45067, 16),
61884 => conv_std_logic_vector(45308, 16),
61885 => conv_std_logic_vector(45549, 16),
61886 => conv_std_logic_vector(45790, 16),
61887 => conv_std_logic_vector(46031, 16),
61888 => conv_std_logic_vector(46272, 16),
61889 => conv_std_logic_vector(46513, 16),
61890 => conv_std_logic_vector(46754, 16),
61891 => conv_std_logic_vector(46995, 16),
61892 => conv_std_logic_vector(47236, 16),
61893 => conv_std_logic_vector(47477, 16),
61894 => conv_std_logic_vector(47718, 16),
61895 => conv_std_logic_vector(47959, 16),
61896 => conv_std_logic_vector(48200, 16),
61897 => conv_std_logic_vector(48441, 16),
61898 => conv_std_logic_vector(48682, 16),
61899 => conv_std_logic_vector(48923, 16),
61900 => conv_std_logic_vector(49164, 16),
61901 => conv_std_logic_vector(49405, 16),
61902 => conv_std_logic_vector(49646, 16),
61903 => conv_std_logic_vector(49887, 16),
61904 => conv_std_logic_vector(50128, 16),
61905 => conv_std_logic_vector(50369, 16),
61906 => conv_std_logic_vector(50610, 16),
61907 => conv_std_logic_vector(50851, 16),
61908 => conv_std_logic_vector(51092, 16),
61909 => conv_std_logic_vector(51333, 16),
61910 => conv_std_logic_vector(51574, 16),
61911 => conv_std_logic_vector(51815, 16),
61912 => conv_std_logic_vector(52056, 16),
61913 => conv_std_logic_vector(52297, 16),
61914 => conv_std_logic_vector(52538, 16),
61915 => conv_std_logic_vector(52779, 16),
61916 => conv_std_logic_vector(53020, 16),
61917 => conv_std_logic_vector(53261, 16),
61918 => conv_std_logic_vector(53502, 16),
61919 => conv_std_logic_vector(53743, 16),
61920 => conv_std_logic_vector(53984, 16),
61921 => conv_std_logic_vector(54225, 16),
61922 => conv_std_logic_vector(54466, 16),
61923 => conv_std_logic_vector(54707, 16),
61924 => conv_std_logic_vector(54948, 16),
61925 => conv_std_logic_vector(55189, 16),
61926 => conv_std_logic_vector(55430, 16),
61927 => conv_std_logic_vector(55671, 16),
61928 => conv_std_logic_vector(55912, 16),
61929 => conv_std_logic_vector(56153, 16),
61930 => conv_std_logic_vector(56394, 16),
61931 => conv_std_logic_vector(56635, 16),
61932 => conv_std_logic_vector(56876, 16),
61933 => conv_std_logic_vector(57117, 16),
61934 => conv_std_logic_vector(57358, 16),
61935 => conv_std_logic_vector(57599, 16),
61936 => conv_std_logic_vector(57840, 16),
61937 => conv_std_logic_vector(58081, 16),
61938 => conv_std_logic_vector(58322, 16),
61939 => conv_std_logic_vector(58563, 16),
61940 => conv_std_logic_vector(58804, 16),
61941 => conv_std_logic_vector(59045, 16),
61942 => conv_std_logic_vector(59286, 16),
61943 => conv_std_logic_vector(59527, 16),
61944 => conv_std_logic_vector(59768, 16),
61945 => conv_std_logic_vector(60009, 16),
61946 => conv_std_logic_vector(60250, 16),
61947 => conv_std_logic_vector(60491, 16),
61948 => conv_std_logic_vector(60732, 16),
61949 => conv_std_logic_vector(60973, 16),
61950 => conv_std_logic_vector(61214, 16),
61951 => conv_std_logic_vector(61455, 16),
61952 => conv_std_logic_vector(0, 16),
61953 => conv_std_logic_vector(242, 16),
61954 => conv_std_logic_vector(484, 16),
61955 => conv_std_logic_vector(726, 16),
61956 => conv_std_logic_vector(968, 16),
61957 => conv_std_logic_vector(1210, 16),
61958 => conv_std_logic_vector(1452, 16),
61959 => conv_std_logic_vector(1694, 16),
61960 => conv_std_logic_vector(1936, 16),
61961 => conv_std_logic_vector(2178, 16),
61962 => conv_std_logic_vector(2420, 16),
61963 => conv_std_logic_vector(2662, 16),
61964 => conv_std_logic_vector(2904, 16),
61965 => conv_std_logic_vector(3146, 16),
61966 => conv_std_logic_vector(3388, 16),
61967 => conv_std_logic_vector(3630, 16),
61968 => conv_std_logic_vector(3872, 16),
61969 => conv_std_logic_vector(4114, 16),
61970 => conv_std_logic_vector(4356, 16),
61971 => conv_std_logic_vector(4598, 16),
61972 => conv_std_logic_vector(4840, 16),
61973 => conv_std_logic_vector(5082, 16),
61974 => conv_std_logic_vector(5324, 16),
61975 => conv_std_logic_vector(5566, 16),
61976 => conv_std_logic_vector(5808, 16),
61977 => conv_std_logic_vector(6050, 16),
61978 => conv_std_logic_vector(6292, 16),
61979 => conv_std_logic_vector(6534, 16),
61980 => conv_std_logic_vector(6776, 16),
61981 => conv_std_logic_vector(7018, 16),
61982 => conv_std_logic_vector(7260, 16),
61983 => conv_std_logic_vector(7502, 16),
61984 => conv_std_logic_vector(7744, 16),
61985 => conv_std_logic_vector(7986, 16),
61986 => conv_std_logic_vector(8228, 16),
61987 => conv_std_logic_vector(8470, 16),
61988 => conv_std_logic_vector(8712, 16),
61989 => conv_std_logic_vector(8954, 16),
61990 => conv_std_logic_vector(9196, 16),
61991 => conv_std_logic_vector(9438, 16),
61992 => conv_std_logic_vector(9680, 16),
61993 => conv_std_logic_vector(9922, 16),
61994 => conv_std_logic_vector(10164, 16),
61995 => conv_std_logic_vector(10406, 16),
61996 => conv_std_logic_vector(10648, 16),
61997 => conv_std_logic_vector(10890, 16),
61998 => conv_std_logic_vector(11132, 16),
61999 => conv_std_logic_vector(11374, 16),
62000 => conv_std_logic_vector(11616, 16),
62001 => conv_std_logic_vector(11858, 16),
62002 => conv_std_logic_vector(12100, 16),
62003 => conv_std_logic_vector(12342, 16),
62004 => conv_std_logic_vector(12584, 16),
62005 => conv_std_logic_vector(12826, 16),
62006 => conv_std_logic_vector(13068, 16),
62007 => conv_std_logic_vector(13310, 16),
62008 => conv_std_logic_vector(13552, 16),
62009 => conv_std_logic_vector(13794, 16),
62010 => conv_std_logic_vector(14036, 16),
62011 => conv_std_logic_vector(14278, 16),
62012 => conv_std_logic_vector(14520, 16),
62013 => conv_std_logic_vector(14762, 16),
62014 => conv_std_logic_vector(15004, 16),
62015 => conv_std_logic_vector(15246, 16),
62016 => conv_std_logic_vector(15488, 16),
62017 => conv_std_logic_vector(15730, 16),
62018 => conv_std_logic_vector(15972, 16),
62019 => conv_std_logic_vector(16214, 16),
62020 => conv_std_logic_vector(16456, 16),
62021 => conv_std_logic_vector(16698, 16),
62022 => conv_std_logic_vector(16940, 16),
62023 => conv_std_logic_vector(17182, 16),
62024 => conv_std_logic_vector(17424, 16),
62025 => conv_std_logic_vector(17666, 16),
62026 => conv_std_logic_vector(17908, 16),
62027 => conv_std_logic_vector(18150, 16),
62028 => conv_std_logic_vector(18392, 16),
62029 => conv_std_logic_vector(18634, 16),
62030 => conv_std_logic_vector(18876, 16),
62031 => conv_std_logic_vector(19118, 16),
62032 => conv_std_logic_vector(19360, 16),
62033 => conv_std_logic_vector(19602, 16),
62034 => conv_std_logic_vector(19844, 16),
62035 => conv_std_logic_vector(20086, 16),
62036 => conv_std_logic_vector(20328, 16),
62037 => conv_std_logic_vector(20570, 16),
62038 => conv_std_logic_vector(20812, 16),
62039 => conv_std_logic_vector(21054, 16),
62040 => conv_std_logic_vector(21296, 16),
62041 => conv_std_logic_vector(21538, 16),
62042 => conv_std_logic_vector(21780, 16),
62043 => conv_std_logic_vector(22022, 16),
62044 => conv_std_logic_vector(22264, 16),
62045 => conv_std_logic_vector(22506, 16),
62046 => conv_std_logic_vector(22748, 16),
62047 => conv_std_logic_vector(22990, 16),
62048 => conv_std_logic_vector(23232, 16),
62049 => conv_std_logic_vector(23474, 16),
62050 => conv_std_logic_vector(23716, 16),
62051 => conv_std_logic_vector(23958, 16),
62052 => conv_std_logic_vector(24200, 16),
62053 => conv_std_logic_vector(24442, 16),
62054 => conv_std_logic_vector(24684, 16),
62055 => conv_std_logic_vector(24926, 16),
62056 => conv_std_logic_vector(25168, 16),
62057 => conv_std_logic_vector(25410, 16),
62058 => conv_std_logic_vector(25652, 16),
62059 => conv_std_logic_vector(25894, 16),
62060 => conv_std_logic_vector(26136, 16),
62061 => conv_std_logic_vector(26378, 16),
62062 => conv_std_logic_vector(26620, 16),
62063 => conv_std_logic_vector(26862, 16),
62064 => conv_std_logic_vector(27104, 16),
62065 => conv_std_logic_vector(27346, 16),
62066 => conv_std_logic_vector(27588, 16),
62067 => conv_std_logic_vector(27830, 16),
62068 => conv_std_logic_vector(28072, 16),
62069 => conv_std_logic_vector(28314, 16),
62070 => conv_std_logic_vector(28556, 16),
62071 => conv_std_logic_vector(28798, 16),
62072 => conv_std_logic_vector(29040, 16),
62073 => conv_std_logic_vector(29282, 16),
62074 => conv_std_logic_vector(29524, 16),
62075 => conv_std_logic_vector(29766, 16),
62076 => conv_std_logic_vector(30008, 16),
62077 => conv_std_logic_vector(30250, 16),
62078 => conv_std_logic_vector(30492, 16),
62079 => conv_std_logic_vector(30734, 16),
62080 => conv_std_logic_vector(30976, 16),
62081 => conv_std_logic_vector(31218, 16),
62082 => conv_std_logic_vector(31460, 16),
62083 => conv_std_logic_vector(31702, 16),
62084 => conv_std_logic_vector(31944, 16),
62085 => conv_std_logic_vector(32186, 16),
62086 => conv_std_logic_vector(32428, 16),
62087 => conv_std_logic_vector(32670, 16),
62088 => conv_std_logic_vector(32912, 16),
62089 => conv_std_logic_vector(33154, 16),
62090 => conv_std_logic_vector(33396, 16),
62091 => conv_std_logic_vector(33638, 16),
62092 => conv_std_logic_vector(33880, 16),
62093 => conv_std_logic_vector(34122, 16),
62094 => conv_std_logic_vector(34364, 16),
62095 => conv_std_logic_vector(34606, 16),
62096 => conv_std_logic_vector(34848, 16),
62097 => conv_std_logic_vector(35090, 16),
62098 => conv_std_logic_vector(35332, 16),
62099 => conv_std_logic_vector(35574, 16),
62100 => conv_std_logic_vector(35816, 16),
62101 => conv_std_logic_vector(36058, 16),
62102 => conv_std_logic_vector(36300, 16),
62103 => conv_std_logic_vector(36542, 16),
62104 => conv_std_logic_vector(36784, 16),
62105 => conv_std_logic_vector(37026, 16),
62106 => conv_std_logic_vector(37268, 16),
62107 => conv_std_logic_vector(37510, 16),
62108 => conv_std_logic_vector(37752, 16),
62109 => conv_std_logic_vector(37994, 16),
62110 => conv_std_logic_vector(38236, 16),
62111 => conv_std_logic_vector(38478, 16),
62112 => conv_std_logic_vector(38720, 16),
62113 => conv_std_logic_vector(38962, 16),
62114 => conv_std_logic_vector(39204, 16),
62115 => conv_std_logic_vector(39446, 16),
62116 => conv_std_logic_vector(39688, 16),
62117 => conv_std_logic_vector(39930, 16),
62118 => conv_std_logic_vector(40172, 16),
62119 => conv_std_logic_vector(40414, 16),
62120 => conv_std_logic_vector(40656, 16),
62121 => conv_std_logic_vector(40898, 16),
62122 => conv_std_logic_vector(41140, 16),
62123 => conv_std_logic_vector(41382, 16),
62124 => conv_std_logic_vector(41624, 16),
62125 => conv_std_logic_vector(41866, 16),
62126 => conv_std_logic_vector(42108, 16),
62127 => conv_std_logic_vector(42350, 16),
62128 => conv_std_logic_vector(42592, 16),
62129 => conv_std_logic_vector(42834, 16),
62130 => conv_std_logic_vector(43076, 16),
62131 => conv_std_logic_vector(43318, 16),
62132 => conv_std_logic_vector(43560, 16),
62133 => conv_std_logic_vector(43802, 16),
62134 => conv_std_logic_vector(44044, 16),
62135 => conv_std_logic_vector(44286, 16),
62136 => conv_std_logic_vector(44528, 16),
62137 => conv_std_logic_vector(44770, 16),
62138 => conv_std_logic_vector(45012, 16),
62139 => conv_std_logic_vector(45254, 16),
62140 => conv_std_logic_vector(45496, 16),
62141 => conv_std_logic_vector(45738, 16),
62142 => conv_std_logic_vector(45980, 16),
62143 => conv_std_logic_vector(46222, 16),
62144 => conv_std_logic_vector(46464, 16),
62145 => conv_std_logic_vector(46706, 16),
62146 => conv_std_logic_vector(46948, 16),
62147 => conv_std_logic_vector(47190, 16),
62148 => conv_std_logic_vector(47432, 16),
62149 => conv_std_logic_vector(47674, 16),
62150 => conv_std_logic_vector(47916, 16),
62151 => conv_std_logic_vector(48158, 16),
62152 => conv_std_logic_vector(48400, 16),
62153 => conv_std_logic_vector(48642, 16),
62154 => conv_std_logic_vector(48884, 16),
62155 => conv_std_logic_vector(49126, 16),
62156 => conv_std_logic_vector(49368, 16),
62157 => conv_std_logic_vector(49610, 16),
62158 => conv_std_logic_vector(49852, 16),
62159 => conv_std_logic_vector(50094, 16),
62160 => conv_std_logic_vector(50336, 16),
62161 => conv_std_logic_vector(50578, 16),
62162 => conv_std_logic_vector(50820, 16),
62163 => conv_std_logic_vector(51062, 16),
62164 => conv_std_logic_vector(51304, 16),
62165 => conv_std_logic_vector(51546, 16),
62166 => conv_std_logic_vector(51788, 16),
62167 => conv_std_logic_vector(52030, 16),
62168 => conv_std_logic_vector(52272, 16),
62169 => conv_std_logic_vector(52514, 16),
62170 => conv_std_logic_vector(52756, 16),
62171 => conv_std_logic_vector(52998, 16),
62172 => conv_std_logic_vector(53240, 16),
62173 => conv_std_logic_vector(53482, 16),
62174 => conv_std_logic_vector(53724, 16),
62175 => conv_std_logic_vector(53966, 16),
62176 => conv_std_logic_vector(54208, 16),
62177 => conv_std_logic_vector(54450, 16),
62178 => conv_std_logic_vector(54692, 16),
62179 => conv_std_logic_vector(54934, 16),
62180 => conv_std_logic_vector(55176, 16),
62181 => conv_std_logic_vector(55418, 16),
62182 => conv_std_logic_vector(55660, 16),
62183 => conv_std_logic_vector(55902, 16),
62184 => conv_std_logic_vector(56144, 16),
62185 => conv_std_logic_vector(56386, 16),
62186 => conv_std_logic_vector(56628, 16),
62187 => conv_std_logic_vector(56870, 16),
62188 => conv_std_logic_vector(57112, 16),
62189 => conv_std_logic_vector(57354, 16),
62190 => conv_std_logic_vector(57596, 16),
62191 => conv_std_logic_vector(57838, 16),
62192 => conv_std_logic_vector(58080, 16),
62193 => conv_std_logic_vector(58322, 16),
62194 => conv_std_logic_vector(58564, 16),
62195 => conv_std_logic_vector(58806, 16),
62196 => conv_std_logic_vector(59048, 16),
62197 => conv_std_logic_vector(59290, 16),
62198 => conv_std_logic_vector(59532, 16),
62199 => conv_std_logic_vector(59774, 16),
62200 => conv_std_logic_vector(60016, 16),
62201 => conv_std_logic_vector(60258, 16),
62202 => conv_std_logic_vector(60500, 16),
62203 => conv_std_logic_vector(60742, 16),
62204 => conv_std_logic_vector(60984, 16),
62205 => conv_std_logic_vector(61226, 16),
62206 => conv_std_logic_vector(61468, 16),
62207 => conv_std_logic_vector(61710, 16),
62208 => conv_std_logic_vector(0, 16),
62209 => conv_std_logic_vector(243, 16),
62210 => conv_std_logic_vector(486, 16),
62211 => conv_std_logic_vector(729, 16),
62212 => conv_std_logic_vector(972, 16),
62213 => conv_std_logic_vector(1215, 16),
62214 => conv_std_logic_vector(1458, 16),
62215 => conv_std_logic_vector(1701, 16),
62216 => conv_std_logic_vector(1944, 16),
62217 => conv_std_logic_vector(2187, 16),
62218 => conv_std_logic_vector(2430, 16),
62219 => conv_std_logic_vector(2673, 16),
62220 => conv_std_logic_vector(2916, 16),
62221 => conv_std_logic_vector(3159, 16),
62222 => conv_std_logic_vector(3402, 16),
62223 => conv_std_logic_vector(3645, 16),
62224 => conv_std_logic_vector(3888, 16),
62225 => conv_std_logic_vector(4131, 16),
62226 => conv_std_logic_vector(4374, 16),
62227 => conv_std_logic_vector(4617, 16),
62228 => conv_std_logic_vector(4860, 16),
62229 => conv_std_logic_vector(5103, 16),
62230 => conv_std_logic_vector(5346, 16),
62231 => conv_std_logic_vector(5589, 16),
62232 => conv_std_logic_vector(5832, 16),
62233 => conv_std_logic_vector(6075, 16),
62234 => conv_std_logic_vector(6318, 16),
62235 => conv_std_logic_vector(6561, 16),
62236 => conv_std_logic_vector(6804, 16),
62237 => conv_std_logic_vector(7047, 16),
62238 => conv_std_logic_vector(7290, 16),
62239 => conv_std_logic_vector(7533, 16),
62240 => conv_std_logic_vector(7776, 16),
62241 => conv_std_logic_vector(8019, 16),
62242 => conv_std_logic_vector(8262, 16),
62243 => conv_std_logic_vector(8505, 16),
62244 => conv_std_logic_vector(8748, 16),
62245 => conv_std_logic_vector(8991, 16),
62246 => conv_std_logic_vector(9234, 16),
62247 => conv_std_logic_vector(9477, 16),
62248 => conv_std_logic_vector(9720, 16),
62249 => conv_std_logic_vector(9963, 16),
62250 => conv_std_logic_vector(10206, 16),
62251 => conv_std_logic_vector(10449, 16),
62252 => conv_std_logic_vector(10692, 16),
62253 => conv_std_logic_vector(10935, 16),
62254 => conv_std_logic_vector(11178, 16),
62255 => conv_std_logic_vector(11421, 16),
62256 => conv_std_logic_vector(11664, 16),
62257 => conv_std_logic_vector(11907, 16),
62258 => conv_std_logic_vector(12150, 16),
62259 => conv_std_logic_vector(12393, 16),
62260 => conv_std_logic_vector(12636, 16),
62261 => conv_std_logic_vector(12879, 16),
62262 => conv_std_logic_vector(13122, 16),
62263 => conv_std_logic_vector(13365, 16),
62264 => conv_std_logic_vector(13608, 16),
62265 => conv_std_logic_vector(13851, 16),
62266 => conv_std_logic_vector(14094, 16),
62267 => conv_std_logic_vector(14337, 16),
62268 => conv_std_logic_vector(14580, 16),
62269 => conv_std_logic_vector(14823, 16),
62270 => conv_std_logic_vector(15066, 16),
62271 => conv_std_logic_vector(15309, 16),
62272 => conv_std_logic_vector(15552, 16),
62273 => conv_std_logic_vector(15795, 16),
62274 => conv_std_logic_vector(16038, 16),
62275 => conv_std_logic_vector(16281, 16),
62276 => conv_std_logic_vector(16524, 16),
62277 => conv_std_logic_vector(16767, 16),
62278 => conv_std_logic_vector(17010, 16),
62279 => conv_std_logic_vector(17253, 16),
62280 => conv_std_logic_vector(17496, 16),
62281 => conv_std_logic_vector(17739, 16),
62282 => conv_std_logic_vector(17982, 16),
62283 => conv_std_logic_vector(18225, 16),
62284 => conv_std_logic_vector(18468, 16),
62285 => conv_std_logic_vector(18711, 16),
62286 => conv_std_logic_vector(18954, 16),
62287 => conv_std_logic_vector(19197, 16),
62288 => conv_std_logic_vector(19440, 16),
62289 => conv_std_logic_vector(19683, 16),
62290 => conv_std_logic_vector(19926, 16),
62291 => conv_std_logic_vector(20169, 16),
62292 => conv_std_logic_vector(20412, 16),
62293 => conv_std_logic_vector(20655, 16),
62294 => conv_std_logic_vector(20898, 16),
62295 => conv_std_logic_vector(21141, 16),
62296 => conv_std_logic_vector(21384, 16),
62297 => conv_std_logic_vector(21627, 16),
62298 => conv_std_logic_vector(21870, 16),
62299 => conv_std_logic_vector(22113, 16),
62300 => conv_std_logic_vector(22356, 16),
62301 => conv_std_logic_vector(22599, 16),
62302 => conv_std_logic_vector(22842, 16),
62303 => conv_std_logic_vector(23085, 16),
62304 => conv_std_logic_vector(23328, 16),
62305 => conv_std_logic_vector(23571, 16),
62306 => conv_std_logic_vector(23814, 16),
62307 => conv_std_logic_vector(24057, 16),
62308 => conv_std_logic_vector(24300, 16),
62309 => conv_std_logic_vector(24543, 16),
62310 => conv_std_logic_vector(24786, 16),
62311 => conv_std_logic_vector(25029, 16),
62312 => conv_std_logic_vector(25272, 16),
62313 => conv_std_logic_vector(25515, 16),
62314 => conv_std_logic_vector(25758, 16),
62315 => conv_std_logic_vector(26001, 16),
62316 => conv_std_logic_vector(26244, 16),
62317 => conv_std_logic_vector(26487, 16),
62318 => conv_std_logic_vector(26730, 16),
62319 => conv_std_logic_vector(26973, 16),
62320 => conv_std_logic_vector(27216, 16),
62321 => conv_std_logic_vector(27459, 16),
62322 => conv_std_logic_vector(27702, 16),
62323 => conv_std_logic_vector(27945, 16),
62324 => conv_std_logic_vector(28188, 16),
62325 => conv_std_logic_vector(28431, 16),
62326 => conv_std_logic_vector(28674, 16),
62327 => conv_std_logic_vector(28917, 16),
62328 => conv_std_logic_vector(29160, 16),
62329 => conv_std_logic_vector(29403, 16),
62330 => conv_std_logic_vector(29646, 16),
62331 => conv_std_logic_vector(29889, 16),
62332 => conv_std_logic_vector(30132, 16),
62333 => conv_std_logic_vector(30375, 16),
62334 => conv_std_logic_vector(30618, 16),
62335 => conv_std_logic_vector(30861, 16),
62336 => conv_std_logic_vector(31104, 16),
62337 => conv_std_logic_vector(31347, 16),
62338 => conv_std_logic_vector(31590, 16),
62339 => conv_std_logic_vector(31833, 16),
62340 => conv_std_logic_vector(32076, 16),
62341 => conv_std_logic_vector(32319, 16),
62342 => conv_std_logic_vector(32562, 16),
62343 => conv_std_logic_vector(32805, 16),
62344 => conv_std_logic_vector(33048, 16),
62345 => conv_std_logic_vector(33291, 16),
62346 => conv_std_logic_vector(33534, 16),
62347 => conv_std_logic_vector(33777, 16),
62348 => conv_std_logic_vector(34020, 16),
62349 => conv_std_logic_vector(34263, 16),
62350 => conv_std_logic_vector(34506, 16),
62351 => conv_std_logic_vector(34749, 16),
62352 => conv_std_logic_vector(34992, 16),
62353 => conv_std_logic_vector(35235, 16),
62354 => conv_std_logic_vector(35478, 16),
62355 => conv_std_logic_vector(35721, 16),
62356 => conv_std_logic_vector(35964, 16),
62357 => conv_std_logic_vector(36207, 16),
62358 => conv_std_logic_vector(36450, 16),
62359 => conv_std_logic_vector(36693, 16),
62360 => conv_std_logic_vector(36936, 16),
62361 => conv_std_logic_vector(37179, 16),
62362 => conv_std_logic_vector(37422, 16),
62363 => conv_std_logic_vector(37665, 16),
62364 => conv_std_logic_vector(37908, 16),
62365 => conv_std_logic_vector(38151, 16),
62366 => conv_std_logic_vector(38394, 16),
62367 => conv_std_logic_vector(38637, 16),
62368 => conv_std_logic_vector(38880, 16),
62369 => conv_std_logic_vector(39123, 16),
62370 => conv_std_logic_vector(39366, 16),
62371 => conv_std_logic_vector(39609, 16),
62372 => conv_std_logic_vector(39852, 16),
62373 => conv_std_logic_vector(40095, 16),
62374 => conv_std_logic_vector(40338, 16),
62375 => conv_std_logic_vector(40581, 16),
62376 => conv_std_logic_vector(40824, 16),
62377 => conv_std_logic_vector(41067, 16),
62378 => conv_std_logic_vector(41310, 16),
62379 => conv_std_logic_vector(41553, 16),
62380 => conv_std_logic_vector(41796, 16),
62381 => conv_std_logic_vector(42039, 16),
62382 => conv_std_logic_vector(42282, 16),
62383 => conv_std_logic_vector(42525, 16),
62384 => conv_std_logic_vector(42768, 16),
62385 => conv_std_logic_vector(43011, 16),
62386 => conv_std_logic_vector(43254, 16),
62387 => conv_std_logic_vector(43497, 16),
62388 => conv_std_logic_vector(43740, 16),
62389 => conv_std_logic_vector(43983, 16),
62390 => conv_std_logic_vector(44226, 16),
62391 => conv_std_logic_vector(44469, 16),
62392 => conv_std_logic_vector(44712, 16),
62393 => conv_std_logic_vector(44955, 16),
62394 => conv_std_logic_vector(45198, 16),
62395 => conv_std_logic_vector(45441, 16),
62396 => conv_std_logic_vector(45684, 16),
62397 => conv_std_logic_vector(45927, 16),
62398 => conv_std_logic_vector(46170, 16),
62399 => conv_std_logic_vector(46413, 16),
62400 => conv_std_logic_vector(46656, 16),
62401 => conv_std_logic_vector(46899, 16),
62402 => conv_std_logic_vector(47142, 16),
62403 => conv_std_logic_vector(47385, 16),
62404 => conv_std_logic_vector(47628, 16),
62405 => conv_std_logic_vector(47871, 16),
62406 => conv_std_logic_vector(48114, 16),
62407 => conv_std_logic_vector(48357, 16),
62408 => conv_std_logic_vector(48600, 16),
62409 => conv_std_logic_vector(48843, 16),
62410 => conv_std_logic_vector(49086, 16),
62411 => conv_std_logic_vector(49329, 16),
62412 => conv_std_logic_vector(49572, 16),
62413 => conv_std_logic_vector(49815, 16),
62414 => conv_std_logic_vector(50058, 16),
62415 => conv_std_logic_vector(50301, 16),
62416 => conv_std_logic_vector(50544, 16),
62417 => conv_std_logic_vector(50787, 16),
62418 => conv_std_logic_vector(51030, 16),
62419 => conv_std_logic_vector(51273, 16),
62420 => conv_std_logic_vector(51516, 16),
62421 => conv_std_logic_vector(51759, 16),
62422 => conv_std_logic_vector(52002, 16),
62423 => conv_std_logic_vector(52245, 16),
62424 => conv_std_logic_vector(52488, 16),
62425 => conv_std_logic_vector(52731, 16),
62426 => conv_std_logic_vector(52974, 16),
62427 => conv_std_logic_vector(53217, 16),
62428 => conv_std_logic_vector(53460, 16),
62429 => conv_std_logic_vector(53703, 16),
62430 => conv_std_logic_vector(53946, 16),
62431 => conv_std_logic_vector(54189, 16),
62432 => conv_std_logic_vector(54432, 16),
62433 => conv_std_logic_vector(54675, 16),
62434 => conv_std_logic_vector(54918, 16),
62435 => conv_std_logic_vector(55161, 16),
62436 => conv_std_logic_vector(55404, 16),
62437 => conv_std_logic_vector(55647, 16),
62438 => conv_std_logic_vector(55890, 16),
62439 => conv_std_logic_vector(56133, 16),
62440 => conv_std_logic_vector(56376, 16),
62441 => conv_std_logic_vector(56619, 16),
62442 => conv_std_logic_vector(56862, 16),
62443 => conv_std_logic_vector(57105, 16),
62444 => conv_std_logic_vector(57348, 16),
62445 => conv_std_logic_vector(57591, 16),
62446 => conv_std_logic_vector(57834, 16),
62447 => conv_std_logic_vector(58077, 16),
62448 => conv_std_logic_vector(58320, 16),
62449 => conv_std_logic_vector(58563, 16),
62450 => conv_std_logic_vector(58806, 16),
62451 => conv_std_logic_vector(59049, 16),
62452 => conv_std_logic_vector(59292, 16),
62453 => conv_std_logic_vector(59535, 16),
62454 => conv_std_logic_vector(59778, 16),
62455 => conv_std_logic_vector(60021, 16),
62456 => conv_std_logic_vector(60264, 16),
62457 => conv_std_logic_vector(60507, 16),
62458 => conv_std_logic_vector(60750, 16),
62459 => conv_std_logic_vector(60993, 16),
62460 => conv_std_logic_vector(61236, 16),
62461 => conv_std_logic_vector(61479, 16),
62462 => conv_std_logic_vector(61722, 16),
62463 => conv_std_logic_vector(61965, 16),
62464 => conv_std_logic_vector(0, 16),
62465 => conv_std_logic_vector(244, 16),
62466 => conv_std_logic_vector(488, 16),
62467 => conv_std_logic_vector(732, 16),
62468 => conv_std_logic_vector(976, 16),
62469 => conv_std_logic_vector(1220, 16),
62470 => conv_std_logic_vector(1464, 16),
62471 => conv_std_logic_vector(1708, 16),
62472 => conv_std_logic_vector(1952, 16),
62473 => conv_std_logic_vector(2196, 16),
62474 => conv_std_logic_vector(2440, 16),
62475 => conv_std_logic_vector(2684, 16),
62476 => conv_std_logic_vector(2928, 16),
62477 => conv_std_logic_vector(3172, 16),
62478 => conv_std_logic_vector(3416, 16),
62479 => conv_std_logic_vector(3660, 16),
62480 => conv_std_logic_vector(3904, 16),
62481 => conv_std_logic_vector(4148, 16),
62482 => conv_std_logic_vector(4392, 16),
62483 => conv_std_logic_vector(4636, 16),
62484 => conv_std_logic_vector(4880, 16),
62485 => conv_std_logic_vector(5124, 16),
62486 => conv_std_logic_vector(5368, 16),
62487 => conv_std_logic_vector(5612, 16),
62488 => conv_std_logic_vector(5856, 16),
62489 => conv_std_logic_vector(6100, 16),
62490 => conv_std_logic_vector(6344, 16),
62491 => conv_std_logic_vector(6588, 16),
62492 => conv_std_logic_vector(6832, 16),
62493 => conv_std_logic_vector(7076, 16),
62494 => conv_std_logic_vector(7320, 16),
62495 => conv_std_logic_vector(7564, 16),
62496 => conv_std_logic_vector(7808, 16),
62497 => conv_std_logic_vector(8052, 16),
62498 => conv_std_logic_vector(8296, 16),
62499 => conv_std_logic_vector(8540, 16),
62500 => conv_std_logic_vector(8784, 16),
62501 => conv_std_logic_vector(9028, 16),
62502 => conv_std_logic_vector(9272, 16),
62503 => conv_std_logic_vector(9516, 16),
62504 => conv_std_logic_vector(9760, 16),
62505 => conv_std_logic_vector(10004, 16),
62506 => conv_std_logic_vector(10248, 16),
62507 => conv_std_logic_vector(10492, 16),
62508 => conv_std_logic_vector(10736, 16),
62509 => conv_std_logic_vector(10980, 16),
62510 => conv_std_logic_vector(11224, 16),
62511 => conv_std_logic_vector(11468, 16),
62512 => conv_std_logic_vector(11712, 16),
62513 => conv_std_logic_vector(11956, 16),
62514 => conv_std_logic_vector(12200, 16),
62515 => conv_std_logic_vector(12444, 16),
62516 => conv_std_logic_vector(12688, 16),
62517 => conv_std_logic_vector(12932, 16),
62518 => conv_std_logic_vector(13176, 16),
62519 => conv_std_logic_vector(13420, 16),
62520 => conv_std_logic_vector(13664, 16),
62521 => conv_std_logic_vector(13908, 16),
62522 => conv_std_logic_vector(14152, 16),
62523 => conv_std_logic_vector(14396, 16),
62524 => conv_std_logic_vector(14640, 16),
62525 => conv_std_logic_vector(14884, 16),
62526 => conv_std_logic_vector(15128, 16),
62527 => conv_std_logic_vector(15372, 16),
62528 => conv_std_logic_vector(15616, 16),
62529 => conv_std_logic_vector(15860, 16),
62530 => conv_std_logic_vector(16104, 16),
62531 => conv_std_logic_vector(16348, 16),
62532 => conv_std_logic_vector(16592, 16),
62533 => conv_std_logic_vector(16836, 16),
62534 => conv_std_logic_vector(17080, 16),
62535 => conv_std_logic_vector(17324, 16),
62536 => conv_std_logic_vector(17568, 16),
62537 => conv_std_logic_vector(17812, 16),
62538 => conv_std_logic_vector(18056, 16),
62539 => conv_std_logic_vector(18300, 16),
62540 => conv_std_logic_vector(18544, 16),
62541 => conv_std_logic_vector(18788, 16),
62542 => conv_std_logic_vector(19032, 16),
62543 => conv_std_logic_vector(19276, 16),
62544 => conv_std_logic_vector(19520, 16),
62545 => conv_std_logic_vector(19764, 16),
62546 => conv_std_logic_vector(20008, 16),
62547 => conv_std_logic_vector(20252, 16),
62548 => conv_std_logic_vector(20496, 16),
62549 => conv_std_logic_vector(20740, 16),
62550 => conv_std_logic_vector(20984, 16),
62551 => conv_std_logic_vector(21228, 16),
62552 => conv_std_logic_vector(21472, 16),
62553 => conv_std_logic_vector(21716, 16),
62554 => conv_std_logic_vector(21960, 16),
62555 => conv_std_logic_vector(22204, 16),
62556 => conv_std_logic_vector(22448, 16),
62557 => conv_std_logic_vector(22692, 16),
62558 => conv_std_logic_vector(22936, 16),
62559 => conv_std_logic_vector(23180, 16),
62560 => conv_std_logic_vector(23424, 16),
62561 => conv_std_logic_vector(23668, 16),
62562 => conv_std_logic_vector(23912, 16),
62563 => conv_std_logic_vector(24156, 16),
62564 => conv_std_logic_vector(24400, 16),
62565 => conv_std_logic_vector(24644, 16),
62566 => conv_std_logic_vector(24888, 16),
62567 => conv_std_logic_vector(25132, 16),
62568 => conv_std_logic_vector(25376, 16),
62569 => conv_std_logic_vector(25620, 16),
62570 => conv_std_logic_vector(25864, 16),
62571 => conv_std_logic_vector(26108, 16),
62572 => conv_std_logic_vector(26352, 16),
62573 => conv_std_logic_vector(26596, 16),
62574 => conv_std_logic_vector(26840, 16),
62575 => conv_std_logic_vector(27084, 16),
62576 => conv_std_logic_vector(27328, 16),
62577 => conv_std_logic_vector(27572, 16),
62578 => conv_std_logic_vector(27816, 16),
62579 => conv_std_logic_vector(28060, 16),
62580 => conv_std_logic_vector(28304, 16),
62581 => conv_std_logic_vector(28548, 16),
62582 => conv_std_logic_vector(28792, 16),
62583 => conv_std_logic_vector(29036, 16),
62584 => conv_std_logic_vector(29280, 16),
62585 => conv_std_logic_vector(29524, 16),
62586 => conv_std_logic_vector(29768, 16),
62587 => conv_std_logic_vector(30012, 16),
62588 => conv_std_logic_vector(30256, 16),
62589 => conv_std_logic_vector(30500, 16),
62590 => conv_std_logic_vector(30744, 16),
62591 => conv_std_logic_vector(30988, 16),
62592 => conv_std_logic_vector(31232, 16),
62593 => conv_std_logic_vector(31476, 16),
62594 => conv_std_logic_vector(31720, 16),
62595 => conv_std_logic_vector(31964, 16),
62596 => conv_std_logic_vector(32208, 16),
62597 => conv_std_logic_vector(32452, 16),
62598 => conv_std_logic_vector(32696, 16),
62599 => conv_std_logic_vector(32940, 16),
62600 => conv_std_logic_vector(33184, 16),
62601 => conv_std_logic_vector(33428, 16),
62602 => conv_std_logic_vector(33672, 16),
62603 => conv_std_logic_vector(33916, 16),
62604 => conv_std_logic_vector(34160, 16),
62605 => conv_std_logic_vector(34404, 16),
62606 => conv_std_logic_vector(34648, 16),
62607 => conv_std_logic_vector(34892, 16),
62608 => conv_std_logic_vector(35136, 16),
62609 => conv_std_logic_vector(35380, 16),
62610 => conv_std_logic_vector(35624, 16),
62611 => conv_std_logic_vector(35868, 16),
62612 => conv_std_logic_vector(36112, 16),
62613 => conv_std_logic_vector(36356, 16),
62614 => conv_std_logic_vector(36600, 16),
62615 => conv_std_logic_vector(36844, 16),
62616 => conv_std_logic_vector(37088, 16),
62617 => conv_std_logic_vector(37332, 16),
62618 => conv_std_logic_vector(37576, 16),
62619 => conv_std_logic_vector(37820, 16),
62620 => conv_std_logic_vector(38064, 16),
62621 => conv_std_logic_vector(38308, 16),
62622 => conv_std_logic_vector(38552, 16),
62623 => conv_std_logic_vector(38796, 16),
62624 => conv_std_logic_vector(39040, 16),
62625 => conv_std_logic_vector(39284, 16),
62626 => conv_std_logic_vector(39528, 16),
62627 => conv_std_logic_vector(39772, 16),
62628 => conv_std_logic_vector(40016, 16),
62629 => conv_std_logic_vector(40260, 16),
62630 => conv_std_logic_vector(40504, 16),
62631 => conv_std_logic_vector(40748, 16),
62632 => conv_std_logic_vector(40992, 16),
62633 => conv_std_logic_vector(41236, 16),
62634 => conv_std_logic_vector(41480, 16),
62635 => conv_std_logic_vector(41724, 16),
62636 => conv_std_logic_vector(41968, 16),
62637 => conv_std_logic_vector(42212, 16),
62638 => conv_std_logic_vector(42456, 16),
62639 => conv_std_logic_vector(42700, 16),
62640 => conv_std_logic_vector(42944, 16),
62641 => conv_std_logic_vector(43188, 16),
62642 => conv_std_logic_vector(43432, 16),
62643 => conv_std_logic_vector(43676, 16),
62644 => conv_std_logic_vector(43920, 16),
62645 => conv_std_logic_vector(44164, 16),
62646 => conv_std_logic_vector(44408, 16),
62647 => conv_std_logic_vector(44652, 16),
62648 => conv_std_logic_vector(44896, 16),
62649 => conv_std_logic_vector(45140, 16),
62650 => conv_std_logic_vector(45384, 16),
62651 => conv_std_logic_vector(45628, 16),
62652 => conv_std_logic_vector(45872, 16),
62653 => conv_std_logic_vector(46116, 16),
62654 => conv_std_logic_vector(46360, 16),
62655 => conv_std_logic_vector(46604, 16),
62656 => conv_std_logic_vector(46848, 16),
62657 => conv_std_logic_vector(47092, 16),
62658 => conv_std_logic_vector(47336, 16),
62659 => conv_std_logic_vector(47580, 16),
62660 => conv_std_logic_vector(47824, 16),
62661 => conv_std_logic_vector(48068, 16),
62662 => conv_std_logic_vector(48312, 16),
62663 => conv_std_logic_vector(48556, 16),
62664 => conv_std_logic_vector(48800, 16),
62665 => conv_std_logic_vector(49044, 16),
62666 => conv_std_logic_vector(49288, 16),
62667 => conv_std_logic_vector(49532, 16),
62668 => conv_std_logic_vector(49776, 16),
62669 => conv_std_logic_vector(50020, 16),
62670 => conv_std_logic_vector(50264, 16),
62671 => conv_std_logic_vector(50508, 16),
62672 => conv_std_logic_vector(50752, 16),
62673 => conv_std_logic_vector(50996, 16),
62674 => conv_std_logic_vector(51240, 16),
62675 => conv_std_logic_vector(51484, 16),
62676 => conv_std_logic_vector(51728, 16),
62677 => conv_std_logic_vector(51972, 16),
62678 => conv_std_logic_vector(52216, 16),
62679 => conv_std_logic_vector(52460, 16),
62680 => conv_std_logic_vector(52704, 16),
62681 => conv_std_logic_vector(52948, 16),
62682 => conv_std_logic_vector(53192, 16),
62683 => conv_std_logic_vector(53436, 16),
62684 => conv_std_logic_vector(53680, 16),
62685 => conv_std_logic_vector(53924, 16),
62686 => conv_std_logic_vector(54168, 16),
62687 => conv_std_logic_vector(54412, 16),
62688 => conv_std_logic_vector(54656, 16),
62689 => conv_std_logic_vector(54900, 16),
62690 => conv_std_logic_vector(55144, 16),
62691 => conv_std_logic_vector(55388, 16),
62692 => conv_std_logic_vector(55632, 16),
62693 => conv_std_logic_vector(55876, 16),
62694 => conv_std_logic_vector(56120, 16),
62695 => conv_std_logic_vector(56364, 16),
62696 => conv_std_logic_vector(56608, 16),
62697 => conv_std_logic_vector(56852, 16),
62698 => conv_std_logic_vector(57096, 16),
62699 => conv_std_logic_vector(57340, 16),
62700 => conv_std_logic_vector(57584, 16),
62701 => conv_std_logic_vector(57828, 16),
62702 => conv_std_logic_vector(58072, 16),
62703 => conv_std_logic_vector(58316, 16),
62704 => conv_std_logic_vector(58560, 16),
62705 => conv_std_logic_vector(58804, 16),
62706 => conv_std_logic_vector(59048, 16),
62707 => conv_std_logic_vector(59292, 16),
62708 => conv_std_logic_vector(59536, 16),
62709 => conv_std_logic_vector(59780, 16),
62710 => conv_std_logic_vector(60024, 16),
62711 => conv_std_logic_vector(60268, 16),
62712 => conv_std_logic_vector(60512, 16),
62713 => conv_std_logic_vector(60756, 16),
62714 => conv_std_logic_vector(61000, 16),
62715 => conv_std_logic_vector(61244, 16),
62716 => conv_std_logic_vector(61488, 16),
62717 => conv_std_logic_vector(61732, 16),
62718 => conv_std_logic_vector(61976, 16),
62719 => conv_std_logic_vector(62220, 16),
62720 => conv_std_logic_vector(0, 16),
62721 => conv_std_logic_vector(245, 16),
62722 => conv_std_logic_vector(490, 16),
62723 => conv_std_logic_vector(735, 16),
62724 => conv_std_logic_vector(980, 16),
62725 => conv_std_logic_vector(1225, 16),
62726 => conv_std_logic_vector(1470, 16),
62727 => conv_std_logic_vector(1715, 16),
62728 => conv_std_logic_vector(1960, 16),
62729 => conv_std_logic_vector(2205, 16),
62730 => conv_std_logic_vector(2450, 16),
62731 => conv_std_logic_vector(2695, 16),
62732 => conv_std_logic_vector(2940, 16),
62733 => conv_std_logic_vector(3185, 16),
62734 => conv_std_logic_vector(3430, 16),
62735 => conv_std_logic_vector(3675, 16),
62736 => conv_std_logic_vector(3920, 16),
62737 => conv_std_logic_vector(4165, 16),
62738 => conv_std_logic_vector(4410, 16),
62739 => conv_std_logic_vector(4655, 16),
62740 => conv_std_logic_vector(4900, 16),
62741 => conv_std_logic_vector(5145, 16),
62742 => conv_std_logic_vector(5390, 16),
62743 => conv_std_logic_vector(5635, 16),
62744 => conv_std_logic_vector(5880, 16),
62745 => conv_std_logic_vector(6125, 16),
62746 => conv_std_logic_vector(6370, 16),
62747 => conv_std_logic_vector(6615, 16),
62748 => conv_std_logic_vector(6860, 16),
62749 => conv_std_logic_vector(7105, 16),
62750 => conv_std_logic_vector(7350, 16),
62751 => conv_std_logic_vector(7595, 16),
62752 => conv_std_logic_vector(7840, 16),
62753 => conv_std_logic_vector(8085, 16),
62754 => conv_std_logic_vector(8330, 16),
62755 => conv_std_logic_vector(8575, 16),
62756 => conv_std_logic_vector(8820, 16),
62757 => conv_std_logic_vector(9065, 16),
62758 => conv_std_logic_vector(9310, 16),
62759 => conv_std_logic_vector(9555, 16),
62760 => conv_std_logic_vector(9800, 16),
62761 => conv_std_logic_vector(10045, 16),
62762 => conv_std_logic_vector(10290, 16),
62763 => conv_std_logic_vector(10535, 16),
62764 => conv_std_logic_vector(10780, 16),
62765 => conv_std_logic_vector(11025, 16),
62766 => conv_std_logic_vector(11270, 16),
62767 => conv_std_logic_vector(11515, 16),
62768 => conv_std_logic_vector(11760, 16),
62769 => conv_std_logic_vector(12005, 16),
62770 => conv_std_logic_vector(12250, 16),
62771 => conv_std_logic_vector(12495, 16),
62772 => conv_std_logic_vector(12740, 16),
62773 => conv_std_logic_vector(12985, 16),
62774 => conv_std_logic_vector(13230, 16),
62775 => conv_std_logic_vector(13475, 16),
62776 => conv_std_logic_vector(13720, 16),
62777 => conv_std_logic_vector(13965, 16),
62778 => conv_std_logic_vector(14210, 16),
62779 => conv_std_logic_vector(14455, 16),
62780 => conv_std_logic_vector(14700, 16),
62781 => conv_std_logic_vector(14945, 16),
62782 => conv_std_logic_vector(15190, 16),
62783 => conv_std_logic_vector(15435, 16),
62784 => conv_std_logic_vector(15680, 16),
62785 => conv_std_logic_vector(15925, 16),
62786 => conv_std_logic_vector(16170, 16),
62787 => conv_std_logic_vector(16415, 16),
62788 => conv_std_logic_vector(16660, 16),
62789 => conv_std_logic_vector(16905, 16),
62790 => conv_std_logic_vector(17150, 16),
62791 => conv_std_logic_vector(17395, 16),
62792 => conv_std_logic_vector(17640, 16),
62793 => conv_std_logic_vector(17885, 16),
62794 => conv_std_logic_vector(18130, 16),
62795 => conv_std_logic_vector(18375, 16),
62796 => conv_std_logic_vector(18620, 16),
62797 => conv_std_logic_vector(18865, 16),
62798 => conv_std_logic_vector(19110, 16),
62799 => conv_std_logic_vector(19355, 16),
62800 => conv_std_logic_vector(19600, 16),
62801 => conv_std_logic_vector(19845, 16),
62802 => conv_std_logic_vector(20090, 16),
62803 => conv_std_logic_vector(20335, 16),
62804 => conv_std_logic_vector(20580, 16),
62805 => conv_std_logic_vector(20825, 16),
62806 => conv_std_logic_vector(21070, 16),
62807 => conv_std_logic_vector(21315, 16),
62808 => conv_std_logic_vector(21560, 16),
62809 => conv_std_logic_vector(21805, 16),
62810 => conv_std_logic_vector(22050, 16),
62811 => conv_std_logic_vector(22295, 16),
62812 => conv_std_logic_vector(22540, 16),
62813 => conv_std_logic_vector(22785, 16),
62814 => conv_std_logic_vector(23030, 16),
62815 => conv_std_logic_vector(23275, 16),
62816 => conv_std_logic_vector(23520, 16),
62817 => conv_std_logic_vector(23765, 16),
62818 => conv_std_logic_vector(24010, 16),
62819 => conv_std_logic_vector(24255, 16),
62820 => conv_std_logic_vector(24500, 16),
62821 => conv_std_logic_vector(24745, 16),
62822 => conv_std_logic_vector(24990, 16),
62823 => conv_std_logic_vector(25235, 16),
62824 => conv_std_logic_vector(25480, 16),
62825 => conv_std_logic_vector(25725, 16),
62826 => conv_std_logic_vector(25970, 16),
62827 => conv_std_logic_vector(26215, 16),
62828 => conv_std_logic_vector(26460, 16),
62829 => conv_std_logic_vector(26705, 16),
62830 => conv_std_logic_vector(26950, 16),
62831 => conv_std_logic_vector(27195, 16),
62832 => conv_std_logic_vector(27440, 16),
62833 => conv_std_logic_vector(27685, 16),
62834 => conv_std_logic_vector(27930, 16),
62835 => conv_std_logic_vector(28175, 16),
62836 => conv_std_logic_vector(28420, 16),
62837 => conv_std_logic_vector(28665, 16),
62838 => conv_std_logic_vector(28910, 16),
62839 => conv_std_logic_vector(29155, 16),
62840 => conv_std_logic_vector(29400, 16),
62841 => conv_std_logic_vector(29645, 16),
62842 => conv_std_logic_vector(29890, 16),
62843 => conv_std_logic_vector(30135, 16),
62844 => conv_std_logic_vector(30380, 16),
62845 => conv_std_logic_vector(30625, 16),
62846 => conv_std_logic_vector(30870, 16),
62847 => conv_std_logic_vector(31115, 16),
62848 => conv_std_logic_vector(31360, 16),
62849 => conv_std_logic_vector(31605, 16),
62850 => conv_std_logic_vector(31850, 16),
62851 => conv_std_logic_vector(32095, 16),
62852 => conv_std_logic_vector(32340, 16),
62853 => conv_std_logic_vector(32585, 16),
62854 => conv_std_logic_vector(32830, 16),
62855 => conv_std_logic_vector(33075, 16),
62856 => conv_std_logic_vector(33320, 16),
62857 => conv_std_logic_vector(33565, 16),
62858 => conv_std_logic_vector(33810, 16),
62859 => conv_std_logic_vector(34055, 16),
62860 => conv_std_logic_vector(34300, 16),
62861 => conv_std_logic_vector(34545, 16),
62862 => conv_std_logic_vector(34790, 16),
62863 => conv_std_logic_vector(35035, 16),
62864 => conv_std_logic_vector(35280, 16),
62865 => conv_std_logic_vector(35525, 16),
62866 => conv_std_logic_vector(35770, 16),
62867 => conv_std_logic_vector(36015, 16),
62868 => conv_std_logic_vector(36260, 16),
62869 => conv_std_logic_vector(36505, 16),
62870 => conv_std_logic_vector(36750, 16),
62871 => conv_std_logic_vector(36995, 16),
62872 => conv_std_logic_vector(37240, 16),
62873 => conv_std_logic_vector(37485, 16),
62874 => conv_std_logic_vector(37730, 16),
62875 => conv_std_logic_vector(37975, 16),
62876 => conv_std_logic_vector(38220, 16),
62877 => conv_std_logic_vector(38465, 16),
62878 => conv_std_logic_vector(38710, 16),
62879 => conv_std_logic_vector(38955, 16),
62880 => conv_std_logic_vector(39200, 16),
62881 => conv_std_logic_vector(39445, 16),
62882 => conv_std_logic_vector(39690, 16),
62883 => conv_std_logic_vector(39935, 16),
62884 => conv_std_logic_vector(40180, 16),
62885 => conv_std_logic_vector(40425, 16),
62886 => conv_std_logic_vector(40670, 16),
62887 => conv_std_logic_vector(40915, 16),
62888 => conv_std_logic_vector(41160, 16),
62889 => conv_std_logic_vector(41405, 16),
62890 => conv_std_logic_vector(41650, 16),
62891 => conv_std_logic_vector(41895, 16),
62892 => conv_std_logic_vector(42140, 16),
62893 => conv_std_logic_vector(42385, 16),
62894 => conv_std_logic_vector(42630, 16),
62895 => conv_std_logic_vector(42875, 16),
62896 => conv_std_logic_vector(43120, 16),
62897 => conv_std_logic_vector(43365, 16),
62898 => conv_std_logic_vector(43610, 16),
62899 => conv_std_logic_vector(43855, 16),
62900 => conv_std_logic_vector(44100, 16),
62901 => conv_std_logic_vector(44345, 16),
62902 => conv_std_logic_vector(44590, 16),
62903 => conv_std_logic_vector(44835, 16),
62904 => conv_std_logic_vector(45080, 16),
62905 => conv_std_logic_vector(45325, 16),
62906 => conv_std_logic_vector(45570, 16),
62907 => conv_std_logic_vector(45815, 16),
62908 => conv_std_logic_vector(46060, 16),
62909 => conv_std_logic_vector(46305, 16),
62910 => conv_std_logic_vector(46550, 16),
62911 => conv_std_logic_vector(46795, 16),
62912 => conv_std_logic_vector(47040, 16),
62913 => conv_std_logic_vector(47285, 16),
62914 => conv_std_logic_vector(47530, 16),
62915 => conv_std_logic_vector(47775, 16),
62916 => conv_std_logic_vector(48020, 16),
62917 => conv_std_logic_vector(48265, 16),
62918 => conv_std_logic_vector(48510, 16),
62919 => conv_std_logic_vector(48755, 16),
62920 => conv_std_logic_vector(49000, 16),
62921 => conv_std_logic_vector(49245, 16),
62922 => conv_std_logic_vector(49490, 16),
62923 => conv_std_logic_vector(49735, 16),
62924 => conv_std_logic_vector(49980, 16),
62925 => conv_std_logic_vector(50225, 16),
62926 => conv_std_logic_vector(50470, 16),
62927 => conv_std_logic_vector(50715, 16),
62928 => conv_std_logic_vector(50960, 16),
62929 => conv_std_logic_vector(51205, 16),
62930 => conv_std_logic_vector(51450, 16),
62931 => conv_std_logic_vector(51695, 16),
62932 => conv_std_logic_vector(51940, 16),
62933 => conv_std_logic_vector(52185, 16),
62934 => conv_std_logic_vector(52430, 16),
62935 => conv_std_logic_vector(52675, 16),
62936 => conv_std_logic_vector(52920, 16),
62937 => conv_std_logic_vector(53165, 16),
62938 => conv_std_logic_vector(53410, 16),
62939 => conv_std_logic_vector(53655, 16),
62940 => conv_std_logic_vector(53900, 16),
62941 => conv_std_logic_vector(54145, 16),
62942 => conv_std_logic_vector(54390, 16),
62943 => conv_std_logic_vector(54635, 16),
62944 => conv_std_logic_vector(54880, 16),
62945 => conv_std_logic_vector(55125, 16),
62946 => conv_std_logic_vector(55370, 16),
62947 => conv_std_logic_vector(55615, 16),
62948 => conv_std_logic_vector(55860, 16),
62949 => conv_std_logic_vector(56105, 16),
62950 => conv_std_logic_vector(56350, 16),
62951 => conv_std_logic_vector(56595, 16),
62952 => conv_std_logic_vector(56840, 16),
62953 => conv_std_logic_vector(57085, 16),
62954 => conv_std_logic_vector(57330, 16),
62955 => conv_std_logic_vector(57575, 16),
62956 => conv_std_logic_vector(57820, 16),
62957 => conv_std_logic_vector(58065, 16),
62958 => conv_std_logic_vector(58310, 16),
62959 => conv_std_logic_vector(58555, 16),
62960 => conv_std_logic_vector(58800, 16),
62961 => conv_std_logic_vector(59045, 16),
62962 => conv_std_logic_vector(59290, 16),
62963 => conv_std_logic_vector(59535, 16),
62964 => conv_std_logic_vector(59780, 16),
62965 => conv_std_logic_vector(60025, 16),
62966 => conv_std_logic_vector(60270, 16),
62967 => conv_std_logic_vector(60515, 16),
62968 => conv_std_logic_vector(60760, 16),
62969 => conv_std_logic_vector(61005, 16),
62970 => conv_std_logic_vector(61250, 16),
62971 => conv_std_logic_vector(61495, 16),
62972 => conv_std_logic_vector(61740, 16),
62973 => conv_std_logic_vector(61985, 16),
62974 => conv_std_logic_vector(62230, 16),
62975 => conv_std_logic_vector(62475, 16),
62976 => conv_std_logic_vector(0, 16),
62977 => conv_std_logic_vector(246, 16),
62978 => conv_std_logic_vector(492, 16),
62979 => conv_std_logic_vector(738, 16),
62980 => conv_std_logic_vector(984, 16),
62981 => conv_std_logic_vector(1230, 16),
62982 => conv_std_logic_vector(1476, 16),
62983 => conv_std_logic_vector(1722, 16),
62984 => conv_std_logic_vector(1968, 16),
62985 => conv_std_logic_vector(2214, 16),
62986 => conv_std_logic_vector(2460, 16),
62987 => conv_std_logic_vector(2706, 16),
62988 => conv_std_logic_vector(2952, 16),
62989 => conv_std_logic_vector(3198, 16),
62990 => conv_std_logic_vector(3444, 16),
62991 => conv_std_logic_vector(3690, 16),
62992 => conv_std_logic_vector(3936, 16),
62993 => conv_std_logic_vector(4182, 16),
62994 => conv_std_logic_vector(4428, 16),
62995 => conv_std_logic_vector(4674, 16),
62996 => conv_std_logic_vector(4920, 16),
62997 => conv_std_logic_vector(5166, 16),
62998 => conv_std_logic_vector(5412, 16),
62999 => conv_std_logic_vector(5658, 16),
63000 => conv_std_logic_vector(5904, 16),
63001 => conv_std_logic_vector(6150, 16),
63002 => conv_std_logic_vector(6396, 16),
63003 => conv_std_logic_vector(6642, 16),
63004 => conv_std_logic_vector(6888, 16),
63005 => conv_std_logic_vector(7134, 16),
63006 => conv_std_logic_vector(7380, 16),
63007 => conv_std_logic_vector(7626, 16),
63008 => conv_std_logic_vector(7872, 16),
63009 => conv_std_logic_vector(8118, 16),
63010 => conv_std_logic_vector(8364, 16),
63011 => conv_std_logic_vector(8610, 16),
63012 => conv_std_logic_vector(8856, 16),
63013 => conv_std_logic_vector(9102, 16),
63014 => conv_std_logic_vector(9348, 16),
63015 => conv_std_logic_vector(9594, 16),
63016 => conv_std_logic_vector(9840, 16),
63017 => conv_std_logic_vector(10086, 16),
63018 => conv_std_logic_vector(10332, 16),
63019 => conv_std_logic_vector(10578, 16),
63020 => conv_std_logic_vector(10824, 16),
63021 => conv_std_logic_vector(11070, 16),
63022 => conv_std_logic_vector(11316, 16),
63023 => conv_std_logic_vector(11562, 16),
63024 => conv_std_logic_vector(11808, 16),
63025 => conv_std_logic_vector(12054, 16),
63026 => conv_std_logic_vector(12300, 16),
63027 => conv_std_logic_vector(12546, 16),
63028 => conv_std_logic_vector(12792, 16),
63029 => conv_std_logic_vector(13038, 16),
63030 => conv_std_logic_vector(13284, 16),
63031 => conv_std_logic_vector(13530, 16),
63032 => conv_std_logic_vector(13776, 16),
63033 => conv_std_logic_vector(14022, 16),
63034 => conv_std_logic_vector(14268, 16),
63035 => conv_std_logic_vector(14514, 16),
63036 => conv_std_logic_vector(14760, 16),
63037 => conv_std_logic_vector(15006, 16),
63038 => conv_std_logic_vector(15252, 16),
63039 => conv_std_logic_vector(15498, 16),
63040 => conv_std_logic_vector(15744, 16),
63041 => conv_std_logic_vector(15990, 16),
63042 => conv_std_logic_vector(16236, 16),
63043 => conv_std_logic_vector(16482, 16),
63044 => conv_std_logic_vector(16728, 16),
63045 => conv_std_logic_vector(16974, 16),
63046 => conv_std_logic_vector(17220, 16),
63047 => conv_std_logic_vector(17466, 16),
63048 => conv_std_logic_vector(17712, 16),
63049 => conv_std_logic_vector(17958, 16),
63050 => conv_std_logic_vector(18204, 16),
63051 => conv_std_logic_vector(18450, 16),
63052 => conv_std_logic_vector(18696, 16),
63053 => conv_std_logic_vector(18942, 16),
63054 => conv_std_logic_vector(19188, 16),
63055 => conv_std_logic_vector(19434, 16),
63056 => conv_std_logic_vector(19680, 16),
63057 => conv_std_logic_vector(19926, 16),
63058 => conv_std_logic_vector(20172, 16),
63059 => conv_std_logic_vector(20418, 16),
63060 => conv_std_logic_vector(20664, 16),
63061 => conv_std_logic_vector(20910, 16),
63062 => conv_std_logic_vector(21156, 16),
63063 => conv_std_logic_vector(21402, 16),
63064 => conv_std_logic_vector(21648, 16),
63065 => conv_std_logic_vector(21894, 16),
63066 => conv_std_logic_vector(22140, 16),
63067 => conv_std_logic_vector(22386, 16),
63068 => conv_std_logic_vector(22632, 16),
63069 => conv_std_logic_vector(22878, 16),
63070 => conv_std_logic_vector(23124, 16),
63071 => conv_std_logic_vector(23370, 16),
63072 => conv_std_logic_vector(23616, 16),
63073 => conv_std_logic_vector(23862, 16),
63074 => conv_std_logic_vector(24108, 16),
63075 => conv_std_logic_vector(24354, 16),
63076 => conv_std_logic_vector(24600, 16),
63077 => conv_std_logic_vector(24846, 16),
63078 => conv_std_logic_vector(25092, 16),
63079 => conv_std_logic_vector(25338, 16),
63080 => conv_std_logic_vector(25584, 16),
63081 => conv_std_logic_vector(25830, 16),
63082 => conv_std_logic_vector(26076, 16),
63083 => conv_std_logic_vector(26322, 16),
63084 => conv_std_logic_vector(26568, 16),
63085 => conv_std_logic_vector(26814, 16),
63086 => conv_std_logic_vector(27060, 16),
63087 => conv_std_logic_vector(27306, 16),
63088 => conv_std_logic_vector(27552, 16),
63089 => conv_std_logic_vector(27798, 16),
63090 => conv_std_logic_vector(28044, 16),
63091 => conv_std_logic_vector(28290, 16),
63092 => conv_std_logic_vector(28536, 16),
63093 => conv_std_logic_vector(28782, 16),
63094 => conv_std_logic_vector(29028, 16),
63095 => conv_std_logic_vector(29274, 16),
63096 => conv_std_logic_vector(29520, 16),
63097 => conv_std_logic_vector(29766, 16),
63098 => conv_std_logic_vector(30012, 16),
63099 => conv_std_logic_vector(30258, 16),
63100 => conv_std_logic_vector(30504, 16),
63101 => conv_std_logic_vector(30750, 16),
63102 => conv_std_logic_vector(30996, 16),
63103 => conv_std_logic_vector(31242, 16),
63104 => conv_std_logic_vector(31488, 16),
63105 => conv_std_logic_vector(31734, 16),
63106 => conv_std_logic_vector(31980, 16),
63107 => conv_std_logic_vector(32226, 16),
63108 => conv_std_logic_vector(32472, 16),
63109 => conv_std_logic_vector(32718, 16),
63110 => conv_std_logic_vector(32964, 16),
63111 => conv_std_logic_vector(33210, 16),
63112 => conv_std_logic_vector(33456, 16),
63113 => conv_std_logic_vector(33702, 16),
63114 => conv_std_logic_vector(33948, 16),
63115 => conv_std_logic_vector(34194, 16),
63116 => conv_std_logic_vector(34440, 16),
63117 => conv_std_logic_vector(34686, 16),
63118 => conv_std_logic_vector(34932, 16),
63119 => conv_std_logic_vector(35178, 16),
63120 => conv_std_logic_vector(35424, 16),
63121 => conv_std_logic_vector(35670, 16),
63122 => conv_std_logic_vector(35916, 16),
63123 => conv_std_logic_vector(36162, 16),
63124 => conv_std_logic_vector(36408, 16),
63125 => conv_std_logic_vector(36654, 16),
63126 => conv_std_logic_vector(36900, 16),
63127 => conv_std_logic_vector(37146, 16),
63128 => conv_std_logic_vector(37392, 16),
63129 => conv_std_logic_vector(37638, 16),
63130 => conv_std_logic_vector(37884, 16),
63131 => conv_std_logic_vector(38130, 16),
63132 => conv_std_logic_vector(38376, 16),
63133 => conv_std_logic_vector(38622, 16),
63134 => conv_std_logic_vector(38868, 16),
63135 => conv_std_logic_vector(39114, 16),
63136 => conv_std_logic_vector(39360, 16),
63137 => conv_std_logic_vector(39606, 16),
63138 => conv_std_logic_vector(39852, 16),
63139 => conv_std_logic_vector(40098, 16),
63140 => conv_std_logic_vector(40344, 16),
63141 => conv_std_logic_vector(40590, 16),
63142 => conv_std_logic_vector(40836, 16),
63143 => conv_std_logic_vector(41082, 16),
63144 => conv_std_logic_vector(41328, 16),
63145 => conv_std_logic_vector(41574, 16),
63146 => conv_std_logic_vector(41820, 16),
63147 => conv_std_logic_vector(42066, 16),
63148 => conv_std_logic_vector(42312, 16),
63149 => conv_std_logic_vector(42558, 16),
63150 => conv_std_logic_vector(42804, 16),
63151 => conv_std_logic_vector(43050, 16),
63152 => conv_std_logic_vector(43296, 16),
63153 => conv_std_logic_vector(43542, 16),
63154 => conv_std_logic_vector(43788, 16),
63155 => conv_std_logic_vector(44034, 16),
63156 => conv_std_logic_vector(44280, 16),
63157 => conv_std_logic_vector(44526, 16),
63158 => conv_std_logic_vector(44772, 16),
63159 => conv_std_logic_vector(45018, 16),
63160 => conv_std_logic_vector(45264, 16),
63161 => conv_std_logic_vector(45510, 16),
63162 => conv_std_logic_vector(45756, 16),
63163 => conv_std_logic_vector(46002, 16),
63164 => conv_std_logic_vector(46248, 16),
63165 => conv_std_logic_vector(46494, 16),
63166 => conv_std_logic_vector(46740, 16),
63167 => conv_std_logic_vector(46986, 16),
63168 => conv_std_logic_vector(47232, 16),
63169 => conv_std_logic_vector(47478, 16),
63170 => conv_std_logic_vector(47724, 16),
63171 => conv_std_logic_vector(47970, 16),
63172 => conv_std_logic_vector(48216, 16),
63173 => conv_std_logic_vector(48462, 16),
63174 => conv_std_logic_vector(48708, 16),
63175 => conv_std_logic_vector(48954, 16),
63176 => conv_std_logic_vector(49200, 16),
63177 => conv_std_logic_vector(49446, 16),
63178 => conv_std_logic_vector(49692, 16),
63179 => conv_std_logic_vector(49938, 16),
63180 => conv_std_logic_vector(50184, 16),
63181 => conv_std_logic_vector(50430, 16),
63182 => conv_std_logic_vector(50676, 16),
63183 => conv_std_logic_vector(50922, 16),
63184 => conv_std_logic_vector(51168, 16),
63185 => conv_std_logic_vector(51414, 16),
63186 => conv_std_logic_vector(51660, 16),
63187 => conv_std_logic_vector(51906, 16),
63188 => conv_std_logic_vector(52152, 16),
63189 => conv_std_logic_vector(52398, 16),
63190 => conv_std_logic_vector(52644, 16),
63191 => conv_std_logic_vector(52890, 16),
63192 => conv_std_logic_vector(53136, 16),
63193 => conv_std_logic_vector(53382, 16),
63194 => conv_std_logic_vector(53628, 16),
63195 => conv_std_logic_vector(53874, 16),
63196 => conv_std_logic_vector(54120, 16),
63197 => conv_std_logic_vector(54366, 16),
63198 => conv_std_logic_vector(54612, 16),
63199 => conv_std_logic_vector(54858, 16),
63200 => conv_std_logic_vector(55104, 16),
63201 => conv_std_logic_vector(55350, 16),
63202 => conv_std_logic_vector(55596, 16),
63203 => conv_std_logic_vector(55842, 16),
63204 => conv_std_logic_vector(56088, 16),
63205 => conv_std_logic_vector(56334, 16),
63206 => conv_std_logic_vector(56580, 16),
63207 => conv_std_logic_vector(56826, 16),
63208 => conv_std_logic_vector(57072, 16),
63209 => conv_std_logic_vector(57318, 16),
63210 => conv_std_logic_vector(57564, 16),
63211 => conv_std_logic_vector(57810, 16),
63212 => conv_std_logic_vector(58056, 16),
63213 => conv_std_logic_vector(58302, 16),
63214 => conv_std_logic_vector(58548, 16),
63215 => conv_std_logic_vector(58794, 16),
63216 => conv_std_logic_vector(59040, 16),
63217 => conv_std_logic_vector(59286, 16),
63218 => conv_std_logic_vector(59532, 16),
63219 => conv_std_logic_vector(59778, 16),
63220 => conv_std_logic_vector(60024, 16),
63221 => conv_std_logic_vector(60270, 16),
63222 => conv_std_logic_vector(60516, 16),
63223 => conv_std_logic_vector(60762, 16),
63224 => conv_std_logic_vector(61008, 16),
63225 => conv_std_logic_vector(61254, 16),
63226 => conv_std_logic_vector(61500, 16),
63227 => conv_std_logic_vector(61746, 16),
63228 => conv_std_logic_vector(61992, 16),
63229 => conv_std_logic_vector(62238, 16),
63230 => conv_std_logic_vector(62484, 16),
63231 => conv_std_logic_vector(62730, 16),
63232 => conv_std_logic_vector(0, 16),
63233 => conv_std_logic_vector(247, 16),
63234 => conv_std_logic_vector(494, 16),
63235 => conv_std_logic_vector(741, 16),
63236 => conv_std_logic_vector(988, 16),
63237 => conv_std_logic_vector(1235, 16),
63238 => conv_std_logic_vector(1482, 16),
63239 => conv_std_logic_vector(1729, 16),
63240 => conv_std_logic_vector(1976, 16),
63241 => conv_std_logic_vector(2223, 16),
63242 => conv_std_logic_vector(2470, 16),
63243 => conv_std_logic_vector(2717, 16),
63244 => conv_std_logic_vector(2964, 16),
63245 => conv_std_logic_vector(3211, 16),
63246 => conv_std_logic_vector(3458, 16),
63247 => conv_std_logic_vector(3705, 16),
63248 => conv_std_logic_vector(3952, 16),
63249 => conv_std_logic_vector(4199, 16),
63250 => conv_std_logic_vector(4446, 16),
63251 => conv_std_logic_vector(4693, 16),
63252 => conv_std_logic_vector(4940, 16),
63253 => conv_std_logic_vector(5187, 16),
63254 => conv_std_logic_vector(5434, 16),
63255 => conv_std_logic_vector(5681, 16),
63256 => conv_std_logic_vector(5928, 16),
63257 => conv_std_logic_vector(6175, 16),
63258 => conv_std_logic_vector(6422, 16),
63259 => conv_std_logic_vector(6669, 16),
63260 => conv_std_logic_vector(6916, 16),
63261 => conv_std_logic_vector(7163, 16),
63262 => conv_std_logic_vector(7410, 16),
63263 => conv_std_logic_vector(7657, 16),
63264 => conv_std_logic_vector(7904, 16),
63265 => conv_std_logic_vector(8151, 16),
63266 => conv_std_logic_vector(8398, 16),
63267 => conv_std_logic_vector(8645, 16),
63268 => conv_std_logic_vector(8892, 16),
63269 => conv_std_logic_vector(9139, 16),
63270 => conv_std_logic_vector(9386, 16),
63271 => conv_std_logic_vector(9633, 16),
63272 => conv_std_logic_vector(9880, 16),
63273 => conv_std_logic_vector(10127, 16),
63274 => conv_std_logic_vector(10374, 16),
63275 => conv_std_logic_vector(10621, 16),
63276 => conv_std_logic_vector(10868, 16),
63277 => conv_std_logic_vector(11115, 16),
63278 => conv_std_logic_vector(11362, 16),
63279 => conv_std_logic_vector(11609, 16),
63280 => conv_std_logic_vector(11856, 16),
63281 => conv_std_logic_vector(12103, 16),
63282 => conv_std_logic_vector(12350, 16),
63283 => conv_std_logic_vector(12597, 16),
63284 => conv_std_logic_vector(12844, 16),
63285 => conv_std_logic_vector(13091, 16),
63286 => conv_std_logic_vector(13338, 16),
63287 => conv_std_logic_vector(13585, 16),
63288 => conv_std_logic_vector(13832, 16),
63289 => conv_std_logic_vector(14079, 16),
63290 => conv_std_logic_vector(14326, 16),
63291 => conv_std_logic_vector(14573, 16),
63292 => conv_std_logic_vector(14820, 16),
63293 => conv_std_logic_vector(15067, 16),
63294 => conv_std_logic_vector(15314, 16),
63295 => conv_std_logic_vector(15561, 16),
63296 => conv_std_logic_vector(15808, 16),
63297 => conv_std_logic_vector(16055, 16),
63298 => conv_std_logic_vector(16302, 16),
63299 => conv_std_logic_vector(16549, 16),
63300 => conv_std_logic_vector(16796, 16),
63301 => conv_std_logic_vector(17043, 16),
63302 => conv_std_logic_vector(17290, 16),
63303 => conv_std_logic_vector(17537, 16),
63304 => conv_std_logic_vector(17784, 16),
63305 => conv_std_logic_vector(18031, 16),
63306 => conv_std_logic_vector(18278, 16),
63307 => conv_std_logic_vector(18525, 16),
63308 => conv_std_logic_vector(18772, 16),
63309 => conv_std_logic_vector(19019, 16),
63310 => conv_std_logic_vector(19266, 16),
63311 => conv_std_logic_vector(19513, 16),
63312 => conv_std_logic_vector(19760, 16),
63313 => conv_std_logic_vector(20007, 16),
63314 => conv_std_logic_vector(20254, 16),
63315 => conv_std_logic_vector(20501, 16),
63316 => conv_std_logic_vector(20748, 16),
63317 => conv_std_logic_vector(20995, 16),
63318 => conv_std_logic_vector(21242, 16),
63319 => conv_std_logic_vector(21489, 16),
63320 => conv_std_logic_vector(21736, 16),
63321 => conv_std_logic_vector(21983, 16),
63322 => conv_std_logic_vector(22230, 16),
63323 => conv_std_logic_vector(22477, 16),
63324 => conv_std_logic_vector(22724, 16),
63325 => conv_std_logic_vector(22971, 16),
63326 => conv_std_logic_vector(23218, 16),
63327 => conv_std_logic_vector(23465, 16),
63328 => conv_std_logic_vector(23712, 16),
63329 => conv_std_logic_vector(23959, 16),
63330 => conv_std_logic_vector(24206, 16),
63331 => conv_std_logic_vector(24453, 16),
63332 => conv_std_logic_vector(24700, 16),
63333 => conv_std_logic_vector(24947, 16),
63334 => conv_std_logic_vector(25194, 16),
63335 => conv_std_logic_vector(25441, 16),
63336 => conv_std_logic_vector(25688, 16),
63337 => conv_std_logic_vector(25935, 16),
63338 => conv_std_logic_vector(26182, 16),
63339 => conv_std_logic_vector(26429, 16),
63340 => conv_std_logic_vector(26676, 16),
63341 => conv_std_logic_vector(26923, 16),
63342 => conv_std_logic_vector(27170, 16),
63343 => conv_std_logic_vector(27417, 16),
63344 => conv_std_logic_vector(27664, 16),
63345 => conv_std_logic_vector(27911, 16),
63346 => conv_std_logic_vector(28158, 16),
63347 => conv_std_logic_vector(28405, 16),
63348 => conv_std_logic_vector(28652, 16),
63349 => conv_std_logic_vector(28899, 16),
63350 => conv_std_logic_vector(29146, 16),
63351 => conv_std_logic_vector(29393, 16),
63352 => conv_std_logic_vector(29640, 16),
63353 => conv_std_logic_vector(29887, 16),
63354 => conv_std_logic_vector(30134, 16),
63355 => conv_std_logic_vector(30381, 16),
63356 => conv_std_logic_vector(30628, 16),
63357 => conv_std_logic_vector(30875, 16),
63358 => conv_std_logic_vector(31122, 16),
63359 => conv_std_logic_vector(31369, 16),
63360 => conv_std_logic_vector(31616, 16),
63361 => conv_std_logic_vector(31863, 16),
63362 => conv_std_logic_vector(32110, 16),
63363 => conv_std_logic_vector(32357, 16),
63364 => conv_std_logic_vector(32604, 16),
63365 => conv_std_logic_vector(32851, 16),
63366 => conv_std_logic_vector(33098, 16),
63367 => conv_std_logic_vector(33345, 16),
63368 => conv_std_logic_vector(33592, 16),
63369 => conv_std_logic_vector(33839, 16),
63370 => conv_std_logic_vector(34086, 16),
63371 => conv_std_logic_vector(34333, 16),
63372 => conv_std_logic_vector(34580, 16),
63373 => conv_std_logic_vector(34827, 16),
63374 => conv_std_logic_vector(35074, 16),
63375 => conv_std_logic_vector(35321, 16),
63376 => conv_std_logic_vector(35568, 16),
63377 => conv_std_logic_vector(35815, 16),
63378 => conv_std_logic_vector(36062, 16),
63379 => conv_std_logic_vector(36309, 16),
63380 => conv_std_logic_vector(36556, 16),
63381 => conv_std_logic_vector(36803, 16),
63382 => conv_std_logic_vector(37050, 16),
63383 => conv_std_logic_vector(37297, 16),
63384 => conv_std_logic_vector(37544, 16),
63385 => conv_std_logic_vector(37791, 16),
63386 => conv_std_logic_vector(38038, 16),
63387 => conv_std_logic_vector(38285, 16),
63388 => conv_std_logic_vector(38532, 16),
63389 => conv_std_logic_vector(38779, 16),
63390 => conv_std_logic_vector(39026, 16),
63391 => conv_std_logic_vector(39273, 16),
63392 => conv_std_logic_vector(39520, 16),
63393 => conv_std_logic_vector(39767, 16),
63394 => conv_std_logic_vector(40014, 16),
63395 => conv_std_logic_vector(40261, 16),
63396 => conv_std_logic_vector(40508, 16),
63397 => conv_std_logic_vector(40755, 16),
63398 => conv_std_logic_vector(41002, 16),
63399 => conv_std_logic_vector(41249, 16),
63400 => conv_std_logic_vector(41496, 16),
63401 => conv_std_logic_vector(41743, 16),
63402 => conv_std_logic_vector(41990, 16),
63403 => conv_std_logic_vector(42237, 16),
63404 => conv_std_logic_vector(42484, 16),
63405 => conv_std_logic_vector(42731, 16),
63406 => conv_std_logic_vector(42978, 16),
63407 => conv_std_logic_vector(43225, 16),
63408 => conv_std_logic_vector(43472, 16),
63409 => conv_std_logic_vector(43719, 16),
63410 => conv_std_logic_vector(43966, 16),
63411 => conv_std_logic_vector(44213, 16),
63412 => conv_std_logic_vector(44460, 16),
63413 => conv_std_logic_vector(44707, 16),
63414 => conv_std_logic_vector(44954, 16),
63415 => conv_std_logic_vector(45201, 16),
63416 => conv_std_logic_vector(45448, 16),
63417 => conv_std_logic_vector(45695, 16),
63418 => conv_std_logic_vector(45942, 16),
63419 => conv_std_logic_vector(46189, 16),
63420 => conv_std_logic_vector(46436, 16),
63421 => conv_std_logic_vector(46683, 16),
63422 => conv_std_logic_vector(46930, 16),
63423 => conv_std_logic_vector(47177, 16),
63424 => conv_std_logic_vector(47424, 16),
63425 => conv_std_logic_vector(47671, 16),
63426 => conv_std_logic_vector(47918, 16),
63427 => conv_std_logic_vector(48165, 16),
63428 => conv_std_logic_vector(48412, 16),
63429 => conv_std_logic_vector(48659, 16),
63430 => conv_std_logic_vector(48906, 16),
63431 => conv_std_logic_vector(49153, 16),
63432 => conv_std_logic_vector(49400, 16),
63433 => conv_std_logic_vector(49647, 16),
63434 => conv_std_logic_vector(49894, 16),
63435 => conv_std_logic_vector(50141, 16),
63436 => conv_std_logic_vector(50388, 16),
63437 => conv_std_logic_vector(50635, 16),
63438 => conv_std_logic_vector(50882, 16),
63439 => conv_std_logic_vector(51129, 16),
63440 => conv_std_logic_vector(51376, 16),
63441 => conv_std_logic_vector(51623, 16),
63442 => conv_std_logic_vector(51870, 16),
63443 => conv_std_logic_vector(52117, 16),
63444 => conv_std_logic_vector(52364, 16),
63445 => conv_std_logic_vector(52611, 16),
63446 => conv_std_logic_vector(52858, 16),
63447 => conv_std_logic_vector(53105, 16),
63448 => conv_std_logic_vector(53352, 16),
63449 => conv_std_logic_vector(53599, 16),
63450 => conv_std_logic_vector(53846, 16),
63451 => conv_std_logic_vector(54093, 16),
63452 => conv_std_logic_vector(54340, 16),
63453 => conv_std_logic_vector(54587, 16),
63454 => conv_std_logic_vector(54834, 16),
63455 => conv_std_logic_vector(55081, 16),
63456 => conv_std_logic_vector(55328, 16),
63457 => conv_std_logic_vector(55575, 16),
63458 => conv_std_logic_vector(55822, 16),
63459 => conv_std_logic_vector(56069, 16),
63460 => conv_std_logic_vector(56316, 16),
63461 => conv_std_logic_vector(56563, 16),
63462 => conv_std_logic_vector(56810, 16),
63463 => conv_std_logic_vector(57057, 16),
63464 => conv_std_logic_vector(57304, 16),
63465 => conv_std_logic_vector(57551, 16),
63466 => conv_std_logic_vector(57798, 16),
63467 => conv_std_logic_vector(58045, 16),
63468 => conv_std_logic_vector(58292, 16),
63469 => conv_std_logic_vector(58539, 16),
63470 => conv_std_logic_vector(58786, 16),
63471 => conv_std_logic_vector(59033, 16),
63472 => conv_std_logic_vector(59280, 16),
63473 => conv_std_logic_vector(59527, 16),
63474 => conv_std_logic_vector(59774, 16),
63475 => conv_std_logic_vector(60021, 16),
63476 => conv_std_logic_vector(60268, 16),
63477 => conv_std_logic_vector(60515, 16),
63478 => conv_std_logic_vector(60762, 16),
63479 => conv_std_logic_vector(61009, 16),
63480 => conv_std_logic_vector(61256, 16),
63481 => conv_std_logic_vector(61503, 16),
63482 => conv_std_logic_vector(61750, 16),
63483 => conv_std_logic_vector(61997, 16),
63484 => conv_std_logic_vector(62244, 16),
63485 => conv_std_logic_vector(62491, 16),
63486 => conv_std_logic_vector(62738, 16),
63487 => conv_std_logic_vector(62985, 16),
63488 => conv_std_logic_vector(0, 16),
63489 => conv_std_logic_vector(248, 16),
63490 => conv_std_logic_vector(496, 16),
63491 => conv_std_logic_vector(744, 16),
63492 => conv_std_logic_vector(992, 16),
63493 => conv_std_logic_vector(1240, 16),
63494 => conv_std_logic_vector(1488, 16),
63495 => conv_std_logic_vector(1736, 16),
63496 => conv_std_logic_vector(1984, 16),
63497 => conv_std_logic_vector(2232, 16),
63498 => conv_std_logic_vector(2480, 16),
63499 => conv_std_logic_vector(2728, 16),
63500 => conv_std_logic_vector(2976, 16),
63501 => conv_std_logic_vector(3224, 16),
63502 => conv_std_logic_vector(3472, 16),
63503 => conv_std_logic_vector(3720, 16),
63504 => conv_std_logic_vector(3968, 16),
63505 => conv_std_logic_vector(4216, 16),
63506 => conv_std_logic_vector(4464, 16),
63507 => conv_std_logic_vector(4712, 16),
63508 => conv_std_logic_vector(4960, 16),
63509 => conv_std_logic_vector(5208, 16),
63510 => conv_std_logic_vector(5456, 16),
63511 => conv_std_logic_vector(5704, 16),
63512 => conv_std_logic_vector(5952, 16),
63513 => conv_std_logic_vector(6200, 16),
63514 => conv_std_logic_vector(6448, 16),
63515 => conv_std_logic_vector(6696, 16),
63516 => conv_std_logic_vector(6944, 16),
63517 => conv_std_logic_vector(7192, 16),
63518 => conv_std_logic_vector(7440, 16),
63519 => conv_std_logic_vector(7688, 16),
63520 => conv_std_logic_vector(7936, 16),
63521 => conv_std_logic_vector(8184, 16),
63522 => conv_std_logic_vector(8432, 16),
63523 => conv_std_logic_vector(8680, 16),
63524 => conv_std_logic_vector(8928, 16),
63525 => conv_std_logic_vector(9176, 16),
63526 => conv_std_logic_vector(9424, 16),
63527 => conv_std_logic_vector(9672, 16),
63528 => conv_std_logic_vector(9920, 16),
63529 => conv_std_logic_vector(10168, 16),
63530 => conv_std_logic_vector(10416, 16),
63531 => conv_std_logic_vector(10664, 16),
63532 => conv_std_logic_vector(10912, 16),
63533 => conv_std_logic_vector(11160, 16),
63534 => conv_std_logic_vector(11408, 16),
63535 => conv_std_logic_vector(11656, 16),
63536 => conv_std_logic_vector(11904, 16),
63537 => conv_std_logic_vector(12152, 16),
63538 => conv_std_logic_vector(12400, 16),
63539 => conv_std_logic_vector(12648, 16),
63540 => conv_std_logic_vector(12896, 16),
63541 => conv_std_logic_vector(13144, 16),
63542 => conv_std_logic_vector(13392, 16),
63543 => conv_std_logic_vector(13640, 16),
63544 => conv_std_logic_vector(13888, 16),
63545 => conv_std_logic_vector(14136, 16),
63546 => conv_std_logic_vector(14384, 16),
63547 => conv_std_logic_vector(14632, 16),
63548 => conv_std_logic_vector(14880, 16),
63549 => conv_std_logic_vector(15128, 16),
63550 => conv_std_logic_vector(15376, 16),
63551 => conv_std_logic_vector(15624, 16),
63552 => conv_std_logic_vector(15872, 16),
63553 => conv_std_logic_vector(16120, 16),
63554 => conv_std_logic_vector(16368, 16),
63555 => conv_std_logic_vector(16616, 16),
63556 => conv_std_logic_vector(16864, 16),
63557 => conv_std_logic_vector(17112, 16),
63558 => conv_std_logic_vector(17360, 16),
63559 => conv_std_logic_vector(17608, 16),
63560 => conv_std_logic_vector(17856, 16),
63561 => conv_std_logic_vector(18104, 16),
63562 => conv_std_logic_vector(18352, 16),
63563 => conv_std_logic_vector(18600, 16),
63564 => conv_std_logic_vector(18848, 16),
63565 => conv_std_logic_vector(19096, 16),
63566 => conv_std_logic_vector(19344, 16),
63567 => conv_std_logic_vector(19592, 16),
63568 => conv_std_logic_vector(19840, 16),
63569 => conv_std_logic_vector(20088, 16),
63570 => conv_std_logic_vector(20336, 16),
63571 => conv_std_logic_vector(20584, 16),
63572 => conv_std_logic_vector(20832, 16),
63573 => conv_std_logic_vector(21080, 16),
63574 => conv_std_logic_vector(21328, 16),
63575 => conv_std_logic_vector(21576, 16),
63576 => conv_std_logic_vector(21824, 16),
63577 => conv_std_logic_vector(22072, 16),
63578 => conv_std_logic_vector(22320, 16),
63579 => conv_std_logic_vector(22568, 16),
63580 => conv_std_logic_vector(22816, 16),
63581 => conv_std_logic_vector(23064, 16),
63582 => conv_std_logic_vector(23312, 16),
63583 => conv_std_logic_vector(23560, 16),
63584 => conv_std_logic_vector(23808, 16),
63585 => conv_std_logic_vector(24056, 16),
63586 => conv_std_logic_vector(24304, 16),
63587 => conv_std_logic_vector(24552, 16),
63588 => conv_std_logic_vector(24800, 16),
63589 => conv_std_logic_vector(25048, 16),
63590 => conv_std_logic_vector(25296, 16),
63591 => conv_std_logic_vector(25544, 16),
63592 => conv_std_logic_vector(25792, 16),
63593 => conv_std_logic_vector(26040, 16),
63594 => conv_std_logic_vector(26288, 16),
63595 => conv_std_logic_vector(26536, 16),
63596 => conv_std_logic_vector(26784, 16),
63597 => conv_std_logic_vector(27032, 16),
63598 => conv_std_logic_vector(27280, 16),
63599 => conv_std_logic_vector(27528, 16),
63600 => conv_std_logic_vector(27776, 16),
63601 => conv_std_logic_vector(28024, 16),
63602 => conv_std_logic_vector(28272, 16),
63603 => conv_std_logic_vector(28520, 16),
63604 => conv_std_logic_vector(28768, 16),
63605 => conv_std_logic_vector(29016, 16),
63606 => conv_std_logic_vector(29264, 16),
63607 => conv_std_logic_vector(29512, 16),
63608 => conv_std_logic_vector(29760, 16),
63609 => conv_std_logic_vector(30008, 16),
63610 => conv_std_logic_vector(30256, 16),
63611 => conv_std_logic_vector(30504, 16),
63612 => conv_std_logic_vector(30752, 16),
63613 => conv_std_logic_vector(31000, 16),
63614 => conv_std_logic_vector(31248, 16),
63615 => conv_std_logic_vector(31496, 16),
63616 => conv_std_logic_vector(31744, 16),
63617 => conv_std_logic_vector(31992, 16),
63618 => conv_std_logic_vector(32240, 16),
63619 => conv_std_logic_vector(32488, 16),
63620 => conv_std_logic_vector(32736, 16),
63621 => conv_std_logic_vector(32984, 16),
63622 => conv_std_logic_vector(33232, 16),
63623 => conv_std_logic_vector(33480, 16),
63624 => conv_std_logic_vector(33728, 16),
63625 => conv_std_logic_vector(33976, 16),
63626 => conv_std_logic_vector(34224, 16),
63627 => conv_std_logic_vector(34472, 16),
63628 => conv_std_logic_vector(34720, 16),
63629 => conv_std_logic_vector(34968, 16),
63630 => conv_std_logic_vector(35216, 16),
63631 => conv_std_logic_vector(35464, 16),
63632 => conv_std_logic_vector(35712, 16),
63633 => conv_std_logic_vector(35960, 16),
63634 => conv_std_logic_vector(36208, 16),
63635 => conv_std_logic_vector(36456, 16),
63636 => conv_std_logic_vector(36704, 16),
63637 => conv_std_logic_vector(36952, 16),
63638 => conv_std_logic_vector(37200, 16),
63639 => conv_std_logic_vector(37448, 16),
63640 => conv_std_logic_vector(37696, 16),
63641 => conv_std_logic_vector(37944, 16),
63642 => conv_std_logic_vector(38192, 16),
63643 => conv_std_logic_vector(38440, 16),
63644 => conv_std_logic_vector(38688, 16),
63645 => conv_std_logic_vector(38936, 16),
63646 => conv_std_logic_vector(39184, 16),
63647 => conv_std_logic_vector(39432, 16),
63648 => conv_std_logic_vector(39680, 16),
63649 => conv_std_logic_vector(39928, 16),
63650 => conv_std_logic_vector(40176, 16),
63651 => conv_std_logic_vector(40424, 16),
63652 => conv_std_logic_vector(40672, 16),
63653 => conv_std_logic_vector(40920, 16),
63654 => conv_std_logic_vector(41168, 16),
63655 => conv_std_logic_vector(41416, 16),
63656 => conv_std_logic_vector(41664, 16),
63657 => conv_std_logic_vector(41912, 16),
63658 => conv_std_logic_vector(42160, 16),
63659 => conv_std_logic_vector(42408, 16),
63660 => conv_std_logic_vector(42656, 16),
63661 => conv_std_logic_vector(42904, 16),
63662 => conv_std_logic_vector(43152, 16),
63663 => conv_std_logic_vector(43400, 16),
63664 => conv_std_logic_vector(43648, 16),
63665 => conv_std_logic_vector(43896, 16),
63666 => conv_std_logic_vector(44144, 16),
63667 => conv_std_logic_vector(44392, 16),
63668 => conv_std_logic_vector(44640, 16),
63669 => conv_std_logic_vector(44888, 16),
63670 => conv_std_logic_vector(45136, 16),
63671 => conv_std_logic_vector(45384, 16),
63672 => conv_std_logic_vector(45632, 16),
63673 => conv_std_logic_vector(45880, 16),
63674 => conv_std_logic_vector(46128, 16),
63675 => conv_std_logic_vector(46376, 16),
63676 => conv_std_logic_vector(46624, 16),
63677 => conv_std_logic_vector(46872, 16),
63678 => conv_std_logic_vector(47120, 16),
63679 => conv_std_logic_vector(47368, 16),
63680 => conv_std_logic_vector(47616, 16),
63681 => conv_std_logic_vector(47864, 16),
63682 => conv_std_logic_vector(48112, 16),
63683 => conv_std_logic_vector(48360, 16),
63684 => conv_std_logic_vector(48608, 16),
63685 => conv_std_logic_vector(48856, 16),
63686 => conv_std_logic_vector(49104, 16),
63687 => conv_std_logic_vector(49352, 16),
63688 => conv_std_logic_vector(49600, 16),
63689 => conv_std_logic_vector(49848, 16),
63690 => conv_std_logic_vector(50096, 16),
63691 => conv_std_logic_vector(50344, 16),
63692 => conv_std_logic_vector(50592, 16),
63693 => conv_std_logic_vector(50840, 16),
63694 => conv_std_logic_vector(51088, 16),
63695 => conv_std_logic_vector(51336, 16),
63696 => conv_std_logic_vector(51584, 16),
63697 => conv_std_logic_vector(51832, 16),
63698 => conv_std_logic_vector(52080, 16),
63699 => conv_std_logic_vector(52328, 16),
63700 => conv_std_logic_vector(52576, 16),
63701 => conv_std_logic_vector(52824, 16),
63702 => conv_std_logic_vector(53072, 16),
63703 => conv_std_logic_vector(53320, 16),
63704 => conv_std_logic_vector(53568, 16),
63705 => conv_std_logic_vector(53816, 16),
63706 => conv_std_logic_vector(54064, 16),
63707 => conv_std_logic_vector(54312, 16),
63708 => conv_std_logic_vector(54560, 16),
63709 => conv_std_logic_vector(54808, 16),
63710 => conv_std_logic_vector(55056, 16),
63711 => conv_std_logic_vector(55304, 16),
63712 => conv_std_logic_vector(55552, 16),
63713 => conv_std_logic_vector(55800, 16),
63714 => conv_std_logic_vector(56048, 16),
63715 => conv_std_logic_vector(56296, 16),
63716 => conv_std_logic_vector(56544, 16),
63717 => conv_std_logic_vector(56792, 16),
63718 => conv_std_logic_vector(57040, 16),
63719 => conv_std_logic_vector(57288, 16),
63720 => conv_std_logic_vector(57536, 16),
63721 => conv_std_logic_vector(57784, 16),
63722 => conv_std_logic_vector(58032, 16),
63723 => conv_std_logic_vector(58280, 16),
63724 => conv_std_logic_vector(58528, 16),
63725 => conv_std_logic_vector(58776, 16),
63726 => conv_std_logic_vector(59024, 16),
63727 => conv_std_logic_vector(59272, 16),
63728 => conv_std_logic_vector(59520, 16),
63729 => conv_std_logic_vector(59768, 16),
63730 => conv_std_logic_vector(60016, 16),
63731 => conv_std_logic_vector(60264, 16),
63732 => conv_std_logic_vector(60512, 16),
63733 => conv_std_logic_vector(60760, 16),
63734 => conv_std_logic_vector(61008, 16),
63735 => conv_std_logic_vector(61256, 16),
63736 => conv_std_logic_vector(61504, 16),
63737 => conv_std_logic_vector(61752, 16),
63738 => conv_std_logic_vector(62000, 16),
63739 => conv_std_logic_vector(62248, 16),
63740 => conv_std_logic_vector(62496, 16),
63741 => conv_std_logic_vector(62744, 16),
63742 => conv_std_logic_vector(62992, 16),
63743 => conv_std_logic_vector(63240, 16),
63744 => conv_std_logic_vector(0, 16),
63745 => conv_std_logic_vector(249, 16),
63746 => conv_std_logic_vector(498, 16),
63747 => conv_std_logic_vector(747, 16),
63748 => conv_std_logic_vector(996, 16),
63749 => conv_std_logic_vector(1245, 16),
63750 => conv_std_logic_vector(1494, 16),
63751 => conv_std_logic_vector(1743, 16),
63752 => conv_std_logic_vector(1992, 16),
63753 => conv_std_logic_vector(2241, 16),
63754 => conv_std_logic_vector(2490, 16),
63755 => conv_std_logic_vector(2739, 16),
63756 => conv_std_logic_vector(2988, 16),
63757 => conv_std_logic_vector(3237, 16),
63758 => conv_std_logic_vector(3486, 16),
63759 => conv_std_logic_vector(3735, 16),
63760 => conv_std_logic_vector(3984, 16),
63761 => conv_std_logic_vector(4233, 16),
63762 => conv_std_logic_vector(4482, 16),
63763 => conv_std_logic_vector(4731, 16),
63764 => conv_std_logic_vector(4980, 16),
63765 => conv_std_logic_vector(5229, 16),
63766 => conv_std_logic_vector(5478, 16),
63767 => conv_std_logic_vector(5727, 16),
63768 => conv_std_logic_vector(5976, 16),
63769 => conv_std_logic_vector(6225, 16),
63770 => conv_std_logic_vector(6474, 16),
63771 => conv_std_logic_vector(6723, 16),
63772 => conv_std_logic_vector(6972, 16),
63773 => conv_std_logic_vector(7221, 16),
63774 => conv_std_logic_vector(7470, 16),
63775 => conv_std_logic_vector(7719, 16),
63776 => conv_std_logic_vector(7968, 16),
63777 => conv_std_logic_vector(8217, 16),
63778 => conv_std_logic_vector(8466, 16),
63779 => conv_std_logic_vector(8715, 16),
63780 => conv_std_logic_vector(8964, 16),
63781 => conv_std_logic_vector(9213, 16),
63782 => conv_std_logic_vector(9462, 16),
63783 => conv_std_logic_vector(9711, 16),
63784 => conv_std_logic_vector(9960, 16),
63785 => conv_std_logic_vector(10209, 16),
63786 => conv_std_logic_vector(10458, 16),
63787 => conv_std_logic_vector(10707, 16),
63788 => conv_std_logic_vector(10956, 16),
63789 => conv_std_logic_vector(11205, 16),
63790 => conv_std_logic_vector(11454, 16),
63791 => conv_std_logic_vector(11703, 16),
63792 => conv_std_logic_vector(11952, 16),
63793 => conv_std_logic_vector(12201, 16),
63794 => conv_std_logic_vector(12450, 16),
63795 => conv_std_logic_vector(12699, 16),
63796 => conv_std_logic_vector(12948, 16),
63797 => conv_std_logic_vector(13197, 16),
63798 => conv_std_logic_vector(13446, 16),
63799 => conv_std_logic_vector(13695, 16),
63800 => conv_std_logic_vector(13944, 16),
63801 => conv_std_logic_vector(14193, 16),
63802 => conv_std_logic_vector(14442, 16),
63803 => conv_std_logic_vector(14691, 16),
63804 => conv_std_logic_vector(14940, 16),
63805 => conv_std_logic_vector(15189, 16),
63806 => conv_std_logic_vector(15438, 16),
63807 => conv_std_logic_vector(15687, 16),
63808 => conv_std_logic_vector(15936, 16),
63809 => conv_std_logic_vector(16185, 16),
63810 => conv_std_logic_vector(16434, 16),
63811 => conv_std_logic_vector(16683, 16),
63812 => conv_std_logic_vector(16932, 16),
63813 => conv_std_logic_vector(17181, 16),
63814 => conv_std_logic_vector(17430, 16),
63815 => conv_std_logic_vector(17679, 16),
63816 => conv_std_logic_vector(17928, 16),
63817 => conv_std_logic_vector(18177, 16),
63818 => conv_std_logic_vector(18426, 16),
63819 => conv_std_logic_vector(18675, 16),
63820 => conv_std_logic_vector(18924, 16),
63821 => conv_std_logic_vector(19173, 16),
63822 => conv_std_logic_vector(19422, 16),
63823 => conv_std_logic_vector(19671, 16),
63824 => conv_std_logic_vector(19920, 16),
63825 => conv_std_logic_vector(20169, 16),
63826 => conv_std_logic_vector(20418, 16),
63827 => conv_std_logic_vector(20667, 16),
63828 => conv_std_logic_vector(20916, 16),
63829 => conv_std_logic_vector(21165, 16),
63830 => conv_std_logic_vector(21414, 16),
63831 => conv_std_logic_vector(21663, 16),
63832 => conv_std_logic_vector(21912, 16),
63833 => conv_std_logic_vector(22161, 16),
63834 => conv_std_logic_vector(22410, 16),
63835 => conv_std_logic_vector(22659, 16),
63836 => conv_std_logic_vector(22908, 16),
63837 => conv_std_logic_vector(23157, 16),
63838 => conv_std_logic_vector(23406, 16),
63839 => conv_std_logic_vector(23655, 16),
63840 => conv_std_logic_vector(23904, 16),
63841 => conv_std_logic_vector(24153, 16),
63842 => conv_std_logic_vector(24402, 16),
63843 => conv_std_logic_vector(24651, 16),
63844 => conv_std_logic_vector(24900, 16),
63845 => conv_std_logic_vector(25149, 16),
63846 => conv_std_logic_vector(25398, 16),
63847 => conv_std_logic_vector(25647, 16),
63848 => conv_std_logic_vector(25896, 16),
63849 => conv_std_logic_vector(26145, 16),
63850 => conv_std_logic_vector(26394, 16),
63851 => conv_std_logic_vector(26643, 16),
63852 => conv_std_logic_vector(26892, 16),
63853 => conv_std_logic_vector(27141, 16),
63854 => conv_std_logic_vector(27390, 16),
63855 => conv_std_logic_vector(27639, 16),
63856 => conv_std_logic_vector(27888, 16),
63857 => conv_std_logic_vector(28137, 16),
63858 => conv_std_logic_vector(28386, 16),
63859 => conv_std_logic_vector(28635, 16),
63860 => conv_std_logic_vector(28884, 16),
63861 => conv_std_logic_vector(29133, 16),
63862 => conv_std_logic_vector(29382, 16),
63863 => conv_std_logic_vector(29631, 16),
63864 => conv_std_logic_vector(29880, 16),
63865 => conv_std_logic_vector(30129, 16),
63866 => conv_std_logic_vector(30378, 16),
63867 => conv_std_logic_vector(30627, 16),
63868 => conv_std_logic_vector(30876, 16),
63869 => conv_std_logic_vector(31125, 16),
63870 => conv_std_logic_vector(31374, 16),
63871 => conv_std_logic_vector(31623, 16),
63872 => conv_std_logic_vector(31872, 16),
63873 => conv_std_logic_vector(32121, 16),
63874 => conv_std_logic_vector(32370, 16),
63875 => conv_std_logic_vector(32619, 16),
63876 => conv_std_logic_vector(32868, 16),
63877 => conv_std_logic_vector(33117, 16),
63878 => conv_std_logic_vector(33366, 16),
63879 => conv_std_logic_vector(33615, 16),
63880 => conv_std_logic_vector(33864, 16),
63881 => conv_std_logic_vector(34113, 16),
63882 => conv_std_logic_vector(34362, 16),
63883 => conv_std_logic_vector(34611, 16),
63884 => conv_std_logic_vector(34860, 16),
63885 => conv_std_logic_vector(35109, 16),
63886 => conv_std_logic_vector(35358, 16),
63887 => conv_std_logic_vector(35607, 16),
63888 => conv_std_logic_vector(35856, 16),
63889 => conv_std_logic_vector(36105, 16),
63890 => conv_std_logic_vector(36354, 16),
63891 => conv_std_logic_vector(36603, 16),
63892 => conv_std_logic_vector(36852, 16),
63893 => conv_std_logic_vector(37101, 16),
63894 => conv_std_logic_vector(37350, 16),
63895 => conv_std_logic_vector(37599, 16),
63896 => conv_std_logic_vector(37848, 16),
63897 => conv_std_logic_vector(38097, 16),
63898 => conv_std_logic_vector(38346, 16),
63899 => conv_std_logic_vector(38595, 16),
63900 => conv_std_logic_vector(38844, 16),
63901 => conv_std_logic_vector(39093, 16),
63902 => conv_std_logic_vector(39342, 16),
63903 => conv_std_logic_vector(39591, 16),
63904 => conv_std_logic_vector(39840, 16),
63905 => conv_std_logic_vector(40089, 16),
63906 => conv_std_logic_vector(40338, 16),
63907 => conv_std_logic_vector(40587, 16),
63908 => conv_std_logic_vector(40836, 16),
63909 => conv_std_logic_vector(41085, 16),
63910 => conv_std_logic_vector(41334, 16),
63911 => conv_std_logic_vector(41583, 16),
63912 => conv_std_logic_vector(41832, 16),
63913 => conv_std_logic_vector(42081, 16),
63914 => conv_std_logic_vector(42330, 16),
63915 => conv_std_logic_vector(42579, 16),
63916 => conv_std_logic_vector(42828, 16),
63917 => conv_std_logic_vector(43077, 16),
63918 => conv_std_logic_vector(43326, 16),
63919 => conv_std_logic_vector(43575, 16),
63920 => conv_std_logic_vector(43824, 16),
63921 => conv_std_logic_vector(44073, 16),
63922 => conv_std_logic_vector(44322, 16),
63923 => conv_std_logic_vector(44571, 16),
63924 => conv_std_logic_vector(44820, 16),
63925 => conv_std_logic_vector(45069, 16),
63926 => conv_std_logic_vector(45318, 16),
63927 => conv_std_logic_vector(45567, 16),
63928 => conv_std_logic_vector(45816, 16),
63929 => conv_std_logic_vector(46065, 16),
63930 => conv_std_logic_vector(46314, 16),
63931 => conv_std_logic_vector(46563, 16),
63932 => conv_std_logic_vector(46812, 16),
63933 => conv_std_logic_vector(47061, 16),
63934 => conv_std_logic_vector(47310, 16),
63935 => conv_std_logic_vector(47559, 16),
63936 => conv_std_logic_vector(47808, 16),
63937 => conv_std_logic_vector(48057, 16),
63938 => conv_std_logic_vector(48306, 16),
63939 => conv_std_logic_vector(48555, 16),
63940 => conv_std_logic_vector(48804, 16),
63941 => conv_std_logic_vector(49053, 16),
63942 => conv_std_logic_vector(49302, 16),
63943 => conv_std_logic_vector(49551, 16),
63944 => conv_std_logic_vector(49800, 16),
63945 => conv_std_logic_vector(50049, 16),
63946 => conv_std_logic_vector(50298, 16),
63947 => conv_std_logic_vector(50547, 16),
63948 => conv_std_logic_vector(50796, 16),
63949 => conv_std_logic_vector(51045, 16),
63950 => conv_std_logic_vector(51294, 16),
63951 => conv_std_logic_vector(51543, 16),
63952 => conv_std_logic_vector(51792, 16),
63953 => conv_std_logic_vector(52041, 16),
63954 => conv_std_logic_vector(52290, 16),
63955 => conv_std_logic_vector(52539, 16),
63956 => conv_std_logic_vector(52788, 16),
63957 => conv_std_logic_vector(53037, 16),
63958 => conv_std_logic_vector(53286, 16),
63959 => conv_std_logic_vector(53535, 16),
63960 => conv_std_logic_vector(53784, 16),
63961 => conv_std_logic_vector(54033, 16),
63962 => conv_std_logic_vector(54282, 16),
63963 => conv_std_logic_vector(54531, 16),
63964 => conv_std_logic_vector(54780, 16),
63965 => conv_std_logic_vector(55029, 16),
63966 => conv_std_logic_vector(55278, 16),
63967 => conv_std_logic_vector(55527, 16),
63968 => conv_std_logic_vector(55776, 16),
63969 => conv_std_logic_vector(56025, 16),
63970 => conv_std_logic_vector(56274, 16),
63971 => conv_std_logic_vector(56523, 16),
63972 => conv_std_logic_vector(56772, 16),
63973 => conv_std_logic_vector(57021, 16),
63974 => conv_std_logic_vector(57270, 16),
63975 => conv_std_logic_vector(57519, 16),
63976 => conv_std_logic_vector(57768, 16),
63977 => conv_std_logic_vector(58017, 16),
63978 => conv_std_logic_vector(58266, 16),
63979 => conv_std_logic_vector(58515, 16),
63980 => conv_std_logic_vector(58764, 16),
63981 => conv_std_logic_vector(59013, 16),
63982 => conv_std_logic_vector(59262, 16),
63983 => conv_std_logic_vector(59511, 16),
63984 => conv_std_logic_vector(59760, 16),
63985 => conv_std_logic_vector(60009, 16),
63986 => conv_std_logic_vector(60258, 16),
63987 => conv_std_logic_vector(60507, 16),
63988 => conv_std_logic_vector(60756, 16),
63989 => conv_std_logic_vector(61005, 16),
63990 => conv_std_logic_vector(61254, 16),
63991 => conv_std_logic_vector(61503, 16),
63992 => conv_std_logic_vector(61752, 16),
63993 => conv_std_logic_vector(62001, 16),
63994 => conv_std_logic_vector(62250, 16),
63995 => conv_std_logic_vector(62499, 16),
63996 => conv_std_logic_vector(62748, 16),
63997 => conv_std_logic_vector(62997, 16),
63998 => conv_std_logic_vector(63246, 16),
63999 => conv_std_logic_vector(63495, 16),
64000 => conv_std_logic_vector(0, 16),
64001 => conv_std_logic_vector(250, 16),
64002 => conv_std_logic_vector(500, 16),
64003 => conv_std_logic_vector(750, 16),
64004 => conv_std_logic_vector(1000, 16),
64005 => conv_std_logic_vector(1250, 16),
64006 => conv_std_logic_vector(1500, 16),
64007 => conv_std_logic_vector(1750, 16),
64008 => conv_std_logic_vector(2000, 16),
64009 => conv_std_logic_vector(2250, 16),
64010 => conv_std_logic_vector(2500, 16),
64011 => conv_std_logic_vector(2750, 16),
64012 => conv_std_logic_vector(3000, 16),
64013 => conv_std_logic_vector(3250, 16),
64014 => conv_std_logic_vector(3500, 16),
64015 => conv_std_logic_vector(3750, 16),
64016 => conv_std_logic_vector(4000, 16),
64017 => conv_std_logic_vector(4250, 16),
64018 => conv_std_logic_vector(4500, 16),
64019 => conv_std_logic_vector(4750, 16),
64020 => conv_std_logic_vector(5000, 16),
64021 => conv_std_logic_vector(5250, 16),
64022 => conv_std_logic_vector(5500, 16),
64023 => conv_std_logic_vector(5750, 16),
64024 => conv_std_logic_vector(6000, 16),
64025 => conv_std_logic_vector(6250, 16),
64026 => conv_std_logic_vector(6500, 16),
64027 => conv_std_logic_vector(6750, 16),
64028 => conv_std_logic_vector(7000, 16),
64029 => conv_std_logic_vector(7250, 16),
64030 => conv_std_logic_vector(7500, 16),
64031 => conv_std_logic_vector(7750, 16),
64032 => conv_std_logic_vector(8000, 16),
64033 => conv_std_logic_vector(8250, 16),
64034 => conv_std_logic_vector(8500, 16),
64035 => conv_std_logic_vector(8750, 16),
64036 => conv_std_logic_vector(9000, 16),
64037 => conv_std_logic_vector(9250, 16),
64038 => conv_std_logic_vector(9500, 16),
64039 => conv_std_logic_vector(9750, 16),
64040 => conv_std_logic_vector(10000, 16),
64041 => conv_std_logic_vector(10250, 16),
64042 => conv_std_logic_vector(10500, 16),
64043 => conv_std_logic_vector(10750, 16),
64044 => conv_std_logic_vector(11000, 16),
64045 => conv_std_logic_vector(11250, 16),
64046 => conv_std_logic_vector(11500, 16),
64047 => conv_std_logic_vector(11750, 16),
64048 => conv_std_logic_vector(12000, 16),
64049 => conv_std_logic_vector(12250, 16),
64050 => conv_std_logic_vector(12500, 16),
64051 => conv_std_logic_vector(12750, 16),
64052 => conv_std_logic_vector(13000, 16),
64053 => conv_std_logic_vector(13250, 16),
64054 => conv_std_logic_vector(13500, 16),
64055 => conv_std_logic_vector(13750, 16),
64056 => conv_std_logic_vector(14000, 16),
64057 => conv_std_logic_vector(14250, 16),
64058 => conv_std_logic_vector(14500, 16),
64059 => conv_std_logic_vector(14750, 16),
64060 => conv_std_logic_vector(15000, 16),
64061 => conv_std_logic_vector(15250, 16),
64062 => conv_std_logic_vector(15500, 16),
64063 => conv_std_logic_vector(15750, 16),
64064 => conv_std_logic_vector(16000, 16),
64065 => conv_std_logic_vector(16250, 16),
64066 => conv_std_logic_vector(16500, 16),
64067 => conv_std_logic_vector(16750, 16),
64068 => conv_std_logic_vector(17000, 16),
64069 => conv_std_logic_vector(17250, 16),
64070 => conv_std_logic_vector(17500, 16),
64071 => conv_std_logic_vector(17750, 16),
64072 => conv_std_logic_vector(18000, 16),
64073 => conv_std_logic_vector(18250, 16),
64074 => conv_std_logic_vector(18500, 16),
64075 => conv_std_logic_vector(18750, 16),
64076 => conv_std_logic_vector(19000, 16),
64077 => conv_std_logic_vector(19250, 16),
64078 => conv_std_logic_vector(19500, 16),
64079 => conv_std_logic_vector(19750, 16),
64080 => conv_std_logic_vector(20000, 16),
64081 => conv_std_logic_vector(20250, 16),
64082 => conv_std_logic_vector(20500, 16),
64083 => conv_std_logic_vector(20750, 16),
64084 => conv_std_logic_vector(21000, 16),
64085 => conv_std_logic_vector(21250, 16),
64086 => conv_std_logic_vector(21500, 16),
64087 => conv_std_logic_vector(21750, 16),
64088 => conv_std_logic_vector(22000, 16),
64089 => conv_std_logic_vector(22250, 16),
64090 => conv_std_logic_vector(22500, 16),
64091 => conv_std_logic_vector(22750, 16),
64092 => conv_std_logic_vector(23000, 16),
64093 => conv_std_logic_vector(23250, 16),
64094 => conv_std_logic_vector(23500, 16),
64095 => conv_std_logic_vector(23750, 16),
64096 => conv_std_logic_vector(24000, 16),
64097 => conv_std_logic_vector(24250, 16),
64098 => conv_std_logic_vector(24500, 16),
64099 => conv_std_logic_vector(24750, 16),
64100 => conv_std_logic_vector(25000, 16),
64101 => conv_std_logic_vector(25250, 16),
64102 => conv_std_logic_vector(25500, 16),
64103 => conv_std_logic_vector(25750, 16),
64104 => conv_std_logic_vector(26000, 16),
64105 => conv_std_logic_vector(26250, 16),
64106 => conv_std_logic_vector(26500, 16),
64107 => conv_std_logic_vector(26750, 16),
64108 => conv_std_logic_vector(27000, 16),
64109 => conv_std_logic_vector(27250, 16),
64110 => conv_std_logic_vector(27500, 16),
64111 => conv_std_logic_vector(27750, 16),
64112 => conv_std_logic_vector(28000, 16),
64113 => conv_std_logic_vector(28250, 16),
64114 => conv_std_logic_vector(28500, 16),
64115 => conv_std_logic_vector(28750, 16),
64116 => conv_std_logic_vector(29000, 16),
64117 => conv_std_logic_vector(29250, 16),
64118 => conv_std_logic_vector(29500, 16),
64119 => conv_std_logic_vector(29750, 16),
64120 => conv_std_logic_vector(30000, 16),
64121 => conv_std_logic_vector(30250, 16),
64122 => conv_std_logic_vector(30500, 16),
64123 => conv_std_logic_vector(30750, 16),
64124 => conv_std_logic_vector(31000, 16),
64125 => conv_std_logic_vector(31250, 16),
64126 => conv_std_logic_vector(31500, 16),
64127 => conv_std_logic_vector(31750, 16),
64128 => conv_std_logic_vector(32000, 16),
64129 => conv_std_logic_vector(32250, 16),
64130 => conv_std_logic_vector(32500, 16),
64131 => conv_std_logic_vector(32750, 16),
64132 => conv_std_logic_vector(33000, 16),
64133 => conv_std_logic_vector(33250, 16),
64134 => conv_std_logic_vector(33500, 16),
64135 => conv_std_logic_vector(33750, 16),
64136 => conv_std_logic_vector(34000, 16),
64137 => conv_std_logic_vector(34250, 16),
64138 => conv_std_logic_vector(34500, 16),
64139 => conv_std_logic_vector(34750, 16),
64140 => conv_std_logic_vector(35000, 16),
64141 => conv_std_logic_vector(35250, 16),
64142 => conv_std_logic_vector(35500, 16),
64143 => conv_std_logic_vector(35750, 16),
64144 => conv_std_logic_vector(36000, 16),
64145 => conv_std_logic_vector(36250, 16),
64146 => conv_std_logic_vector(36500, 16),
64147 => conv_std_logic_vector(36750, 16),
64148 => conv_std_logic_vector(37000, 16),
64149 => conv_std_logic_vector(37250, 16),
64150 => conv_std_logic_vector(37500, 16),
64151 => conv_std_logic_vector(37750, 16),
64152 => conv_std_logic_vector(38000, 16),
64153 => conv_std_logic_vector(38250, 16),
64154 => conv_std_logic_vector(38500, 16),
64155 => conv_std_logic_vector(38750, 16),
64156 => conv_std_logic_vector(39000, 16),
64157 => conv_std_logic_vector(39250, 16),
64158 => conv_std_logic_vector(39500, 16),
64159 => conv_std_logic_vector(39750, 16),
64160 => conv_std_logic_vector(40000, 16),
64161 => conv_std_logic_vector(40250, 16),
64162 => conv_std_logic_vector(40500, 16),
64163 => conv_std_logic_vector(40750, 16),
64164 => conv_std_logic_vector(41000, 16),
64165 => conv_std_logic_vector(41250, 16),
64166 => conv_std_logic_vector(41500, 16),
64167 => conv_std_logic_vector(41750, 16),
64168 => conv_std_logic_vector(42000, 16),
64169 => conv_std_logic_vector(42250, 16),
64170 => conv_std_logic_vector(42500, 16),
64171 => conv_std_logic_vector(42750, 16),
64172 => conv_std_logic_vector(43000, 16),
64173 => conv_std_logic_vector(43250, 16),
64174 => conv_std_logic_vector(43500, 16),
64175 => conv_std_logic_vector(43750, 16),
64176 => conv_std_logic_vector(44000, 16),
64177 => conv_std_logic_vector(44250, 16),
64178 => conv_std_logic_vector(44500, 16),
64179 => conv_std_logic_vector(44750, 16),
64180 => conv_std_logic_vector(45000, 16),
64181 => conv_std_logic_vector(45250, 16),
64182 => conv_std_logic_vector(45500, 16),
64183 => conv_std_logic_vector(45750, 16),
64184 => conv_std_logic_vector(46000, 16),
64185 => conv_std_logic_vector(46250, 16),
64186 => conv_std_logic_vector(46500, 16),
64187 => conv_std_logic_vector(46750, 16),
64188 => conv_std_logic_vector(47000, 16),
64189 => conv_std_logic_vector(47250, 16),
64190 => conv_std_logic_vector(47500, 16),
64191 => conv_std_logic_vector(47750, 16),
64192 => conv_std_logic_vector(48000, 16),
64193 => conv_std_logic_vector(48250, 16),
64194 => conv_std_logic_vector(48500, 16),
64195 => conv_std_logic_vector(48750, 16),
64196 => conv_std_logic_vector(49000, 16),
64197 => conv_std_logic_vector(49250, 16),
64198 => conv_std_logic_vector(49500, 16),
64199 => conv_std_logic_vector(49750, 16),
64200 => conv_std_logic_vector(50000, 16),
64201 => conv_std_logic_vector(50250, 16),
64202 => conv_std_logic_vector(50500, 16),
64203 => conv_std_logic_vector(50750, 16),
64204 => conv_std_logic_vector(51000, 16),
64205 => conv_std_logic_vector(51250, 16),
64206 => conv_std_logic_vector(51500, 16),
64207 => conv_std_logic_vector(51750, 16),
64208 => conv_std_logic_vector(52000, 16),
64209 => conv_std_logic_vector(52250, 16),
64210 => conv_std_logic_vector(52500, 16),
64211 => conv_std_logic_vector(52750, 16),
64212 => conv_std_logic_vector(53000, 16),
64213 => conv_std_logic_vector(53250, 16),
64214 => conv_std_logic_vector(53500, 16),
64215 => conv_std_logic_vector(53750, 16),
64216 => conv_std_logic_vector(54000, 16),
64217 => conv_std_logic_vector(54250, 16),
64218 => conv_std_logic_vector(54500, 16),
64219 => conv_std_logic_vector(54750, 16),
64220 => conv_std_logic_vector(55000, 16),
64221 => conv_std_logic_vector(55250, 16),
64222 => conv_std_logic_vector(55500, 16),
64223 => conv_std_logic_vector(55750, 16),
64224 => conv_std_logic_vector(56000, 16),
64225 => conv_std_logic_vector(56250, 16),
64226 => conv_std_logic_vector(56500, 16),
64227 => conv_std_logic_vector(56750, 16),
64228 => conv_std_logic_vector(57000, 16),
64229 => conv_std_logic_vector(57250, 16),
64230 => conv_std_logic_vector(57500, 16),
64231 => conv_std_logic_vector(57750, 16),
64232 => conv_std_logic_vector(58000, 16),
64233 => conv_std_logic_vector(58250, 16),
64234 => conv_std_logic_vector(58500, 16),
64235 => conv_std_logic_vector(58750, 16),
64236 => conv_std_logic_vector(59000, 16),
64237 => conv_std_logic_vector(59250, 16),
64238 => conv_std_logic_vector(59500, 16),
64239 => conv_std_logic_vector(59750, 16),
64240 => conv_std_logic_vector(60000, 16),
64241 => conv_std_logic_vector(60250, 16),
64242 => conv_std_logic_vector(60500, 16),
64243 => conv_std_logic_vector(60750, 16),
64244 => conv_std_logic_vector(61000, 16),
64245 => conv_std_logic_vector(61250, 16),
64246 => conv_std_logic_vector(61500, 16),
64247 => conv_std_logic_vector(61750, 16),
64248 => conv_std_logic_vector(62000, 16),
64249 => conv_std_logic_vector(62250, 16),
64250 => conv_std_logic_vector(62500, 16),
64251 => conv_std_logic_vector(62750, 16),
64252 => conv_std_logic_vector(63000, 16),
64253 => conv_std_logic_vector(63250, 16),
64254 => conv_std_logic_vector(63500, 16),
64255 => conv_std_logic_vector(63750, 16),
64256 => conv_std_logic_vector(0, 16),
64257 => conv_std_logic_vector(251, 16),
64258 => conv_std_logic_vector(502, 16),
64259 => conv_std_logic_vector(753, 16),
64260 => conv_std_logic_vector(1004, 16),
64261 => conv_std_logic_vector(1255, 16),
64262 => conv_std_logic_vector(1506, 16),
64263 => conv_std_logic_vector(1757, 16),
64264 => conv_std_logic_vector(2008, 16),
64265 => conv_std_logic_vector(2259, 16),
64266 => conv_std_logic_vector(2510, 16),
64267 => conv_std_logic_vector(2761, 16),
64268 => conv_std_logic_vector(3012, 16),
64269 => conv_std_logic_vector(3263, 16),
64270 => conv_std_logic_vector(3514, 16),
64271 => conv_std_logic_vector(3765, 16),
64272 => conv_std_logic_vector(4016, 16),
64273 => conv_std_logic_vector(4267, 16),
64274 => conv_std_logic_vector(4518, 16),
64275 => conv_std_logic_vector(4769, 16),
64276 => conv_std_logic_vector(5020, 16),
64277 => conv_std_logic_vector(5271, 16),
64278 => conv_std_logic_vector(5522, 16),
64279 => conv_std_logic_vector(5773, 16),
64280 => conv_std_logic_vector(6024, 16),
64281 => conv_std_logic_vector(6275, 16),
64282 => conv_std_logic_vector(6526, 16),
64283 => conv_std_logic_vector(6777, 16),
64284 => conv_std_logic_vector(7028, 16),
64285 => conv_std_logic_vector(7279, 16),
64286 => conv_std_logic_vector(7530, 16),
64287 => conv_std_logic_vector(7781, 16),
64288 => conv_std_logic_vector(8032, 16),
64289 => conv_std_logic_vector(8283, 16),
64290 => conv_std_logic_vector(8534, 16),
64291 => conv_std_logic_vector(8785, 16),
64292 => conv_std_logic_vector(9036, 16),
64293 => conv_std_logic_vector(9287, 16),
64294 => conv_std_logic_vector(9538, 16),
64295 => conv_std_logic_vector(9789, 16),
64296 => conv_std_logic_vector(10040, 16),
64297 => conv_std_logic_vector(10291, 16),
64298 => conv_std_logic_vector(10542, 16),
64299 => conv_std_logic_vector(10793, 16),
64300 => conv_std_logic_vector(11044, 16),
64301 => conv_std_logic_vector(11295, 16),
64302 => conv_std_logic_vector(11546, 16),
64303 => conv_std_logic_vector(11797, 16),
64304 => conv_std_logic_vector(12048, 16),
64305 => conv_std_logic_vector(12299, 16),
64306 => conv_std_logic_vector(12550, 16),
64307 => conv_std_logic_vector(12801, 16),
64308 => conv_std_logic_vector(13052, 16),
64309 => conv_std_logic_vector(13303, 16),
64310 => conv_std_logic_vector(13554, 16),
64311 => conv_std_logic_vector(13805, 16),
64312 => conv_std_logic_vector(14056, 16),
64313 => conv_std_logic_vector(14307, 16),
64314 => conv_std_logic_vector(14558, 16),
64315 => conv_std_logic_vector(14809, 16),
64316 => conv_std_logic_vector(15060, 16),
64317 => conv_std_logic_vector(15311, 16),
64318 => conv_std_logic_vector(15562, 16),
64319 => conv_std_logic_vector(15813, 16),
64320 => conv_std_logic_vector(16064, 16),
64321 => conv_std_logic_vector(16315, 16),
64322 => conv_std_logic_vector(16566, 16),
64323 => conv_std_logic_vector(16817, 16),
64324 => conv_std_logic_vector(17068, 16),
64325 => conv_std_logic_vector(17319, 16),
64326 => conv_std_logic_vector(17570, 16),
64327 => conv_std_logic_vector(17821, 16),
64328 => conv_std_logic_vector(18072, 16),
64329 => conv_std_logic_vector(18323, 16),
64330 => conv_std_logic_vector(18574, 16),
64331 => conv_std_logic_vector(18825, 16),
64332 => conv_std_logic_vector(19076, 16),
64333 => conv_std_logic_vector(19327, 16),
64334 => conv_std_logic_vector(19578, 16),
64335 => conv_std_logic_vector(19829, 16),
64336 => conv_std_logic_vector(20080, 16),
64337 => conv_std_logic_vector(20331, 16),
64338 => conv_std_logic_vector(20582, 16),
64339 => conv_std_logic_vector(20833, 16),
64340 => conv_std_logic_vector(21084, 16),
64341 => conv_std_logic_vector(21335, 16),
64342 => conv_std_logic_vector(21586, 16),
64343 => conv_std_logic_vector(21837, 16),
64344 => conv_std_logic_vector(22088, 16),
64345 => conv_std_logic_vector(22339, 16),
64346 => conv_std_logic_vector(22590, 16),
64347 => conv_std_logic_vector(22841, 16),
64348 => conv_std_logic_vector(23092, 16),
64349 => conv_std_logic_vector(23343, 16),
64350 => conv_std_logic_vector(23594, 16),
64351 => conv_std_logic_vector(23845, 16),
64352 => conv_std_logic_vector(24096, 16),
64353 => conv_std_logic_vector(24347, 16),
64354 => conv_std_logic_vector(24598, 16),
64355 => conv_std_logic_vector(24849, 16),
64356 => conv_std_logic_vector(25100, 16),
64357 => conv_std_logic_vector(25351, 16),
64358 => conv_std_logic_vector(25602, 16),
64359 => conv_std_logic_vector(25853, 16),
64360 => conv_std_logic_vector(26104, 16),
64361 => conv_std_logic_vector(26355, 16),
64362 => conv_std_logic_vector(26606, 16),
64363 => conv_std_logic_vector(26857, 16),
64364 => conv_std_logic_vector(27108, 16),
64365 => conv_std_logic_vector(27359, 16),
64366 => conv_std_logic_vector(27610, 16),
64367 => conv_std_logic_vector(27861, 16),
64368 => conv_std_logic_vector(28112, 16),
64369 => conv_std_logic_vector(28363, 16),
64370 => conv_std_logic_vector(28614, 16),
64371 => conv_std_logic_vector(28865, 16),
64372 => conv_std_logic_vector(29116, 16),
64373 => conv_std_logic_vector(29367, 16),
64374 => conv_std_logic_vector(29618, 16),
64375 => conv_std_logic_vector(29869, 16),
64376 => conv_std_logic_vector(30120, 16),
64377 => conv_std_logic_vector(30371, 16),
64378 => conv_std_logic_vector(30622, 16),
64379 => conv_std_logic_vector(30873, 16),
64380 => conv_std_logic_vector(31124, 16),
64381 => conv_std_logic_vector(31375, 16),
64382 => conv_std_logic_vector(31626, 16),
64383 => conv_std_logic_vector(31877, 16),
64384 => conv_std_logic_vector(32128, 16),
64385 => conv_std_logic_vector(32379, 16),
64386 => conv_std_logic_vector(32630, 16),
64387 => conv_std_logic_vector(32881, 16),
64388 => conv_std_logic_vector(33132, 16),
64389 => conv_std_logic_vector(33383, 16),
64390 => conv_std_logic_vector(33634, 16),
64391 => conv_std_logic_vector(33885, 16),
64392 => conv_std_logic_vector(34136, 16),
64393 => conv_std_logic_vector(34387, 16),
64394 => conv_std_logic_vector(34638, 16),
64395 => conv_std_logic_vector(34889, 16),
64396 => conv_std_logic_vector(35140, 16),
64397 => conv_std_logic_vector(35391, 16),
64398 => conv_std_logic_vector(35642, 16),
64399 => conv_std_logic_vector(35893, 16),
64400 => conv_std_logic_vector(36144, 16),
64401 => conv_std_logic_vector(36395, 16),
64402 => conv_std_logic_vector(36646, 16),
64403 => conv_std_logic_vector(36897, 16),
64404 => conv_std_logic_vector(37148, 16),
64405 => conv_std_logic_vector(37399, 16),
64406 => conv_std_logic_vector(37650, 16),
64407 => conv_std_logic_vector(37901, 16),
64408 => conv_std_logic_vector(38152, 16),
64409 => conv_std_logic_vector(38403, 16),
64410 => conv_std_logic_vector(38654, 16),
64411 => conv_std_logic_vector(38905, 16),
64412 => conv_std_logic_vector(39156, 16),
64413 => conv_std_logic_vector(39407, 16),
64414 => conv_std_logic_vector(39658, 16),
64415 => conv_std_logic_vector(39909, 16),
64416 => conv_std_logic_vector(40160, 16),
64417 => conv_std_logic_vector(40411, 16),
64418 => conv_std_logic_vector(40662, 16),
64419 => conv_std_logic_vector(40913, 16),
64420 => conv_std_logic_vector(41164, 16),
64421 => conv_std_logic_vector(41415, 16),
64422 => conv_std_logic_vector(41666, 16),
64423 => conv_std_logic_vector(41917, 16),
64424 => conv_std_logic_vector(42168, 16),
64425 => conv_std_logic_vector(42419, 16),
64426 => conv_std_logic_vector(42670, 16),
64427 => conv_std_logic_vector(42921, 16),
64428 => conv_std_logic_vector(43172, 16),
64429 => conv_std_logic_vector(43423, 16),
64430 => conv_std_logic_vector(43674, 16),
64431 => conv_std_logic_vector(43925, 16),
64432 => conv_std_logic_vector(44176, 16),
64433 => conv_std_logic_vector(44427, 16),
64434 => conv_std_logic_vector(44678, 16),
64435 => conv_std_logic_vector(44929, 16),
64436 => conv_std_logic_vector(45180, 16),
64437 => conv_std_logic_vector(45431, 16),
64438 => conv_std_logic_vector(45682, 16),
64439 => conv_std_logic_vector(45933, 16),
64440 => conv_std_logic_vector(46184, 16),
64441 => conv_std_logic_vector(46435, 16),
64442 => conv_std_logic_vector(46686, 16),
64443 => conv_std_logic_vector(46937, 16),
64444 => conv_std_logic_vector(47188, 16),
64445 => conv_std_logic_vector(47439, 16),
64446 => conv_std_logic_vector(47690, 16),
64447 => conv_std_logic_vector(47941, 16),
64448 => conv_std_logic_vector(48192, 16),
64449 => conv_std_logic_vector(48443, 16),
64450 => conv_std_logic_vector(48694, 16),
64451 => conv_std_logic_vector(48945, 16),
64452 => conv_std_logic_vector(49196, 16),
64453 => conv_std_logic_vector(49447, 16),
64454 => conv_std_logic_vector(49698, 16),
64455 => conv_std_logic_vector(49949, 16),
64456 => conv_std_logic_vector(50200, 16),
64457 => conv_std_logic_vector(50451, 16),
64458 => conv_std_logic_vector(50702, 16),
64459 => conv_std_logic_vector(50953, 16),
64460 => conv_std_logic_vector(51204, 16),
64461 => conv_std_logic_vector(51455, 16),
64462 => conv_std_logic_vector(51706, 16),
64463 => conv_std_logic_vector(51957, 16),
64464 => conv_std_logic_vector(52208, 16),
64465 => conv_std_logic_vector(52459, 16),
64466 => conv_std_logic_vector(52710, 16),
64467 => conv_std_logic_vector(52961, 16),
64468 => conv_std_logic_vector(53212, 16),
64469 => conv_std_logic_vector(53463, 16),
64470 => conv_std_logic_vector(53714, 16),
64471 => conv_std_logic_vector(53965, 16),
64472 => conv_std_logic_vector(54216, 16),
64473 => conv_std_logic_vector(54467, 16),
64474 => conv_std_logic_vector(54718, 16),
64475 => conv_std_logic_vector(54969, 16),
64476 => conv_std_logic_vector(55220, 16),
64477 => conv_std_logic_vector(55471, 16),
64478 => conv_std_logic_vector(55722, 16),
64479 => conv_std_logic_vector(55973, 16),
64480 => conv_std_logic_vector(56224, 16),
64481 => conv_std_logic_vector(56475, 16),
64482 => conv_std_logic_vector(56726, 16),
64483 => conv_std_logic_vector(56977, 16),
64484 => conv_std_logic_vector(57228, 16),
64485 => conv_std_logic_vector(57479, 16),
64486 => conv_std_logic_vector(57730, 16),
64487 => conv_std_logic_vector(57981, 16),
64488 => conv_std_logic_vector(58232, 16),
64489 => conv_std_logic_vector(58483, 16),
64490 => conv_std_logic_vector(58734, 16),
64491 => conv_std_logic_vector(58985, 16),
64492 => conv_std_logic_vector(59236, 16),
64493 => conv_std_logic_vector(59487, 16),
64494 => conv_std_logic_vector(59738, 16),
64495 => conv_std_logic_vector(59989, 16),
64496 => conv_std_logic_vector(60240, 16),
64497 => conv_std_logic_vector(60491, 16),
64498 => conv_std_logic_vector(60742, 16),
64499 => conv_std_logic_vector(60993, 16),
64500 => conv_std_logic_vector(61244, 16),
64501 => conv_std_logic_vector(61495, 16),
64502 => conv_std_logic_vector(61746, 16),
64503 => conv_std_logic_vector(61997, 16),
64504 => conv_std_logic_vector(62248, 16),
64505 => conv_std_logic_vector(62499, 16),
64506 => conv_std_logic_vector(62750, 16),
64507 => conv_std_logic_vector(63001, 16),
64508 => conv_std_logic_vector(63252, 16),
64509 => conv_std_logic_vector(63503, 16),
64510 => conv_std_logic_vector(63754, 16),
64511 => conv_std_logic_vector(64005, 16),
64512 => conv_std_logic_vector(0, 16),
64513 => conv_std_logic_vector(252, 16),
64514 => conv_std_logic_vector(504, 16),
64515 => conv_std_logic_vector(756, 16),
64516 => conv_std_logic_vector(1008, 16),
64517 => conv_std_logic_vector(1260, 16),
64518 => conv_std_logic_vector(1512, 16),
64519 => conv_std_logic_vector(1764, 16),
64520 => conv_std_logic_vector(2016, 16),
64521 => conv_std_logic_vector(2268, 16),
64522 => conv_std_logic_vector(2520, 16),
64523 => conv_std_logic_vector(2772, 16),
64524 => conv_std_logic_vector(3024, 16),
64525 => conv_std_logic_vector(3276, 16),
64526 => conv_std_logic_vector(3528, 16),
64527 => conv_std_logic_vector(3780, 16),
64528 => conv_std_logic_vector(4032, 16),
64529 => conv_std_logic_vector(4284, 16),
64530 => conv_std_logic_vector(4536, 16),
64531 => conv_std_logic_vector(4788, 16),
64532 => conv_std_logic_vector(5040, 16),
64533 => conv_std_logic_vector(5292, 16),
64534 => conv_std_logic_vector(5544, 16),
64535 => conv_std_logic_vector(5796, 16),
64536 => conv_std_logic_vector(6048, 16),
64537 => conv_std_logic_vector(6300, 16),
64538 => conv_std_logic_vector(6552, 16),
64539 => conv_std_logic_vector(6804, 16),
64540 => conv_std_logic_vector(7056, 16),
64541 => conv_std_logic_vector(7308, 16),
64542 => conv_std_logic_vector(7560, 16),
64543 => conv_std_logic_vector(7812, 16),
64544 => conv_std_logic_vector(8064, 16),
64545 => conv_std_logic_vector(8316, 16),
64546 => conv_std_logic_vector(8568, 16),
64547 => conv_std_logic_vector(8820, 16),
64548 => conv_std_logic_vector(9072, 16),
64549 => conv_std_logic_vector(9324, 16),
64550 => conv_std_logic_vector(9576, 16),
64551 => conv_std_logic_vector(9828, 16),
64552 => conv_std_logic_vector(10080, 16),
64553 => conv_std_logic_vector(10332, 16),
64554 => conv_std_logic_vector(10584, 16),
64555 => conv_std_logic_vector(10836, 16),
64556 => conv_std_logic_vector(11088, 16),
64557 => conv_std_logic_vector(11340, 16),
64558 => conv_std_logic_vector(11592, 16),
64559 => conv_std_logic_vector(11844, 16),
64560 => conv_std_logic_vector(12096, 16),
64561 => conv_std_logic_vector(12348, 16),
64562 => conv_std_logic_vector(12600, 16),
64563 => conv_std_logic_vector(12852, 16),
64564 => conv_std_logic_vector(13104, 16),
64565 => conv_std_logic_vector(13356, 16),
64566 => conv_std_logic_vector(13608, 16),
64567 => conv_std_logic_vector(13860, 16),
64568 => conv_std_logic_vector(14112, 16),
64569 => conv_std_logic_vector(14364, 16),
64570 => conv_std_logic_vector(14616, 16),
64571 => conv_std_logic_vector(14868, 16),
64572 => conv_std_logic_vector(15120, 16),
64573 => conv_std_logic_vector(15372, 16),
64574 => conv_std_logic_vector(15624, 16),
64575 => conv_std_logic_vector(15876, 16),
64576 => conv_std_logic_vector(16128, 16),
64577 => conv_std_logic_vector(16380, 16),
64578 => conv_std_logic_vector(16632, 16),
64579 => conv_std_logic_vector(16884, 16),
64580 => conv_std_logic_vector(17136, 16),
64581 => conv_std_logic_vector(17388, 16),
64582 => conv_std_logic_vector(17640, 16),
64583 => conv_std_logic_vector(17892, 16),
64584 => conv_std_logic_vector(18144, 16),
64585 => conv_std_logic_vector(18396, 16),
64586 => conv_std_logic_vector(18648, 16),
64587 => conv_std_logic_vector(18900, 16),
64588 => conv_std_logic_vector(19152, 16),
64589 => conv_std_logic_vector(19404, 16),
64590 => conv_std_logic_vector(19656, 16),
64591 => conv_std_logic_vector(19908, 16),
64592 => conv_std_logic_vector(20160, 16),
64593 => conv_std_logic_vector(20412, 16),
64594 => conv_std_logic_vector(20664, 16),
64595 => conv_std_logic_vector(20916, 16),
64596 => conv_std_logic_vector(21168, 16),
64597 => conv_std_logic_vector(21420, 16),
64598 => conv_std_logic_vector(21672, 16),
64599 => conv_std_logic_vector(21924, 16),
64600 => conv_std_logic_vector(22176, 16),
64601 => conv_std_logic_vector(22428, 16),
64602 => conv_std_logic_vector(22680, 16),
64603 => conv_std_logic_vector(22932, 16),
64604 => conv_std_logic_vector(23184, 16),
64605 => conv_std_logic_vector(23436, 16),
64606 => conv_std_logic_vector(23688, 16),
64607 => conv_std_logic_vector(23940, 16),
64608 => conv_std_logic_vector(24192, 16),
64609 => conv_std_logic_vector(24444, 16),
64610 => conv_std_logic_vector(24696, 16),
64611 => conv_std_logic_vector(24948, 16),
64612 => conv_std_logic_vector(25200, 16),
64613 => conv_std_logic_vector(25452, 16),
64614 => conv_std_logic_vector(25704, 16),
64615 => conv_std_logic_vector(25956, 16),
64616 => conv_std_logic_vector(26208, 16),
64617 => conv_std_logic_vector(26460, 16),
64618 => conv_std_logic_vector(26712, 16),
64619 => conv_std_logic_vector(26964, 16),
64620 => conv_std_logic_vector(27216, 16),
64621 => conv_std_logic_vector(27468, 16),
64622 => conv_std_logic_vector(27720, 16),
64623 => conv_std_logic_vector(27972, 16),
64624 => conv_std_logic_vector(28224, 16),
64625 => conv_std_logic_vector(28476, 16),
64626 => conv_std_logic_vector(28728, 16),
64627 => conv_std_logic_vector(28980, 16),
64628 => conv_std_logic_vector(29232, 16),
64629 => conv_std_logic_vector(29484, 16),
64630 => conv_std_logic_vector(29736, 16),
64631 => conv_std_logic_vector(29988, 16),
64632 => conv_std_logic_vector(30240, 16),
64633 => conv_std_logic_vector(30492, 16),
64634 => conv_std_logic_vector(30744, 16),
64635 => conv_std_logic_vector(30996, 16),
64636 => conv_std_logic_vector(31248, 16),
64637 => conv_std_logic_vector(31500, 16),
64638 => conv_std_logic_vector(31752, 16),
64639 => conv_std_logic_vector(32004, 16),
64640 => conv_std_logic_vector(32256, 16),
64641 => conv_std_logic_vector(32508, 16),
64642 => conv_std_logic_vector(32760, 16),
64643 => conv_std_logic_vector(33012, 16),
64644 => conv_std_logic_vector(33264, 16),
64645 => conv_std_logic_vector(33516, 16),
64646 => conv_std_logic_vector(33768, 16),
64647 => conv_std_logic_vector(34020, 16),
64648 => conv_std_logic_vector(34272, 16),
64649 => conv_std_logic_vector(34524, 16),
64650 => conv_std_logic_vector(34776, 16),
64651 => conv_std_logic_vector(35028, 16),
64652 => conv_std_logic_vector(35280, 16),
64653 => conv_std_logic_vector(35532, 16),
64654 => conv_std_logic_vector(35784, 16),
64655 => conv_std_logic_vector(36036, 16),
64656 => conv_std_logic_vector(36288, 16),
64657 => conv_std_logic_vector(36540, 16),
64658 => conv_std_logic_vector(36792, 16),
64659 => conv_std_logic_vector(37044, 16),
64660 => conv_std_logic_vector(37296, 16),
64661 => conv_std_logic_vector(37548, 16),
64662 => conv_std_logic_vector(37800, 16),
64663 => conv_std_logic_vector(38052, 16),
64664 => conv_std_logic_vector(38304, 16),
64665 => conv_std_logic_vector(38556, 16),
64666 => conv_std_logic_vector(38808, 16),
64667 => conv_std_logic_vector(39060, 16),
64668 => conv_std_logic_vector(39312, 16),
64669 => conv_std_logic_vector(39564, 16),
64670 => conv_std_logic_vector(39816, 16),
64671 => conv_std_logic_vector(40068, 16),
64672 => conv_std_logic_vector(40320, 16),
64673 => conv_std_logic_vector(40572, 16),
64674 => conv_std_logic_vector(40824, 16),
64675 => conv_std_logic_vector(41076, 16),
64676 => conv_std_logic_vector(41328, 16),
64677 => conv_std_logic_vector(41580, 16),
64678 => conv_std_logic_vector(41832, 16),
64679 => conv_std_logic_vector(42084, 16),
64680 => conv_std_logic_vector(42336, 16),
64681 => conv_std_logic_vector(42588, 16),
64682 => conv_std_logic_vector(42840, 16),
64683 => conv_std_logic_vector(43092, 16),
64684 => conv_std_logic_vector(43344, 16),
64685 => conv_std_logic_vector(43596, 16),
64686 => conv_std_logic_vector(43848, 16),
64687 => conv_std_logic_vector(44100, 16),
64688 => conv_std_logic_vector(44352, 16),
64689 => conv_std_logic_vector(44604, 16),
64690 => conv_std_logic_vector(44856, 16),
64691 => conv_std_logic_vector(45108, 16),
64692 => conv_std_logic_vector(45360, 16),
64693 => conv_std_logic_vector(45612, 16),
64694 => conv_std_logic_vector(45864, 16),
64695 => conv_std_logic_vector(46116, 16),
64696 => conv_std_logic_vector(46368, 16),
64697 => conv_std_logic_vector(46620, 16),
64698 => conv_std_logic_vector(46872, 16),
64699 => conv_std_logic_vector(47124, 16),
64700 => conv_std_logic_vector(47376, 16),
64701 => conv_std_logic_vector(47628, 16),
64702 => conv_std_logic_vector(47880, 16),
64703 => conv_std_logic_vector(48132, 16),
64704 => conv_std_logic_vector(48384, 16),
64705 => conv_std_logic_vector(48636, 16),
64706 => conv_std_logic_vector(48888, 16),
64707 => conv_std_logic_vector(49140, 16),
64708 => conv_std_logic_vector(49392, 16),
64709 => conv_std_logic_vector(49644, 16),
64710 => conv_std_logic_vector(49896, 16),
64711 => conv_std_logic_vector(50148, 16),
64712 => conv_std_logic_vector(50400, 16),
64713 => conv_std_logic_vector(50652, 16),
64714 => conv_std_logic_vector(50904, 16),
64715 => conv_std_logic_vector(51156, 16),
64716 => conv_std_logic_vector(51408, 16),
64717 => conv_std_logic_vector(51660, 16),
64718 => conv_std_logic_vector(51912, 16),
64719 => conv_std_logic_vector(52164, 16),
64720 => conv_std_logic_vector(52416, 16),
64721 => conv_std_logic_vector(52668, 16),
64722 => conv_std_logic_vector(52920, 16),
64723 => conv_std_logic_vector(53172, 16),
64724 => conv_std_logic_vector(53424, 16),
64725 => conv_std_logic_vector(53676, 16),
64726 => conv_std_logic_vector(53928, 16),
64727 => conv_std_logic_vector(54180, 16),
64728 => conv_std_logic_vector(54432, 16),
64729 => conv_std_logic_vector(54684, 16),
64730 => conv_std_logic_vector(54936, 16),
64731 => conv_std_logic_vector(55188, 16),
64732 => conv_std_logic_vector(55440, 16),
64733 => conv_std_logic_vector(55692, 16),
64734 => conv_std_logic_vector(55944, 16),
64735 => conv_std_logic_vector(56196, 16),
64736 => conv_std_logic_vector(56448, 16),
64737 => conv_std_logic_vector(56700, 16),
64738 => conv_std_logic_vector(56952, 16),
64739 => conv_std_logic_vector(57204, 16),
64740 => conv_std_logic_vector(57456, 16),
64741 => conv_std_logic_vector(57708, 16),
64742 => conv_std_logic_vector(57960, 16),
64743 => conv_std_logic_vector(58212, 16),
64744 => conv_std_logic_vector(58464, 16),
64745 => conv_std_logic_vector(58716, 16),
64746 => conv_std_logic_vector(58968, 16),
64747 => conv_std_logic_vector(59220, 16),
64748 => conv_std_logic_vector(59472, 16),
64749 => conv_std_logic_vector(59724, 16),
64750 => conv_std_logic_vector(59976, 16),
64751 => conv_std_logic_vector(60228, 16),
64752 => conv_std_logic_vector(60480, 16),
64753 => conv_std_logic_vector(60732, 16),
64754 => conv_std_logic_vector(60984, 16),
64755 => conv_std_logic_vector(61236, 16),
64756 => conv_std_logic_vector(61488, 16),
64757 => conv_std_logic_vector(61740, 16),
64758 => conv_std_logic_vector(61992, 16),
64759 => conv_std_logic_vector(62244, 16),
64760 => conv_std_logic_vector(62496, 16),
64761 => conv_std_logic_vector(62748, 16),
64762 => conv_std_logic_vector(63000, 16),
64763 => conv_std_logic_vector(63252, 16),
64764 => conv_std_logic_vector(63504, 16),
64765 => conv_std_logic_vector(63756, 16),
64766 => conv_std_logic_vector(64008, 16),
64767 => conv_std_logic_vector(64260, 16),
64768 => conv_std_logic_vector(0, 16),
64769 => conv_std_logic_vector(253, 16),
64770 => conv_std_logic_vector(506, 16),
64771 => conv_std_logic_vector(759, 16),
64772 => conv_std_logic_vector(1012, 16),
64773 => conv_std_logic_vector(1265, 16),
64774 => conv_std_logic_vector(1518, 16),
64775 => conv_std_logic_vector(1771, 16),
64776 => conv_std_logic_vector(2024, 16),
64777 => conv_std_logic_vector(2277, 16),
64778 => conv_std_logic_vector(2530, 16),
64779 => conv_std_logic_vector(2783, 16),
64780 => conv_std_logic_vector(3036, 16),
64781 => conv_std_logic_vector(3289, 16),
64782 => conv_std_logic_vector(3542, 16),
64783 => conv_std_logic_vector(3795, 16),
64784 => conv_std_logic_vector(4048, 16),
64785 => conv_std_logic_vector(4301, 16),
64786 => conv_std_logic_vector(4554, 16),
64787 => conv_std_logic_vector(4807, 16),
64788 => conv_std_logic_vector(5060, 16),
64789 => conv_std_logic_vector(5313, 16),
64790 => conv_std_logic_vector(5566, 16),
64791 => conv_std_logic_vector(5819, 16),
64792 => conv_std_logic_vector(6072, 16),
64793 => conv_std_logic_vector(6325, 16),
64794 => conv_std_logic_vector(6578, 16),
64795 => conv_std_logic_vector(6831, 16),
64796 => conv_std_logic_vector(7084, 16),
64797 => conv_std_logic_vector(7337, 16),
64798 => conv_std_logic_vector(7590, 16),
64799 => conv_std_logic_vector(7843, 16),
64800 => conv_std_logic_vector(8096, 16),
64801 => conv_std_logic_vector(8349, 16),
64802 => conv_std_logic_vector(8602, 16),
64803 => conv_std_logic_vector(8855, 16),
64804 => conv_std_logic_vector(9108, 16),
64805 => conv_std_logic_vector(9361, 16),
64806 => conv_std_logic_vector(9614, 16),
64807 => conv_std_logic_vector(9867, 16),
64808 => conv_std_logic_vector(10120, 16),
64809 => conv_std_logic_vector(10373, 16),
64810 => conv_std_logic_vector(10626, 16),
64811 => conv_std_logic_vector(10879, 16),
64812 => conv_std_logic_vector(11132, 16),
64813 => conv_std_logic_vector(11385, 16),
64814 => conv_std_logic_vector(11638, 16),
64815 => conv_std_logic_vector(11891, 16),
64816 => conv_std_logic_vector(12144, 16),
64817 => conv_std_logic_vector(12397, 16),
64818 => conv_std_logic_vector(12650, 16),
64819 => conv_std_logic_vector(12903, 16),
64820 => conv_std_logic_vector(13156, 16),
64821 => conv_std_logic_vector(13409, 16),
64822 => conv_std_logic_vector(13662, 16),
64823 => conv_std_logic_vector(13915, 16),
64824 => conv_std_logic_vector(14168, 16),
64825 => conv_std_logic_vector(14421, 16),
64826 => conv_std_logic_vector(14674, 16),
64827 => conv_std_logic_vector(14927, 16),
64828 => conv_std_logic_vector(15180, 16),
64829 => conv_std_logic_vector(15433, 16),
64830 => conv_std_logic_vector(15686, 16),
64831 => conv_std_logic_vector(15939, 16),
64832 => conv_std_logic_vector(16192, 16),
64833 => conv_std_logic_vector(16445, 16),
64834 => conv_std_logic_vector(16698, 16),
64835 => conv_std_logic_vector(16951, 16),
64836 => conv_std_logic_vector(17204, 16),
64837 => conv_std_logic_vector(17457, 16),
64838 => conv_std_logic_vector(17710, 16),
64839 => conv_std_logic_vector(17963, 16),
64840 => conv_std_logic_vector(18216, 16),
64841 => conv_std_logic_vector(18469, 16),
64842 => conv_std_logic_vector(18722, 16),
64843 => conv_std_logic_vector(18975, 16),
64844 => conv_std_logic_vector(19228, 16),
64845 => conv_std_logic_vector(19481, 16),
64846 => conv_std_logic_vector(19734, 16),
64847 => conv_std_logic_vector(19987, 16),
64848 => conv_std_logic_vector(20240, 16),
64849 => conv_std_logic_vector(20493, 16),
64850 => conv_std_logic_vector(20746, 16),
64851 => conv_std_logic_vector(20999, 16),
64852 => conv_std_logic_vector(21252, 16),
64853 => conv_std_logic_vector(21505, 16),
64854 => conv_std_logic_vector(21758, 16),
64855 => conv_std_logic_vector(22011, 16),
64856 => conv_std_logic_vector(22264, 16),
64857 => conv_std_logic_vector(22517, 16),
64858 => conv_std_logic_vector(22770, 16),
64859 => conv_std_logic_vector(23023, 16),
64860 => conv_std_logic_vector(23276, 16),
64861 => conv_std_logic_vector(23529, 16),
64862 => conv_std_logic_vector(23782, 16),
64863 => conv_std_logic_vector(24035, 16),
64864 => conv_std_logic_vector(24288, 16),
64865 => conv_std_logic_vector(24541, 16),
64866 => conv_std_logic_vector(24794, 16),
64867 => conv_std_logic_vector(25047, 16),
64868 => conv_std_logic_vector(25300, 16),
64869 => conv_std_logic_vector(25553, 16),
64870 => conv_std_logic_vector(25806, 16),
64871 => conv_std_logic_vector(26059, 16),
64872 => conv_std_logic_vector(26312, 16),
64873 => conv_std_logic_vector(26565, 16),
64874 => conv_std_logic_vector(26818, 16),
64875 => conv_std_logic_vector(27071, 16),
64876 => conv_std_logic_vector(27324, 16),
64877 => conv_std_logic_vector(27577, 16),
64878 => conv_std_logic_vector(27830, 16),
64879 => conv_std_logic_vector(28083, 16),
64880 => conv_std_logic_vector(28336, 16),
64881 => conv_std_logic_vector(28589, 16),
64882 => conv_std_logic_vector(28842, 16),
64883 => conv_std_logic_vector(29095, 16),
64884 => conv_std_logic_vector(29348, 16),
64885 => conv_std_logic_vector(29601, 16),
64886 => conv_std_logic_vector(29854, 16),
64887 => conv_std_logic_vector(30107, 16),
64888 => conv_std_logic_vector(30360, 16),
64889 => conv_std_logic_vector(30613, 16),
64890 => conv_std_logic_vector(30866, 16),
64891 => conv_std_logic_vector(31119, 16),
64892 => conv_std_logic_vector(31372, 16),
64893 => conv_std_logic_vector(31625, 16),
64894 => conv_std_logic_vector(31878, 16),
64895 => conv_std_logic_vector(32131, 16),
64896 => conv_std_logic_vector(32384, 16),
64897 => conv_std_logic_vector(32637, 16),
64898 => conv_std_logic_vector(32890, 16),
64899 => conv_std_logic_vector(33143, 16),
64900 => conv_std_logic_vector(33396, 16),
64901 => conv_std_logic_vector(33649, 16),
64902 => conv_std_logic_vector(33902, 16),
64903 => conv_std_logic_vector(34155, 16),
64904 => conv_std_logic_vector(34408, 16),
64905 => conv_std_logic_vector(34661, 16),
64906 => conv_std_logic_vector(34914, 16),
64907 => conv_std_logic_vector(35167, 16),
64908 => conv_std_logic_vector(35420, 16),
64909 => conv_std_logic_vector(35673, 16),
64910 => conv_std_logic_vector(35926, 16),
64911 => conv_std_logic_vector(36179, 16),
64912 => conv_std_logic_vector(36432, 16),
64913 => conv_std_logic_vector(36685, 16),
64914 => conv_std_logic_vector(36938, 16),
64915 => conv_std_logic_vector(37191, 16),
64916 => conv_std_logic_vector(37444, 16),
64917 => conv_std_logic_vector(37697, 16),
64918 => conv_std_logic_vector(37950, 16),
64919 => conv_std_logic_vector(38203, 16),
64920 => conv_std_logic_vector(38456, 16),
64921 => conv_std_logic_vector(38709, 16),
64922 => conv_std_logic_vector(38962, 16),
64923 => conv_std_logic_vector(39215, 16),
64924 => conv_std_logic_vector(39468, 16),
64925 => conv_std_logic_vector(39721, 16),
64926 => conv_std_logic_vector(39974, 16),
64927 => conv_std_logic_vector(40227, 16),
64928 => conv_std_logic_vector(40480, 16),
64929 => conv_std_logic_vector(40733, 16),
64930 => conv_std_logic_vector(40986, 16),
64931 => conv_std_logic_vector(41239, 16),
64932 => conv_std_logic_vector(41492, 16),
64933 => conv_std_logic_vector(41745, 16),
64934 => conv_std_logic_vector(41998, 16),
64935 => conv_std_logic_vector(42251, 16),
64936 => conv_std_logic_vector(42504, 16),
64937 => conv_std_logic_vector(42757, 16),
64938 => conv_std_logic_vector(43010, 16),
64939 => conv_std_logic_vector(43263, 16),
64940 => conv_std_logic_vector(43516, 16),
64941 => conv_std_logic_vector(43769, 16),
64942 => conv_std_logic_vector(44022, 16),
64943 => conv_std_logic_vector(44275, 16),
64944 => conv_std_logic_vector(44528, 16),
64945 => conv_std_logic_vector(44781, 16),
64946 => conv_std_logic_vector(45034, 16),
64947 => conv_std_logic_vector(45287, 16),
64948 => conv_std_logic_vector(45540, 16),
64949 => conv_std_logic_vector(45793, 16),
64950 => conv_std_logic_vector(46046, 16),
64951 => conv_std_logic_vector(46299, 16),
64952 => conv_std_logic_vector(46552, 16),
64953 => conv_std_logic_vector(46805, 16),
64954 => conv_std_logic_vector(47058, 16),
64955 => conv_std_logic_vector(47311, 16),
64956 => conv_std_logic_vector(47564, 16),
64957 => conv_std_logic_vector(47817, 16),
64958 => conv_std_logic_vector(48070, 16),
64959 => conv_std_logic_vector(48323, 16),
64960 => conv_std_logic_vector(48576, 16),
64961 => conv_std_logic_vector(48829, 16),
64962 => conv_std_logic_vector(49082, 16),
64963 => conv_std_logic_vector(49335, 16),
64964 => conv_std_logic_vector(49588, 16),
64965 => conv_std_logic_vector(49841, 16),
64966 => conv_std_logic_vector(50094, 16),
64967 => conv_std_logic_vector(50347, 16),
64968 => conv_std_logic_vector(50600, 16),
64969 => conv_std_logic_vector(50853, 16),
64970 => conv_std_logic_vector(51106, 16),
64971 => conv_std_logic_vector(51359, 16),
64972 => conv_std_logic_vector(51612, 16),
64973 => conv_std_logic_vector(51865, 16),
64974 => conv_std_logic_vector(52118, 16),
64975 => conv_std_logic_vector(52371, 16),
64976 => conv_std_logic_vector(52624, 16),
64977 => conv_std_logic_vector(52877, 16),
64978 => conv_std_logic_vector(53130, 16),
64979 => conv_std_logic_vector(53383, 16),
64980 => conv_std_logic_vector(53636, 16),
64981 => conv_std_logic_vector(53889, 16),
64982 => conv_std_logic_vector(54142, 16),
64983 => conv_std_logic_vector(54395, 16),
64984 => conv_std_logic_vector(54648, 16),
64985 => conv_std_logic_vector(54901, 16),
64986 => conv_std_logic_vector(55154, 16),
64987 => conv_std_logic_vector(55407, 16),
64988 => conv_std_logic_vector(55660, 16),
64989 => conv_std_logic_vector(55913, 16),
64990 => conv_std_logic_vector(56166, 16),
64991 => conv_std_logic_vector(56419, 16),
64992 => conv_std_logic_vector(56672, 16),
64993 => conv_std_logic_vector(56925, 16),
64994 => conv_std_logic_vector(57178, 16),
64995 => conv_std_logic_vector(57431, 16),
64996 => conv_std_logic_vector(57684, 16),
64997 => conv_std_logic_vector(57937, 16),
64998 => conv_std_logic_vector(58190, 16),
64999 => conv_std_logic_vector(58443, 16),
65000 => conv_std_logic_vector(58696, 16),
65001 => conv_std_logic_vector(58949, 16),
65002 => conv_std_logic_vector(59202, 16),
65003 => conv_std_logic_vector(59455, 16),
65004 => conv_std_logic_vector(59708, 16),
65005 => conv_std_logic_vector(59961, 16),
65006 => conv_std_logic_vector(60214, 16),
65007 => conv_std_logic_vector(60467, 16),
65008 => conv_std_logic_vector(60720, 16),
65009 => conv_std_logic_vector(60973, 16),
65010 => conv_std_logic_vector(61226, 16),
65011 => conv_std_logic_vector(61479, 16),
65012 => conv_std_logic_vector(61732, 16),
65013 => conv_std_logic_vector(61985, 16),
65014 => conv_std_logic_vector(62238, 16),
65015 => conv_std_logic_vector(62491, 16),
65016 => conv_std_logic_vector(62744, 16),
65017 => conv_std_logic_vector(62997, 16),
65018 => conv_std_logic_vector(63250, 16),
65019 => conv_std_logic_vector(63503, 16),
65020 => conv_std_logic_vector(63756, 16),
65021 => conv_std_logic_vector(64009, 16),
65022 => conv_std_logic_vector(64262, 16),
65023 => conv_std_logic_vector(64515, 16),
65024 => conv_std_logic_vector(0, 16),
65025 => conv_std_logic_vector(254, 16),
65026 => conv_std_logic_vector(508, 16),
65027 => conv_std_logic_vector(762, 16),
65028 => conv_std_logic_vector(1016, 16),
65029 => conv_std_logic_vector(1270, 16),
65030 => conv_std_logic_vector(1524, 16),
65031 => conv_std_logic_vector(1778, 16),
65032 => conv_std_logic_vector(2032, 16),
65033 => conv_std_logic_vector(2286, 16),
65034 => conv_std_logic_vector(2540, 16),
65035 => conv_std_logic_vector(2794, 16),
65036 => conv_std_logic_vector(3048, 16),
65037 => conv_std_logic_vector(3302, 16),
65038 => conv_std_logic_vector(3556, 16),
65039 => conv_std_logic_vector(3810, 16),
65040 => conv_std_logic_vector(4064, 16),
65041 => conv_std_logic_vector(4318, 16),
65042 => conv_std_logic_vector(4572, 16),
65043 => conv_std_logic_vector(4826, 16),
65044 => conv_std_logic_vector(5080, 16),
65045 => conv_std_logic_vector(5334, 16),
65046 => conv_std_logic_vector(5588, 16),
65047 => conv_std_logic_vector(5842, 16),
65048 => conv_std_logic_vector(6096, 16),
65049 => conv_std_logic_vector(6350, 16),
65050 => conv_std_logic_vector(6604, 16),
65051 => conv_std_logic_vector(6858, 16),
65052 => conv_std_logic_vector(7112, 16),
65053 => conv_std_logic_vector(7366, 16),
65054 => conv_std_logic_vector(7620, 16),
65055 => conv_std_logic_vector(7874, 16),
65056 => conv_std_logic_vector(8128, 16),
65057 => conv_std_logic_vector(8382, 16),
65058 => conv_std_logic_vector(8636, 16),
65059 => conv_std_logic_vector(8890, 16),
65060 => conv_std_logic_vector(9144, 16),
65061 => conv_std_logic_vector(9398, 16),
65062 => conv_std_logic_vector(9652, 16),
65063 => conv_std_logic_vector(9906, 16),
65064 => conv_std_logic_vector(10160, 16),
65065 => conv_std_logic_vector(10414, 16),
65066 => conv_std_logic_vector(10668, 16),
65067 => conv_std_logic_vector(10922, 16),
65068 => conv_std_logic_vector(11176, 16),
65069 => conv_std_logic_vector(11430, 16),
65070 => conv_std_logic_vector(11684, 16),
65071 => conv_std_logic_vector(11938, 16),
65072 => conv_std_logic_vector(12192, 16),
65073 => conv_std_logic_vector(12446, 16),
65074 => conv_std_logic_vector(12700, 16),
65075 => conv_std_logic_vector(12954, 16),
65076 => conv_std_logic_vector(13208, 16),
65077 => conv_std_logic_vector(13462, 16),
65078 => conv_std_logic_vector(13716, 16),
65079 => conv_std_logic_vector(13970, 16),
65080 => conv_std_logic_vector(14224, 16),
65081 => conv_std_logic_vector(14478, 16),
65082 => conv_std_logic_vector(14732, 16),
65083 => conv_std_logic_vector(14986, 16),
65084 => conv_std_logic_vector(15240, 16),
65085 => conv_std_logic_vector(15494, 16),
65086 => conv_std_logic_vector(15748, 16),
65087 => conv_std_logic_vector(16002, 16),
65088 => conv_std_logic_vector(16256, 16),
65089 => conv_std_logic_vector(16510, 16),
65090 => conv_std_logic_vector(16764, 16),
65091 => conv_std_logic_vector(17018, 16),
65092 => conv_std_logic_vector(17272, 16),
65093 => conv_std_logic_vector(17526, 16),
65094 => conv_std_logic_vector(17780, 16),
65095 => conv_std_logic_vector(18034, 16),
65096 => conv_std_logic_vector(18288, 16),
65097 => conv_std_logic_vector(18542, 16),
65098 => conv_std_logic_vector(18796, 16),
65099 => conv_std_logic_vector(19050, 16),
65100 => conv_std_logic_vector(19304, 16),
65101 => conv_std_logic_vector(19558, 16),
65102 => conv_std_logic_vector(19812, 16),
65103 => conv_std_logic_vector(20066, 16),
65104 => conv_std_logic_vector(20320, 16),
65105 => conv_std_logic_vector(20574, 16),
65106 => conv_std_logic_vector(20828, 16),
65107 => conv_std_logic_vector(21082, 16),
65108 => conv_std_logic_vector(21336, 16),
65109 => conv_std_logic_vector(21590, 16),
65110 => conv_std_logic_vector(21844, 16),
65111 => conv_std_logic_vector(22098, 16),
65112 => conv_std_logic_vector(22352, 16),
65113 => conv_std_logic_vector(22606, 16),
65114 => conv_std_logic_vector(22860, 16),
65115 => conv_std_logic_vector(23114, 16),
65116 => conv_std_logic_vector(23368, 16),
65117 => conv_std_logic_vector(23622, 16),
65118 => conv_std_logic_vector(23876, 16),
65119 => conv_std_logic_vector(24130, 16),
65120 => conv_std_logic_vector(24384, 16),
65121 => conv_std_logic_vector(24638, 16),
65122 => conv_std_logic_vector(24892, 16),
65123 => conv_std_logic_vector(25146, 16),
65124 => conv_std_logic_vector(25400, 16),
65125 => conv_std_logic_vector(25654, 16),
65126 => conv_std_logic_vector(25908, 16),
65127 => conv_std_logic_vector(26162, 16),
65128 => conv_std_logic_vector(26416, 16),
65129 => conv_std_logic_vector(26670, 16),
65130 => conv_std_logic_vector(26924, 16),
65131 => conv_std_logic_vector(27178, 16),
65132 => conv_std_logic_vector(27432, 16),
65133 => conv_std_logic_vector(27686, 16),
65134 => conv_std_logic_vector(27940, 16),
65135 => conv_std_logic_vector(28194, 16),
65136 => conv_std_logic_vector(28448, 16),
65137 => conv_std_logic_vector(28702, 16),
65138 => conv_std_logic_vector(28956, 16),
65139 => conv_std_logic_vector(29210, 16),
65140 => conv_std_logic_vector(29464, 16),
65141 => conv_std_logic_vector(29718, 16),
65142 => conv_std_logic_vector(29972, 16),
65143 => conv_std_logic_vector(30226, 16),
65144 => conv_std_logic_vector(30480, 16),
65145 => conv_std_logic_vector(30734, 16),
65146 => conv_std_logic_vector(30988, 16),
65147 => conv_std_logic_vector(31242, 16),
65148 => conv_std_logic_vector(31496, 16),
65149 => conv_std_logic_vector(31750, 16),
65150 => conv_std_logic_vector(32004, 16),
65151 => conv_std_logic_vector(32258, 16),
65152 => conv_std_logic_vector(32512, 16),
65153 => conv_std_logic_vector(32766, 16),
65154 => conv_std_logic_vector(33020, 16),
65155 => conv_std_logic_vector(33274, 16),
65156 => conv_std_logic_vector(33528, 16),
65157 => conv_std_logic_vector(33782, 16),
65158 => conv_std_logic_vector(34036, 16),
65159 => conv_std_logic_vector(34290, 16),
65160 => conv_std_logic_vector(34544, 16),
65161 => conv_std_logic_vector(34798, 16),
65162 => conv_std_logic_vector(35052, 16),
65163 => conv_std_logic_vector(35306, 16),
65164 => conv_std_logic_vector(35560, 16),
65165 => conv_std_logic_vector(35814, 16),
65166 => conv_std_logic_vector(36068, 16),
65167 => conv_std_logic_vector(36322, 16),
65168 => conv_std_logic_vector(36576, 16),
65169 => conv_std_logic_vector(36830, 16),
65170 => conv_std_logic_vector(37084, 16),
65171 => conv_std_logic_vector(37338, 16),
65172 => conv_std_logic_vector(37592, 16),
65173 => conv_std_logic_vector(37846, 16),
65174 => conv_std_logic_vector(38100, 16),
65175 => conv_std_logic_vector(38354, 16),
65176 => conv_std_logic_vector(38608, 16),
65177 => conv_std_logic_vector(38862, 16),
65178 => conv_std_logic_vector(39116, 16),
65179 => conv_std_logic_vector(39370, 16),
65180 => conv_std_logic_vector(39624, 16),
65181 => conv_std_logic_vector(39878, 16),
65182 => conv_std_logic_vector(40132, 16),
65183 => conv_std_logic_vector(40386, 16),
65184 => conv_std_logic_vector(40640, 16),
65185 => conv_std_logic_vector(40894, 16),
65186 => conv_std_logic_vector(41148, 16),
65187 => conv_std_logic_vector(41402, 16),
65188 => conv_std_logic_vector(41656, 16),
65189 => conv_std_logic_vector(41910, 16),
65190 => conv_std_logic_vector(42164, 16),
65191 => conv_std_logic_vector(42418, 16),
65192 => conv_std_logic_vector(42672, 16),
65193 => conv_std_logic_vector(42926, 16),
65194 => conv_std_logic_vector(43180, 16),
65195 => conv_std_logic_vector(43434, 16),
65196 => conv_std_logic_vector(43688, 16),
65197 => conv_std_logic_vector(43942, 16),
65198 => conv_std_logic_vector(44196, 16),
65199 => conv_std_logic_vector(44450, 16),
65200 => conv_std_logic_vector(44704, 16),
65201 => conv_std_logic_vector(44958, 16),
65202 => conv_std_logic_vector(45212, 16),
65203 => conv_std_logic_vector(45466, 16),
65204 => conv_std_logic_vector(45720, 16),
65205 => conv_std_logic_vector(45974, 16),
65206 => conv_std_logic_vector(46228, 16),
65207 => conv_std_logic_vector(46482, 16),
65208 => conv_std_logic_vector(46736, 16),
65209 => conv_std_logic_vector(46990, 16),
65210 => conv_std_logic_vector(47244, 16),
65211 => conv_std_logic_vector(47498, 16),
65212 => conv_std_logic_vector(47752, 16),
65213 => conv_std_logic_vector(48006, 16),
65214 => conv_std_logic_vector(48260, 16),
65215 => conv_std_logic_vector(48514, 16),
65216 => conv_std_logic_vector(48768, 16),
65217 => conv_std_logic_vector(49022, 16),
65218 => conv_std_logic_vector(49276, 16),
65219 => conv_std_logic_vector(49530, 16),
65220 => conv_std_logic_vector(49784, 16),
65221 => conv_std_logic_vector(50038, 16),
65222 => conv_std_logic_vector(50292, 16),
65223 => conv_std_logic_vector(50546, 16),
65224 => conv_std_logic_vector(50800, 16),
65225 => conv_std_logic_vector(51054, 16),
65226 => conv_std_logic_vector(51308, 16),
65227 => conv_std_logic_vector(51562, 16),
65228 => conv_std_logic_vector(51816, 16),
65229 => conv_std_logic_vector(52070, 16),
65230 => conv_std_logic_vector(52324, 16),
65231 => conv_std_logic_vector(52578, 16),
65232 => conv_std_logic_vector(52832, 16),
65233 => conv_std_logic_vector(53086, 16),
65234 => conv_std_logic_vector(53340, 16),
65235 => conv_std_logic_vector(53594, 16),
65236 => conv_std_logic_vector(53848, 16),
65237 => conv_std_logic_vector(54102, 16),
65238 => conv_std_logic_vector(54356, 16),
65239 => conv_std_logic_vector(54610, 16),
65240 => conv_std_logic_vector(54864, 16),
65241 => conv_std_logic_vector(55118, 16),
65242 => conv_std_logic_vector(55372, 16),
65243 => conv_std_logic_vector(55626, 16),
65244 => conv_std_logic_vector(55880, 16),
65245 => conv_std_logic_vector(56134, 16),
65246 => conv_std_logic_vector(56388, 16),
65247 => conv_std_logic_vector(56642, 16),
65248 => conv_std_logic_vector(56896, 16),
65249 => conv_std_logic_vector(57150, 16),
65250 => conv_std_logic_vector(57404, 16),
65251 => conv_std_logic_vector(57658, 16),
65252 => conv_std_logic_vector(57912, 16),
65253 => conv_std_logic_vector(58166, 16),
65254 => conv_std_logic_vector(58420, 16),
65255 => conv_std_logic_vector(58674, 16),
65256 => conv_std_logic_vector(58928, 16),
65257 => conv_std_logic_vector(59182, 16),
65258 => conv_std_logic_vector(59436, 16),
65259 => conv_std_logic_vector(59690, 16),
65260 => conv_std_logic_vector(59944, 16),
65261 => conv_std_logic_vector(60198, 16),
65262 => conv_std_logic_vector(60452, 16),
65263 => conv_std_logic_vector(60706, 16),
65264 => conv_std_logic_vector(60960, 16),
65265 => conv_std_logic_vector(61214, 16),
65266 => conv_std_logic_vector(61468, 16),
65267 => conv_std_logic_vector(61722, 16),
65268 => conv_std_logic_vector(61976, 16),
65269 => conv_std_logic_vector(62230, 16),
65270 => conv_std_logic_vector(62484, 16),
65271 => conv_std_logic_vector(62738, 16),
65272 => conv_std_logic_vector(62992, 16),
65273 => conv_std_logic_vector(63246, 16),
65274 => conv_std_logic_vector(63500, 16),
65275 => conv_std_logic_vector(63754, 16),
65276 => conv_std_logic_vector(64008, 16),
65277 => conv_std_logic_vector(64262, 16),
65278 => conv_std_logic_vector(64516, 16),
65279 => conv_std_logic_vector(64770, 16),
65280 => conv_std_logic_vector(0, 16),
65281 => conv_std_logic_vector(255, 16),
65282 => conv_std_logic_vector(510, 16),
65283 => conv_std_logic_vector(765, 16),
65284 => conv_std_logic_vector(1020, 16),
65285 => conv_std_logic_vector(1275, 16),
65286 => conv_std_logic_vector(1530, 16),
65287 => conv_std_logic_vector(1785, 16),
65288 => conv_std_logic_vector(2040, 16),
65289 => conv_std_logic_vector(2295, 16),
65290 => conv_std_logic_vector(2550, 16),
65291 => conv_std_logic_vector(2805, 16),
65292 => conv_std_logic_vector(3060, 16),
65293 => conv_std_logic_vector(3315, 16),
65294 => conv_std_logic_vector(3570, 16),
65295 => conv_std_logic_vector(3825, 16),
65296 => conv_std_logic_vector(4080, 16),
65297 => conv_std_logic_vector(4335, 16),
65298 => conv_std_logic_vector(4590, 16),
65299 => conv_std_logic_vector(4845, 16),
65300 => conv_std_logic_vector(5100, 16),
65301 => conv_std_logic_vector(5355, 16),
65302 => conv_std_logic_vector(5610, 16),
65303 => conv_std_logic_vector(5865, 16),
65304 => conv_std_logic_vector(6120, 16),
65305 => conv_std_logic_vector(6375, 16),
65306 => conv_std_logic_vector(6630, 16),
65307 => conv_std_logic_vector(6885, 16),
65308 => conv_std_logic_vector(7140, 16),
65309 => conv_std_logic_vector(7395, 16),
65310 => conv_std_logic_vector(7650, 16),
65311 => conv_std_logic_vector(7905, 16),
65312 => conv_std_logic_vector(8160, 16),
65313 => conv_std_logic_vector(8415, 16),
65314 => conv_std_logic_vector(8670, 16),
65315 => conv_std_logic_vector(8925, 16),
65316 => conv_std_logic_vector(9180, 16),
65317 => conv_std_logic_vector(9435, 16),
65318 => conv_std_logic_vector(9690, 16),
65319 => conv_std_logic_vector(9945, 16),
65320 => conv_std_logic_vector(10200, 16),
65321 => conv_std_logic_vector(10455, 16),
65322 => conv_std_logic_vector(10710, 16),
65323 => conv_std_logic_vector(10965, 16),
65324 => conv_std_logic_vector(11220, 16),
65325 => conv_std_logic_vector(11475, 16),
65326 => conv_std_logic_vector(11730, 16),
65327 => conv_std_logic_vector(11985, 16),
65328 => conv_std_logic_vector(12240, 16),
65329 => conv_std_logic_vector(12495, 16),
65330 => conv_std_logic_vector(12750, 16),
65331 => conv_std_logic_vector(13005, 16),
65332 => conv_std_logic_vector(13260, 16),
65333 => conv_std_logic_vector(13515, 16),
65334 => conv_std_logic_vector(13770, 16),
65335 => conv_std_logic_vector(14025, 16),
65336 => conv_std_logic_vector(14280, 16),
65337 => conv_std_logic_vector(14535, 16),
65338 => conv_std_logic_vector(14790, 16),
65339 => conv_std_logic_vector(15045, 16),
65340 => conv_std_logic_vector(15300, 16),
65341 => conv_std_logic_vector(15555, 16),
65342 => conv_std_logic_vector(15810, 16),
65343 => conv_std_logic_vector(16065, 16),
65344 => conv_std_logic_vector(16320, 16),
65345 => conv_std_logic_vector(16575, 16),
65346 => conv_std_logic_vector(16830, 16),
65347 => conv_std_logic_vector(17085, 16),
65348 => conv_std_logic_vector(17340, 16),
65349 => conv_std_logic_vector(17595, 16),
65350 => conv_std_logic_vector(17850, 16),
65351 => conv_std_logic_vector(18105, 16),
65352 => conv_std_logic_vector(18360, 16),
65353 => conv_std_logic_vector(18615, 16),
65354 => conv_std_logic_vector(18870, 16),
65355 => conv_std_logic_vector(19125, 16),
65356 => conv_std_logic_vector(19380, 16),
65357 => conv_std_logic_vector(19635, 16),
65358 => conv_std_logic_vector(19890, 16),
65359 => conv_std_logic_vector(20145, 16),
65360 => conv_std_logic_vector(20400, 16),
65361 => conv_std_logic_vector(20655, 16),
65362 => conv_std_logic_vector(20910, 16),
65363 => conv_std_logic_vector(21165, 16),
65364 => conv_std_logic_vector(21420, 16),
65365 => conv_std_logic_vector(21675, 16),
65366 => conv_std_logic_vector(21930, 16),
65367 => conv_std_logic_vector(22185, 16),
65368 => conv_std_logic_vector(22440, 16),
65369 => conv_std_logic_vector(22695, 16),
65370 => conv_std_logic_vector(22950, 16),
65371 => conv_std_logic_vector(23205, 16),
65372 => conv_std_logic_vector(23460, 16),
65373 => conv_std_logic_vector(23715, 16),
65374 => conv_std_logic_vector(23970, 16),
65375 => conv_std_logic_vector(24225, 16),
65376 => conv_std_logic_vector(24480, 16),
65377 => conv_std_logic_vector(24735, 16),
65378 => conv_std_logic_vector(24990, 16),
65379 => conv_std_logic_vector(25245, 16),
65380 => conv_std_logic_vector(25500, 16),
65381 => conv_std_logic_vector(25755, 16),
65382 => conv_std_logic_vector(26010, 16),
65383 => conv_std_logic_vector(26265, 16),
65384 => conv_std_logic_vector(26520, 16),
65385 => conv_std_logic_vector(26775, 16),
65386 => conv_std_logic_vector(27030, 16),
65387 => conv_std_logic_vector(27285, 16),
65388 => conv_std_logic_vector(27540, 16),
65389 => conv_std_logic_vector(27795, 16),
65390 => conv_std_logic_vector(28050, 16),
65391 => conv_std_logic_vector(28305, 16),
65392 => conv_std_logic_vector(28560, 16),
65393 => conv_std_logic_vector(28815, 16),
65394 => conv_std_logic_vector(29070, 16),
65395 => conv_std_logic_vector(29325, 16),
65396 => conv_std_logic_vector(29580, 16),
65397 => conv_std_logic_vector(29835, 16),
65398 => conv_std_logic_vector(30090, 16),
65399 => conv_std_logic_vector(30345, 16),
65400 => conv_std_logic_vector(30600, 16),
65401 => conv_std_logic_vector(30855, 16),
65402 => conv_std_logic_vector(31110, 16),
65403 => conv_std_logic_vector(31365, 16),
65404 => conv_std_logic_vector(31620, 16),
65405 => conv_std_logic_vector(31875, 16),
65406 => conv_std_logic_vector(32130, 16),
65407 => conv_std_logic_vector(32385, 16),
65408 => conv_std_logic_vector(32640, 16),
65409 => conv_std_logic_vector(32895, 16),
65410 => conv_std_logic_vector(33150, 16),
65411 => conv_std_logic_vector(33405, 16),
65412 => conv_std_logic_vector(33660, 16),
65413 => conv_std_logic_vector(33915, 16),
65414 => conv_std_logic_vector(34170, 16),
65415 => conv_std_logic_vector(34425, 16),
65416 => conv_std_logic_vector(34680, 16),
65417 => conv_std_logic_vector(34935, 16),
65418 => conv_std_logic_vector(35190, 16),
65419 => conv_std_logic_vector(35445, 16),
65420 => conv_std_logic_vector(35700, 16),
65421 => conv_std_logic_vector(35955, 16),
65422 => conv_std_logic_vector(36210, 16),
65423 => conv_std_logic_vector(36465, 16),
65424 => conv_std_logic_vector(36720, 16),
65425 => conv_std_logic_vector(36975, 16),
65426 => conv_std_logic_vector(37230, 16),
65427 => conv_std_logic_vector(37485, 16),
65428 => conv_std_logic_vector(37740, 16),
65429 => conv_std_logic_vector(37995, 16),
65430 => conv_std_logic_vector(38250, 16),
65431 => conv_std_logic_vector(38505, 16),
65432 => conv_std_logic_vector(38760, 16),
65433 => conv_std_logic_vector(39015, 16),
65434 => conv_std_logic_vector(39270, 16),
65435 => conv_std_logic_vector(39525, 16),
65436 => conv_std_logic_vector(39780, 16),
65437 => conv_std_logic_vector(40035, 16),
65438 => conv_std_logic_vector(40290, 16),
65439 => conv_std_logic_vector(40545, 16),
65440 => conv_std_logic_vector(40800, 16),
65441 => conv_std_logic_vector(41055, 16),
65442 => conv_std_logic_vector(41310, 16),
65443 => conv_std_logic_vector(41565, 16),
65444 => conv_std_logic_vector(41820, 16),
65445 => conv_std_logic_vector(42075, 16),
65446 => conv_std_logic_vector(42330, 16),
65447 => conv_std_logic_vector(42585, 16),
65448 => conv_std_logic_vector(42840, 16),
65449 => conv_std_logic_vector(43095, 16),
65450 => conv_std_logic_vector(43350, 16),
65451 => conv_std_logic_vector(43605, 16),
65452 => conv_std_logic_vector(43860, 16),
65453 => conv_std_logic_vector(44115, 16),
65454 => conv_std_logic_vector(44370, 16),
65455 => conv_std_logic_vector(44625, 16),
65456 => conv_std_logic_vector(44880, 16),
65457 => conv_std_logic_vector(45135, 16),
65458 => conv_std_logic_vector(45390, 16),
65459 => conv_std_logic_vector(45645, 16),
65460 => conv_std_logic_vector(45900, 16),
65461 => conv_std_logic_vector(46155, 16),
65462 => conv_std_logic_vector(46410, 16),
65463 => conv_std_logic_vector(46665, 16),
65464 => conv_std_logic_vector(46920, 16),
65465 => conv_std_logic_vector(47175, 16),
65466 => conv_std_logic_vector(47430, 16),
65467 => conv_std_logic_vector(47685, 16),
65468 => conv_std_logic_vector(47940, 16),
65469 => conv_std_logic_vector(48195, 16),
65470 => conv_std_logic_vector(48450, 16),
65471 => conv_std_logic_vector(48705, 16),
65472 => conv_std_logic_vector(48960, 16),
65473 => conv_std_logic_vector(49215, 16),
65474 => conv_std_logic_vector(49470, 16),
65475 => conv_std_logic_vector(49725, 16),
65476 => conv_std_logic_vector(49980, 16),
65477 => conv_std_logic_vector(50235, 16),
65478 => conv_std_logic_vector(50490, 16),
65479 => conv_std_logic_vector(50745, 16),
65480 => conv_std_logic_vector(51000, 16),
65481 => conv_std_logic_vector(51255, 16),
65482 => conv_std_logic_vector(51510, 16),
65483 => conv_std_logic_vector(51765, 16),
65484 => conv_std_logic_vector(52020, 16),
65485 => conv_std_logic_vector(52275, 16),
65486 => conv_std_logic_vector(52530, 16),
65487 => conv_std_logic_vector(52785, 16),
65488 => conv_std_logic_vector(53040, 16),
65489 => conv_std_logic_vector(53295, 16),
65490 => conv_std_logic_vector(53550, 16),
65491 => conv_std_logic_vector(53805, 16),
65492 => conv_std_logic_vector(54060, 16),
65493 => conv_std_logic_vector(54315, 16),
65494 => conv_std_logic_vector(54570, 16),
65495 => conv_std_logic_vector(54825, 16),
65496 => conv_std_logic_vector(55080, 16),
65497 => conv_std_logic_vector(55335, 16),
65498 => conv_std_logic_vector(55590, 16),
65499 => conv_std_logic_vector(55845, 16),
65500 => conv_std_logic_vector(56100, 16),
65501 => conv_std_logic_vector(56355, 16),
65502 => conv_std_logic_vector(56610, 16),
65503 => conv_std_logic_vector(56865, 16),
65504 => conv_std_logic_vector(57120, 16),
65505 => conv_std_logic_vector(57375, 16),
65506 => conv_std_logic_vector(57630, 16),
65507 => conv_std_logic_vector(57885, 16),
65508 => conv_std_logic_vector(58140, 16),
65509 => conv_std_logic_vector(58395, 16),
65510 => conv_std_logic_vector(58650, 16),
65511 => conv_std_logic_vector(58905, 16),
65512 => conv_std_logic_vector(59160, 16),
65513 => conv_std_logic_vector(59415, 16),
65514 => conv_std_logic_vector(59670, 16),
65515 => conv_std_logic_vector(59925, 16),
65516 => conv_std_logic_vector(60180, 16),
65517 => conv_std_logic_vector(60435, 16),
65518 => conv_std_logic_vector(60690, 16),
65519 => conv_std_logic_vector(60945, 16),
65520 => conv_std_logic_vector(61200, 16),
65521 => conv_std_logic_vector(61455, 16),
65522 => conv_std_logic_vector(61710, 16),
65523 => conv_std_logic_vector(61965, 16),
65524 => conv_std_logic_vector(62220, 16),
65525 => conv_std_logic_vector(62475, 16),
65526 => conv_std_logic_vector(62730, 16),
65527 => conv_std_logic_vector(62985, 16),
65528 => conv_std_logic_vector(63240, 16),
65529 => conv_std_logic_vector(63495, 16),
65530 => conv_std_logic_vector(63750, 16),
65531 => conv_std_logic_vector(64005, 16),
65532 => conv_std_logic_vector(64260, 16),
65533 => conv_std_logic_vector(64515, 16),
65534 => conv_std_logic_vector(64770, 16),
65535 => conv_std_logic_vector(65025, 16),
 OTHERS => conv_std_logic_vector( 0, 16)
  );       

begin
    process(clk)
    begin
       if( clk'event and clk = '1' ) then
          ROM_data <= Content(conv_integer(ROM_addr));
       end if;
    end process;
end a;